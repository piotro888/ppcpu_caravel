// This is the unpowered netlist.
module core1 (i_clk,
    i_disable,
    i_irq,
    i_mc_core_int,
    i_mem_ack,
    i_mem_exception,
    i_req_data_valid,
    i_rst,
    o_c_data_page,
    o_c_instr_long,
    o_c_instr_page,
    o_icache_flush,
    o_mem_long,
    o_mem_req,
    o_mem_we,
    o_req_active,
    o_req_ppl_submit,
    sr_bus_we,
    dbg_in,
    dbg_out,
    dbg_pc,
    dbg_r0,
    i_core_int_sreg,
    i_mem_data,
    i_req_data,
    o_instr_long_addr,
    o_mem_addr,
    o_mem_addr_high,
    o_mem_data,
    o_mem_sel,
    o_req_addr,
    sr_bus_addr,
    sr_bus_data_o);
 input i_clk;
 input i_disable;
 input i_irq;
 input i_mc_core_int;
 input i_mem_ack;
 input i_mem_exception;
 input i_req_data_valid;
 input i_rst;
 output o_c_data_page;
 output o_c_instr_long;
 output o_c_instr_page;
 output o_icache_flush;
 output o_mem_long;
 output o_mem_req;
 output o_mem_we;
 output o_req_active;
 output o_req_ppl_submit;
 output sr_bus_we;
 input [3:0] dbg_in;
 output [35:0] dbg_out;
 output [15:0] dbg_pc;
 output [15:0] dbg_r0;
 input [15:0] i_core_int_sreg;
 input [15:0] i_mem_data;
 input [31:0] i_req_data;
 output [7:0] o_instr_long_addr;
 output [15:0] o_mem_addr;
 output [7:0] o_mem_addr_high;
 output [15:0] o_mem_data;
 output [1:0] o_mem_sel;
 output [15:0] o_req_addr;
 output [15:0] sr_bus_addr;
 output [15:0] sr_bus_data_o;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire \core_1.de_jmp_pred ;
 wire \core_1.dec_alu_carry_en ;
 wire \core_1.dec_alu_flags_ie ;
 wire \core_1.dec_jump_cond_code[0] ;
 wire \core_1.dec_jump_cond_code[1] ;
 wire \core_1.dec_jump_cond_code[2] ;
 wire \core_1.dec_jump_cond_code[3] ;
 wire \core_1.dec_jump_cond_code[4] ;
 wire \core_1.dec_l_reg_sel[0] ;
 wire \core_1.dec_l_reg_sel[1] ;
 wire \core_1.dec_l_reg_sel[2] ;
 wire \core_1.dec_mem_access ;
 wire \core_1.dec_mem_long ;
 wire \core_1.dec_mem_we ;
 wire \core_1.dec_mem_width ;
 wire \core_1.dec_pc_inc ;
 wire \core_1.dec_r_bus_imm ;
 wire \core_1.dec_r_reg_sel[0] ;
 wire \core_1.dec_r_reg_sel[1] ;
 wire \core_1.dec_r_reg_sel[2] ;
 wire \core_1.dec_rf_ie[0] ;
 wire \core_1.dec_rf_ie[1] ;
 wire \core_1.dec_rf_ie[2] ;
 wire \core_1.dec_rf_ie[3] ;
 wire \core_1.dec_rf_ie[4] ;
 wire \core_1.dec_rf_ie[5] ;
 wire \core_1.dec_rf_ie[6] ;
 wire \core_1.dec_rf_ie[7] ;
 wire \core_1.dec_sreg_irt ;
 wire \core_1.dec_sreg_jal_over ;
 wire \core_1.dec_sreg_load ;
 wire \core_1.dec_sreg_store ;
 wire \core_1.dec_sys ;
 wire \core_1.dec_used_operands[0] ;
 wire \core_1.dec_used_operands[1] ;
 wire \core_1.decode.i_flush ;
 wire \core_1.decode.i_imm_pass[0] ;
 wire \core_1.decode.i_imm_pass[10] ;
 wire \core_1.decode.i_imm_pass[11] ;
 wire \core_1.decode.i_imm_pass[12] ;
 wire \core_1.decode.i_imm_pass[13] ;
 wire \core_1.decode.i_imm_pass[14] ;
 wire \core_1.decode.i_imm_pass[15] ;
 wire \core_1.decode.i_imm_pass[1] ;
 wire \core_1.decode.i_imm_pass[2] ;
 wire \core_1.decode.i_imm_pass[3] ;
 wire \core_1.decode.i_imm_pass[4] ;
 wire \core_1.decode.i_imm_pass[5] ;
 wire \core_1.decode.i_imm_pass[6] ;
 wire \core_1.decode.i_imm_pass[7] ;
 wire \core_1.decode.i_imm_pass[8] ;
 wire \core_1.decode.i_imm_pass[9] ;
 wire \core_1.decode.i_instr_l[0] ;
 wire \core_1.decode.i_instr_l[10] ;
 wire \core_1.decode.i_instr_l[11] ;
 wire \core_1.decode.i_instr_l[12] ;
 wire \core_1.decode.i_instr_l[13] ;
 wire \core_1.decode.i_instr_l[14] ;
 wire \core_1.decode.i_instr_l[15] ;
 wire \core_1.decode.i_instr_l[1] ;
 wire \core_1.decode.i_instr_l[2] ;
 wire \core_1.decode.i_instr_l[3] ;
 wire \core_1.decode.i_instr_l[4] ;
 wire \core_1.decode.i_instr_l[5] ;
 wire \core_1.decode.i_instr_l[6] ;
 wire \core_1.decode.i_instr_l[7] ;
 wire \core_1.decode.i_instr_l[8] ;
 wire \core_1.decode.i_instr_l[9] ;
 wire \core_1.decode.i_jmp_pred_pass ;
 wire \core_1.decode.i_submit ;
 wire \core_1.decode.input_valid ;
 wire \core_1.decode.o_submit ;
 wire \core_1.decode.oc_alu_mode[11] ;
 wire \core_1.decode.oc_alu_mode[12] ;
 wire \core_1.decode.oc_alu_mode[13] ;
 wire \core_1.decode.oc_alu_mode[1] ;
 wire \core_1.decode.oc_alu_mode[2] ;
 wire \core_1.decode.oc_alu_mode[3] ;
 wire \core_1.decode.oc_alu_mode[4] ;
 wire \core_1.decode.oc_alu_mode[6] ;
 wire \core_1.decode.oc_alu_mode[7] ;
 wire \core_1.decode.oc_alu_mode[9] ;
 wire \core_1.ew_addr[0] ;
 wire \core_1.ew_addr_high[0] ;
 wire \core_1.ew_data[0] ;
 wire \core_1.ew_data[10] ;
 wire \core_1.ew_data[11] ;
 wire \core_1.ew_data[12] ;
 wire \core_1.ew_data[13] ;
 wire \core_1.ew_data[14] ;
 wire \core_1.ew_data[15] ;
 wire \core_1.ew_data[1] ;
 wire \core_1.ew_data[2] ;
 wire \core_1.ew_data[3] ;
 wire \core_1.ew_data[4] ;
 wire \core_1.ew_data[5] ;
 wire \core_1.ew_data[6] ;
 wire \core_1.ew_data[7] ;
 wire \core_1.ew_data[8] ;
 wire \core_1.ew_data[9] ;
 wire \core_1.ew_mem_access ;
 wire \core_1.ew_mem_width ;
 wire \core_1.ew_reg_ie[0] ;
 wire \core_1.ew_reg_ie[1] ;
 wire \core_1.ew_reg_ie[2] ;
 wire \core_1.ew_reg_ie[3] ;
 wire \core_1.ew_reg_ie[4] ;
 wire \core_1.ew_reg_ie[5] ;
 wire \core_1.ew_reg_ie[6] ;
 wire \core_1.ew_reg_ie[7] ;
 wire \core_1.ew_submit ;
 wire \core_1.execute.alu_flag_reg.o_d[0] ;
 wire \core_1.execute.alu_flag_reg.o_d[1] ;
 wire \core_1.execute.alu_flag_reg.o_d[2] ;
 wire \core_1.execute.alu_flag_reg.o_d[3] ;
 wire \core_1.execute.alu_flag_reg.o_d[4] ;
 wire \core_1.execute.alu_mul_div.cbit[0] ;
 wire \core_1.execute.alu_mul_div.cbit[1] ;
 wire \core_1.execute.alu_mul_div.cbit[2] ;
 wire \core_1.execute.alu_mul_div.cbit[3] ;
 wire \core_1.execute.alu_mul_div.comp ;
 wire \core_1.execute.alu_mul_div.div_cur[0] ;
 wire \core_1.execute.alu_mul_div.div_cur[10] ;
 wire \core_1.execute.alu_mul_div.div_cur[11] ;
 wire \core_1.execute.alu_mul_div.div_cur[12] ;
 wire \core_1.execute.alu_mul_div.div_cur[13] ;
 wire \core_1.execute.alu_mul_div.div_cur[14] ;
 wire \core_1.execute.alu_mul_div.div_cur[15] ;
 wire \core_1.execute.alu_mul_div.div_cur[1] ;
 wire \core_1.execute.alu_mul_div.div_cur[2] ;
 wire \core_1.execute.alu_mul_div.div_cur[3] ;
 wire \core_1.execute.alu_mul_div.div_cur[4] ;
 wire \core_1.execute.alu_mul_div.div_cur[5] ;
 wire \core_1.execute.alu_mul_div.div_cur[6] ;
 wire \core_1.execute.alu_mul_div.div_cur[7] ;
 wire \core_1.execute.alu_mul_div.div_cur[8] ;
 wire \core_1.execute.alu_mul_div.div_cur[9] ;
 wire \core_1.execute.alu_mul_div.div_res[0] ;
 wire \core_1.execute.alu_mul_div.div_res[10] ;
 wire \core_1.execute.alu_mul_div.div_res[11] ;
 wire \core_1.execute.alu_mul_div.div_res[12] ;
 wire \core_1.execute.alu_mul_div.div_res[13] ;
 wire \core_1.execute.alu_mul_div.div_res[14] ;
 wire \core_1.execute.alu_mul_div.div_res[15] ;
 wire \core_1.execute.alu_mul_div.div_res[1] ;
 wire \core_1.execute.alu_mul_div.div_res[2] ;
 wire \core_1.execute.alu_mul_div.div_res[3] ;
 wire \core_1.execute.alu_mul_div.div_res[4] ;
 wire \core_1.execute.alu_mul_div.div_res[5] ;
 wire \core_1.execute.alu_mul_div.div_res[6] ;
 wire \core_1.execute.alu_mul_div.div_res[7] ;
 wire \core_1.execute.alu_mul_div.div_res[8] ;
 wire \core_1.execute.alu_mul_div.div_res[9] ;
 wire \core_1.execute.alu_mul_div.i_div ;
 wire \core_1.execute.alu_mul_div.i_mod ;
 wire \core_1.execute.alu_mul_div.i_mul ;
 wire \core_1.execute.alu_mul_div.mul_res[0] ;
 wire \core_1.execute.alu_mul_div.mul_res[10] ;
 wire \core_1.execute.alu_mul_div.mul_res[11] ;
 wire \core_1.execute.alu_mul_div.mul_res[12] ;
 wire \core_1.execute.alu_mul_div.mul_res[13] ;
 wire \core_1.execute.alu_mul_div.mul_res[14] ;
 wire \core_1.execute.alu_mul_div.mul_res[15] ;
 wire \core_1.execute.alu_mul_div.mul_res[1] ;
 wire \core_1.execute.alu_mul_div.mul_res[2] ;
 wire \core_1.execute.alu_mul_div.mul_res[3] ;
 wire \core_1.execute.alu_mul_div.mul_res[4] ;
 wire \core_1.execute.alu_mul_div.mul_res[5] ;
 wire \core_1.execute.alu_mul_div.mul_res[6] ;
 wire \core_1.execute.alu_mul_div.mul_res[7] ;
 wire \core_1.execute.alu_mul_div.mul_res[8] ;
 wire \core_1.execute.alu_mul_div.mul_res[9] ;
 wire \core_1.execute.hold_valid ;
 wire \core_1.execute.irq_en ;
 wire \core_1.execute.mem_stage_pc[0] ;
 wire \core_1.execute.mem_stage_pc[10] ;
 wire \core_1.execute.mem_stage_pc[11] ;
 wire \core_1.execute.mem_stage_pc[12] ;
 wire \core_1.execute.mem_stage_pc[13] ;
 wire \core_1.execute.mem_stage_pc[14] ;
 wire \core_1.execute.mem_stage_pc[15] ;
 wire \core_1.execute.mem_stage_pc[1] ;
 wire \core_1.execute.mem_stage_pc[2] ;
 wire \core_1.execute.mem_stage_pc[3] ;
 wire \core_1.execute.mem_stage_pc[4] ;
 wire \core_1.execute.mem_stage_pc[5] ;
 wire \core_1.execute.mem_stage_pc[6] ;
 wire \core_1.execute.mem_stage_pc[7] ;
 wire \core_1.execute.mem_stage_pc[8] ;
 wire \core_1.execute.mem_stage_pc[9] ;
 wire \core_1.execute.next_ready_delayed ;
 wire \core_1.execute.pc_high_buff_out[0] ;
 wire \core_1.execute.pc_high_buff_out[1] ;
 wire \core_1.execute.pc_high_buff_out[2] ;
 wire \core_1.execute.pc_high_buff_out[3] ;
 wire \core_1.execute.pc_high_buff_out[4] ;
 wire \core_1.execute.pc_high_buff_out[5] ;
 wire \core_1.execute.pc_high_buff_out[6] ;
 wire \core_1.execute.pc_high_buff_out[7] ;
 wire \core_1.execute.pc_high_out[0] ;
 wire \core_1.execute.pc_high_out[1] ;
 wire \core_1.execute.pc_high_out[2] ;
 wire \core_1.execute.pc_high_out[3] ;
 wire \core_1.execute.pc_high_out[4] ;
 wire \core_1.execute.pc_high_out[5] ;
 wire \core_1.execute.pc_high_out[6] ;
 wire \core_1.execute.pc_high_out[7] ;
 wire \core_1.execute.prev_pc_high[0] ;
 wire \core_1.execute.prev_pc_high[1] ;
 wire \core_1.execute.prev_pc_high[2] ;
 wire \core_1.execute.prev_pc_high[3] ;
 wire \core_1.execute.prev_pc_high[4] ;
 wire \core_1.execute.prev_pc_high[5] ;
 wire \core_1.execute.prev_pc_high[6] ;
 wire \core_1.execute.prev_pc_high[7] ;
 wire \core_1.execute.prev_sys ;
 wire \core_1.execute.rf.reg_outputs[1][0] ;
 wire \core_1.execute.rf.reg_outputs[1][10] ;
 wire \core_1.execute.rf.reg_outputs[1][11] ;
 wire \core_1.execute.rf.reg_outputs[1][12] ;
 wire \core_1.execute.rf.reg_outputs[1][13] ;
 wire \core_1.execute.rf.reg_outputs[1][14] ;
 wire \core_1.execute.rf.reg_outputs[1][15] ;
 wire \core_1.execute.rf.reg_outputs[1][1] ;
 wire \core_1.execute.rf.reg_outputs[1][2] ;
 wire \core_1.execute.rf.reg_outputs[1][3] ;
 wire \core_1.execute.rf.reg_outputs[1][4] ;
 wire \core_1.execute.rf.reg_outputs[1][5] ;
 wire \core_1.execute.rf.reg_outputs[1][6] ;
 wire \core_1.execute.rf.reg_outputs[1][7] ;
 wire \core_1.execute.rf.reg_outputs[1][8] ;
 wire \core_1.execute.rf.reg_outputs[1][9] ;
 wire \core_1.execute.rf.reg_outputs[2][0] ;
 wire \core_1.execute.rf.reg_outputs[2][10] ;
 wire \core_1.execute.rf.reg_outputs[2][11] ;
 wire \core_1.execute.rf.reg_outputs[2][12] ;
 wire \core_1.execute.rf.reg_outputs[2][13] ;
 wire \core_1.execute.rf.reg_outputs[2][14] ;
 wire \core_1.execute.rf.reg_outputs[2][15] ;
 wire \core_1.execute.rf.reg_outputs[2][1] ;
 wire \core_1.execute.rf.reg_outputs[2][2] ;
 wire \core_1.execute.rf.reg_outputs[2][3] ;
 wire \core_1.execute.rf.reg_outputs[2][4] ;
 wire \core_1.execute.rf.reg_outputs[2][5] ;
 wire \core_1.execute.rf.reg_outputs[2][6] ;
 wire \core_1.execute.rf.reg_outputs[2][7] ;
 wire \core_1.execute.rf.reg_outputs[2][8] ;
 wire \core_1.execute.rf.reg_outputs[2][9] ;
 wire \core_1.execute.rf.reg_outputs[3][0] ;
 wire \core_1.execute.rf.reg_outputs[3][10] ;
 wire \core_1.execute.rf.reg_outputs[3][11] ;
 wire \core_1.execute.rf.reg_outputs[3][12] ;
 wire \core_1.execute.rf.reg_outputs[3][13] ;
 wire \core_1.execute.rf.reg_outputs[3][14] ;
 wire \core_1.execute.rf.reg_outputs[3][15] ;
 wire \core_1.execute.rf.reg_outputs[3][1] ;
 wire \core_1.execute.rf.reg_outputs[3][2] ;
 wire \core_1.execute.rf.reg_outputs[3][3] ;
 wire \core_1.execute.rf.reg_outputs[3][4] ;
 wire \core_1.execute.rf.reg_outputs[3][5] ;
 wire \core_1.execute.rf.reg_outputs[3][6] ;
 wire \core_1.execute.rf.reg_outputs[3][7] ;
 wire \core_1.execute.rf.reg_outputs[3][8] ;
 wire \core_1.execute.rf.reg_outputs[3][9] ;
 wire \core_1.execute.rf.reg_outputs[4][0] ;
 wire \core_1.execute.rf.reg_outputs[4][10] ;
 wire \core_1.execute.rf.reg_outputs[4][11] ;
 wire \core_1.execute.rf.reg_outputs[4][12] ;
 wire \core_1.execute.rf.reg_outputs[4][13] ;
 wire \core_1.execute.rf.reg_outputs[4][14] ;
 wire \core_1.execute.rf.reg_outputs[4][15] ;
 wire \core_1.execute.rf.reg_outputs[4][1] ;
 wire \core_1.execute.rf.reg_outputs[4][2] ;
 wire \core_1.execute.rf.reg_outputs[4][3] ;
 wire \core_1.execute.rf.reg_outputs[4][4] ;
 wire \core_1.execute.rf.reg_outputs[4][5] ;
 wire \core_1.execute.rf.reg_outputs[4][6] ;
 wire \core_1.execute.rf.reg_outputs[4][7] ;
 wire \core_1.execute.rf.reg_outputs[4][8] ;
 wire \core_1.execute.rf.reg_outputs[4][9] ;
 wire \core_1.execute.rf.reg_outputs[5][0] ;
 wire \core_1.execute.rf.reg_outputs[5][10] ;
 wire \core_1.execute.rf.reg_outputs[5][11] ;
 wire \core_1.execute.rf.reg_outputs[5][12] ;
 wire \core_1.execute.rf.reg_outputs[5][13] ;
 wire \core_1.execute.rf.reg_outputs[5][14] ;
 wire \core_1.execute.rf.reg_outputs[5][15] ;
 wire \core_1.execute.rf.reg_outputs[5][1] ;
 wire \core_1.execute.rf.reg_outputs[5][2] ;
 wire \core_1.execute.rf.reg_outputs[5][3] ;
 wire \core_1.execute.rf.reg_outputs[5][4] ;
 wire \core_1.execute.rf.reg_outputs[5][5] ;
 wire \core_1.execute.rf.reg_outputs[5][6] ;
 wire \core_1.execute.rf.reg_outputs[5][7] ;
 wire \core_1.execute.rf.reg_outputs[5][8] ;
 wire \core_1.execute.rf.reg_outputs[5][9] ;
 wire \core_1.execute.rf.reg_outputs[6][0] ;
 wire \core_1.execute.rf.reg_outputs[6][10] ;
 wire \core_1.execute.rf.reg_outputs[6][11] ;
 wire \core_1.execute.rf.reg_outputs[6][12] ;
 wire \core_1.execute.rf.reg_outputs[6][13] ;
 wire \core_1.execute.rf.reg_outputs[6][14] ;
 wire \core_1.execute.rf.reg_outputs[6][15] ;
 wire \core_1.execute.rf.reg_outputs[6][1] ;
 wire \core_1.execute.rf.reg_outputs[6][2] ;
 wire \core_1.execute.rf.reg_outputs[6][3] ;
 wire \core_1.execute.rf.reg_outputs[6][4] ;
 wire \core_1.execute.rf.reg_outputs[6][5] ;
 wire \core_1.execute.rf.reg_outputs[6][6] ;
 wire \core_1.execute.rf.reg_outputs[6][7] ;
 wire \core_1.execute.rf.reg_outputs[6][8] ;
 wire \core_1.execute.rf.reg_outputs[6][9] ;
 wire \core_1.execute.rf.reg_outputs[7][0] ;
 wire \core_1.execute.rf.reg_outputs[7][10] ;
 wire \core_1.execute.rf.reg_outputs[7][11] ;
 wire \core_1.execute.rf.reg_outputs[7][12] ;
 wire \core_1.execute.rf.reg_outputs[7][13] ;
 wire \core_1.execute.rf.reg_outputs[7][14] ;
 wire \core_1.execute.rf.reg_outputs[7][15] ;
 wire \core_1.execute.rf.reg_outputs[7][1] ;
 wire \core_1.execute.rf.reg_outputs[7][2] ;
 wire \core_1.execute.rf.reg_outputs[7][3] ;
 wire \core_1.execute.rf.reg_outputs[7][4] ;
 wire \core_1.execute.rf.reg_outputs[7][5] ;
 wire \core_1.execute.rf.reg_outputs[7][6] ;
 wire \core_1.execute.rf.reg_outputs[7][7] ;
 wire \core_1.execute.rf.reg_outputs[7][8] ;
 wire \core_1.execute.rf.reg_outputs[7][9] ;
 wire \core_1.execute.sreg_data_page ;
 wire \core_1.execute.sreg_irq_flags.i_d[2] ;
 wire \core_1.execute.sreg_irq_flags.o_d[0] ;
 wire \core_1.execute.sreg_irq_flags.o_d[1] ;
 wire \core_1.execute.sreg_irq_flags.o_d[2] ;
 wire \core_1.execute.sreg_irq_flags.o_d[3] ;
 wire \core_1.execute.sreg_irq_flags.o_d[4] ;
 wire \core_1.execute.sreg_irq_pc.o_d[0] ;
 wire \core_1.execute.sreg_irq_pc.o_d[10] ;
 wire \core_1.execute.sreg_irq_pc.o_d[11] ;
 wire \core_1.execute.sreg_irq_pc.o_d[12] ;
 wire \core_1.execute.sreg_irq_pc.o_d[13] ;
 wire \core_1.execute.sreg_irq_pc.o_d[14] ;
 wire \core_1.execute.sreg_irq_pc.o_d[15] ;
 wire \core_1.execute.sreg_irq_pc.o_d[1] ;
 wire \core_1.execute.sreg_irq_pc.o_d[2] ;
 wire \core_1.execute.sreg_irq_pc.o_d[3] ;
 wire \core_1.execute.sreg_irq_pc.o_d[4] ;
 wire \core_1.execute.sreg_irq_pc.o_d[5] ;
 wire \core_1.execute.sreg_irq_pc.o_d[6] ;
 wire \core_1.execute.sreg_irq_pc.o_d[7] ;
 wire \core_1.execute.sreg_irq_pc.o_d[8] ;
 wire \core_1.execute.sreg_irq_pc.o_d[9] ;
 wire \core_1.execute.sreg_jtr_buff.o_d[0] ;
 wire \core_1.execute.sreg_jtr_buff.o_d[1] ;
 wire \core_1.execute.sreg_jtr_buff.o_d[2] ;
 wire \core_1.execute.sreg_long_ptr_en ;
 wire \core_1.execute.sreg_priv_control.o_d[0] ;
 wire \core_1.execute.sreg_priv_control.o_d[10] ;
 wire \core_1.execute.sreg_priv_control.o_d[11] ;
 wire \core_1.execute.sreg_priv_control.o_d[12] ;
 wire \core_1.execute.sreg_priv_control.o_d[13] ;
 wire \core_1.execute.sreg_priv_control.o_d[14] ;
 wire \core_1.execute.sreg_priv_control.o_d[15] ;
 wire \core_1.execute.sreg_priv_control.o_d[4] ;
 wire \core_1.execute.sreg_priv_control.o_d[5] ;
 wire \core_1.execute.sreg_priv_control.o_d[6] ;
 wire \core_1.execute.sreg_priv_control.o_d[7] ;
 wire \core_1.execute.sreg_priv_control.o_d[8] ;
 wire \core_1.execute.sreg_priv_control.o_d[9] ;
 wire \core_1.execute.sreg_scratch.o_d[0] ;
 wire \core_1.execute.sreg_scratch.o_d[10] ;
 wire \core_1.execute.sreg_scratch.o_d[11] ;
 wire \core_1.execute.sreg_scratch.o_d[12] ;
 wire \core_1.execute.sreg_scratch.o_d[13] ;
 wire \core_1.execute.sreg_scratch.o_d[14] ;
 wire \core_1.execute.sreg_scratch.o_d[15] ;
 wire \core_1.execute.sreg_scratch.o_d[1] ;
 wire \core_1.execute.sreg_scratch.o_d[2] ;
 wire \core_1.execute.sreg_scratch.o_d[3] ;
 wire \core_1.execute.sreg_scratch.o_d[4] ;
 wire \core_1.execute.sreg_scratch.o_d[5] ;
 wire \core_1.execute.sreg_scratch.o_d[6] ;
 wire \core_1.execute.sreg_scratch.o_d[7] ;
 wire \core_1.execute.sreg_scratch.o_d[8] ;
 wire \core_1.execute.sreg_scratch.o_d[9] ;
 wire \core_1.execute.trap_flag ;
 wire \core_1.fetch.current_req_branch_pred ;
 wire \core_1.fetch.dbg_out ;
 wire \core_1.fetch.flush_event_invalidate ;
 wire \core_1.fetch.out_buffer_data_instr[0] ;
 wire \core_1.fetch.out_buffer_data_instr[10] ;
 wire \core_1.fetch.out_buffer_data_instr[11] ;
 wire \core_1.fetch.out_buffer_data_instr[12] ;
 wire \core_1.fetch.out_buffer_data_instr[13] ;
 wire \core_1.fetch.out_buffer_data_instr[14] ;
 wire \core_1.fetch.out_buffer_data_instr[15] ;
 wire \core_1.fetch.out_buffer_data_instr[16] ;
 wire \core_1.fetch.out_buffer_data_instr[17] ;
 wire \core_1.fetch.out_buffer_data_instr[18] ;
 wire \core_1.fetch.out_buffer_data_instr[19] ;
 wire \core_1.fetch.out_buffer_data_instr[1] ;
 wire \core_1.fetch.out_buffer_data_instr[20] ;
 wire \core_1.fetch.out_buffer_data_instr[21] ;
 wire \core_1.fetch.out_buffer_data_instr[22] ;
 wire \core_1.fetch.out_buffer_data_instr[23] ;
 wire \core_1.fetch.out_buffer_data_instr[24] ;
 wire \core_1.fetch.out_buffer_data_instr[25] ;
 wire \core_1.fetch.out_buffer_data_instr[26] ;
 wire \core_1.fetch.out_buffer_data_instr[27] ;
 wire \core_1.fetch.out_buffer_data_instr[28] ;
 wire \core_1.fetch.out_buffer_data_instr[29] ;
 wire \core_1.fetch.out_buffer_data_instr[2] ;
 wire \core_1.fetch.out_buffer_data_instr[30] ;
 wire \core_1.fetch.out_buffer_data_instr[31] ;
 wire \core_1.fetch.out_buffer_data_instr[3] ;
 wire \core_1.fetch.out_buffer_data_instr[4] ;
 wire \core_1.fetch.out_buffer_data_instr[5] ;
 wire \core_1.fetch.out_buffer_data_instr[6] ;
 wire \core_1.fetch.out_buffer_data_instr[7] ;
 wire \core_1.fetch.out_buffer_data_instr[8] ;
 wire \core_1.fetch.out_buffer_data_instr[9] ;
 wire \core_1.fetch.out_buffer_data_pred ;
 wire \core_1.fetch.out_buffer_valid ;
 wire \core_1.fetch.pc_flush_override ;
 wire \core_1.fetch.pc_reset_override ;
 wire \core_1.fetch.prev_req_branch_pred ;
 wire \core_1.fetch.prev_request_pc[0] ;
 wire \core_1.fetch.prev_request_pc[10] ;
 wire \core_1.fetch.prev_request_pc[11] ;
 wire \core_1.fetch.prev_request_pc[12] ;
 wire \core_1.fetch.prev_request_pc[13] ;
 wire \core_1.fetch.prev_request_pc[14] ;
 wire \core_1.fetch.prev_request_pc[15] ;
 wire \core_1.fetch.prev_request_pc[1] ;
 wire \core_1.fetch.prev_request_pc[2] ;
 wire \core_1.fetch.prev_request_pc[3] ;
 wire \core_1.fetch.prev_request_pc[4] ;
 wire \core_1.fetch.prev_request_pc[5] ;
 wire \core_1.fetch.prev_request_pc[6] ;
 wire \core_1.fetch.prev_request_pc[7] ;
 wire \core_1.fetch.prev_request_pc[8] ;
 wire \core_1.fetch.prev_request_pc[9] ;
 wire \core_1.fetch.submitable ;
 wire net213;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net214;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net215;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire clknet_leaf_0_i_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire clknet_leaf_1_i_clk;
 wire clknet_leaf_2_i_clk;
 wire clknet_leaf_3_i_clk;
 wire clknet_leaf_4_i_clk;
 wire clknet_leaf_5_i_clk;
 wire clknet_leaf_6_i_clk;
 wire clknet_leaf_7_i_clk;
 wire clknet_leaf_8_i_clk;
 wire clknet_leaf_9_i_clk;
 wire clknet_leaf_10_i_clk;
 wire clknet_leaf_11_i_clk;
 wire clknet_leaf_12_i_clk;
 wire clknet_leaf_13_i_clk;
 wire clknet_leaf_14_i_clk;
 wire clknet_leaf_15_i_clk;
 wire clknet_leaf_16_i_clk;
 wire clknet_leaf_17_i_clk;
 wire clknet_leaf_18_i_clk;
 wire clknet_leaf_19_i_clk;
 wire clknet_leaf_20_i_clk;
 wire clknet_leaf_21_i_clk;
 wire clknet_leaf_22_i_clk;
 wire clknet_leaf_23_i_clk;
 wire clknet_leaf_24_i_clk;
 wire clknet_leaf_25_i_clk;
 wire clknet_leaf_26_i_clk;
 wire clknet_leaf_27_i_clk;
 wire clknet_leaf_28_i_clk;
 wire clknet_leaf_29_i_clk;
 wire clknet_leaf_30_i_clk;
 wire clknet_leaf_31_i_clk;
 wire clknet_leaf_32_i_clk;
 wire clknet_leaf_33_i_clk;
 wire clknet_leaf_34_i_clk;
 wire clknet_leaf_35_i_clk;
 wire clknet_leaf_36_i_clk;
 wire clknet_leaf_37_i_clk;
 wire clknet_leaf_38_i_clk;
 wire clknet_leaf_39_i_clk;
 wire clknet_leaf_40_i_clk;
 wire clknet_leaf_41_i_clk;
 wire clknet_leaf_42_i_clk;
 wire clknet_leaf_43_i_clk;
 wire clknet_0_i_clk;
 wire clknet_1_0_0_i_clk;
 wire clknet_1_0_1_i_clk;
 wire clknet_1_1_0_i_clk;
 wire clknet_1_1_1_i_clk;
 wire clknet_2_0_0_i_clk;
 wire clknet_2_1_0_i_clk;
 wire clknet_2_2_0_i_clk;
 wire clknet_2_3_0_i_clk;

 sky130_fd_sc_hd__or3_1 _3331_ (.A(\core_1.dec_r_reg_sel[2] ),
    .B(\core_1.dec_r_reg_sel[0] ),
    .C(\core_1.dec_r_reg_sel[1] ),
    .X(_0515_));
 sky130_fd_sc_hd__buf_4 _3332_ (.A(_0515_),
    .X(_0516_));
 sky130_fd_sc_hd__buf_8 _3333_ (.A(_0516_),
    .X(_0517_));
 sky130_fd_sc_hd__and3b_1 _3334_ (.A_N(\core_1.dec_r_reg_sel[0] ),
    .B(\core_1.dec_r_reg_sel[1] ),
    .C(\core_1.dec_r_reg_sel[2] ),
    .X(_0518_));
 sky130_fd_sc_hd__clkbuf_4 _3335_ (.A(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__clkbuf_2 _3336_ (.A(\core_1.dec_r_reg_sel[2] ),
    .X(_0520_));
 sky130_fd_sc_hd__buf_2 _3337_ (.A(\core_1.dec_r_reg_sel[0] ),
    .X(_0521_));
 sky130_fd_sc_hd__clkbuf_2 _3338_ (.A(_0521_),
    .X(_0522_));
 sky130_fd_sc_hd__buf_2 _3339_ (.A(\core_1.dec_r_reg_sel[1] ),
    .X(_0523_));
 sky130_fd_sc_hd__clkbuf_2 _3340_ (.A(_0523_),
    .X(_0524_));
 sky130_fd_sc_hd__and3_1 _3341_ (.A(_0520_),
    .B(_0522_),
    .C(_0524_),
    .X(_0525_));
 sky130_fd_sc_hd__and3b_1 _3342_ (.A_N(\core_1.dec_r_reg_sel[1] ),
    .B(\core_1.dec_r_reg_sel[0] ),
    .C(\core_1.dec_r_reg_sel[2] ),
    .X(_0526_));
 sky130_fd_sc_hd__buf_4 _3343_ (.A(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__a22o_1 _3344_ (.A1(\core_1.execute.rf.reg_outputs[7][15] ),
    .A2(_0525_),
    .B1(_0527_),
    .B2(\core_1.execute.rf.reg_outputs[5][15] ),
    .X(_0528_));
 sky130_fd_sc_hd__a21o_1 _3345_ (.A1(\core_1.execute.rf.reg_outputs[6][15] ),
    .A2(_0519_),
    .B1(_0528_),
    .X(_0529_));
 sky130_fd_sc_hd__clkbuf_2 _3346_ (.A(\core_1.dec_r_reg_sel[2] ),
    .X(_0530_));
 sky130_fd_sc_hd__nor3b_2 _3347_ (.A(_0530_),
    .B(_0523_),
    .C_N(_0521_),
    .Y(_0531_));
 sky130_fd_sc_hd__buf_4 _3348_ (.A(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__buf_2 _3349_ (.A(\core_1.dec_r_reg_sel[2] ),
    .X(_0533_));
 sky130_fd_sc_hd__buf_2 _3350_ (.A(_0533_),
    .X(_0534_));
 sky130_fd_sc_hd__inv_2 _3351_ (.A(_0534_),
    .Y(_0535_));
 sky130_fd_sc_hd__buf_2 _3352_ (.A(\core_1.dec_r_reg_sel[0] ),
    .X(_0536_));
 sky130_fd_sc_hd__buf_2 _3353_ (.A(\core_1.dec_r_reg_sel[1] ),
    .X(_0537_));
 sky130_fd_sc_hd__nor2_2 _3354_ (.A(_0536_),
    .B(_0537_),
    .Y(_0538_));
 sky130_fd_sc_hd__o21a_1 _3355_ (.A1(\core_1.execute.rf.reg_outputs[4][15] ),
    .A2(_0535_),
    .B1(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__nor3b_2 _3356_ (.A(\core_1.dec_r_reg_sel[2] ),
    .B(\core_1.dec_r_reg_sel[0] ),
    .C_N(\core_1.dec_r_reg_sel[1] ),
    .Y(_0540_));
 sky130_fd_sc_hd__buf_4 _3357_ (.A(_0540_),
    .X(_0541_));
 sky130_fd_sc_hd__and3b_2 _3358_ (.A_N(_0530_),
    .B(_0536_),
    .C(_0537_),
    .X(_0542_));
 sky130_fd_sc_hd__a22o_1 _3359_ (.A1(\core_1.execute.rf.reg_outputs[2][15] ),
    .A2(_0541_),
    .B1(_0542_),
    .B2(\core_1.execute.rf.reg_outputs[3][15] ),
    .X(_0543_));
 sky130_fd_sc_hd__a211o_1 _3360_ (.A1(\core_1.execute.rf.reg_outputs[1][15] ),
    .A2(_0532_),
    .B1(_0539_),
    .C1(_0543_),
    .X(_0544_));
 sky130_fd_sc_hd__o22ai_4 _3361_ (.A1(net94),
    .A2(_0517_),
    .B1(_0529_),
    .B2(_0544_),
    .Y(_0545_));
 sky130_fd_sc_hd__clkinv_4 _3362_ (.A(_0545_),
    .Y(net200));
 sky130_fd_sc_hd__a22o_1 _3363_ (.A1(\core_1.execute.rf.reg_outputs[6][14] ),
    .A2(_0519_),
    .B1(_0525_),
    .B2(\core_1.execute.rf.reg_outputs[7][14] ),
    .X(_0546_));
 sky130_fd_sc_hd__a21oi_1 _3364_ (.A1(\core_1.execute.rf.reg_outputs[5][14] ),
    .A2(_0527_),
    .B1(_0546_),
    .Y(_0547_));
 sky130_fd_sc_hd__buf_2 _3365_ (.A(_0533_),
    .X(_0548_));
 sky130_fd_sc_hd__or2b_1 _3366_ (.A(\core_1.execute.rf.reg_outputs[4][14] ),
    .B_N(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__a22o_1 _3367_ (.A1(\core_1.execute.rf.reg_outputs[3][14] ),
    .A2(_0542_),
    .B1(_0549_),
    .B2(_0538_),
    .X(_0550_));
 sky130_fd_sc_hd__a221oi_2 _3368_ (.A1(\core_1.execute.rf.reg_outputs[2][14] ),
    .A2(_0541_),
    .B1(_0532_),
    .B2(\core_1.execute.rf.reg_outputs[1][14] ),
    .C1(_0550_),
    .Y(_0551_));
 sky130_fd_sc_hd__nor2_1 _3369_ (.A(net93),
    .B(_0517_),
    .Y(_0552_));
 sky130_fd_sc_hd__a21o_4 _3370_ (.A1(_0547_),
    .A2(_0551_),
    .B1(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__clkinv_2 _3371_ (.A(_0553_),
    .Y(net199));
 sky130_fd_sc_hd__nor3b_4 _3372_ (.A(_0521_),
    .B(_0523_),
    .C_N(_0530_),
    .Y(_0554_));
 sky130_fd_sc_hd__buf_2 _3373_ (.A(_0524_),
    .X(_0555_));
 sky130_fd_sc_hd__buf_2 _3374_ (.A(_0536_),
    .X(_0556_));
 sky130_fd_sc_hd__and4bb_1 _3375_ (.A_N(_0548_),
    .B_N(_0555_),
    .C(_0556_),
    .D(\core_1.execute.rf.reg_outputs[1][13] ),
    .X(_0557_));
 sky130_fd_sc_hd__clkbuf_4 _3376_ (.A(_0522_),
    .X(_0558_));
 sky130_fd_sc_hd__and4b_1 _3377_ (.A_N(_0555_),
    .B(_0558_),
    .C(_0548_),
    .D(\core_1.execute.rf.reg_outputs[5][13] ),
    .X(_0559_));
 sky130_fd_sc_hd__and4b_1 _3378_ (.A_N(_0558_),
    .B(_0555_),
    .C(\core_1.execute.rf.reg_outputs[6][13] ),
    .D(_0534_),
    .X(_0560_));
 sky130_fd_sc_hd__a2111o_1 _3379_ (.A1(\core_1.execute.rf.reg_outputs[4][13] ),
    .A2(_0554_),
    .B1(_0557_),
    .C1(_0559_),
    .D1(_0560_),
    .X(_0561_));
 sky130_fd_sc_hd__buf_2 _3380_ (.A(_0523_),
    .X(_0562_));
 sky130_fd_sc_hd__and4b_1 _3381_ (.A_N(_0534_),
    .B(_0558_),
    .C(_0562_),
    .D(\core_1.execute.rf.reg_outputs[3][13] ),
    .X(_0563_));
 sky130_fd_sc_hd__and4_1 _3382_ (.A(\core_1.execute.rf.reg_outputs[7][13] ),
    .B(_0534_),
    .C(_0558_),
    .D(_0555_),
    .X(_0564_));
 sky130_fd_sc_hd__nor3_1 _3383_ (.A(\core_1.dec_r_reg_sel[2] ),
    .B(_0521_),
    .C(_0523_),
    .Y(_0565_));
 sky130_fd_sc_hd__buf_4 _3384_ (.A(_0565_),
    .X(_0566_));
 sky130_fd_sc_hd__a2111o_1 _3385_ (.A1(\core_1.execute.rf.reg_outputs[2][13] ),
    .A2(_0541_),
    .B1(_0563_),
    .C1(_0564_),
    .D1(_0566_),
    .X(_0567_));
 sky130_fd_sc_hd__o22ai_4 _3386_ (.A1(net92),
    .A2(_0517_),
    .B1(_0561_),
    .B2(_0567_),
    .Y(_0568_));
 sky130_fd_sc_hd__clkinv_4 _3387_ (.A(_0568_),
    .Y(net198));
 sky130_fd_sc_hd__a22o_1 _3388_ (.A1(\core_1.execute.rf.reg_outputs[5][12] ),
    .A2(_0527_),
    .B1(_0554_),
    .B2(\core_1.execute.rf.reg_outputs[4][12] ),
    .X(_0569_));
 sky130_fd_sc_hd__a22o_1 _3389_ (.A1(\core_1.execute.rf.reg_outputs[6][12] ),
    .A2(_0519_),
    .B1(_0532_),
    .B2(\core_1.execute.rf.reg_outputs[1][12] ),
    .X(_0570_));
 sky130_fd_sc_hd__and4b_1 _3390_ (.A_N(_0534_),
    .B(_0558_),
    .C(_0555_),
    .D(\core_1.execute.rf.reg_outputs[3][12] ),
    .X(_0571_));
 sky130_fd_sc_hd__and4_1 _3391_ (.A(\core_1.execute.rf.reg_outputs[7][12] ),
    .B(_0534_),
    .C(_0558_),
    .D(_0555_),
    .X(_0572_));
 sky130_fd_sc_hd__a2111o_1 _3392_ (.A1(\core_1.execute.rf.reg_outputs[2][12] ),
    .A2(_0541_),
    .B1(_0571_),
    .C1(_0572_),
    .D1(_0566_),
    .X(_0573_));
 sky130_fd_sc_hd__or2_1 _3393_ (.A(net91),
    .B(_0517_),
    .X(_0574_));
 sky130_fd_sc_hd__o31ai_4 _3394_ (.A1(_0569_),
    .A2(_0570_),
    .A3(_0573_),
    .B1(_0574_),
    .Y(_0575_));
 sky130_fd_sc_hd__inv_2 _3395_ (.A(_0575_),
    .Y(net197));
 sky130_fd_sc_hd__a22o_1 _3396_ (.A1(\core_1.execute.rf.reg_outputs[5][11] ),
    .A2(_0527_),
    .B1(_0554_),
    .B2(\core_1.execute.rf.reg_outputs[4][11] ),
    .X(_0576_));
 sky130_fd_sc_hd__a22o_1 _3397_ (.A1(\core_1.execute.rf.reg_outputs[6][11] ),
    .A2(_0519_),
    .B1(_0531_),
    .B2(\core_1.execute.rf.reg_outputs[1][11] ),
    .X(_0577_));
 sky130_fd_sc_hd__and4b_1 _3398_ (.A_N(_0530_),
    .B(_0521_),
    .C(_0523_),
    .D(\core_1.execute.rf.reg_outputs[3][11] ),
    .X(_0578_));
 sky130_fd_sc_hd__and4_1 _3399_ (.A(\core_1.execute.rf.reg_outputs[7][11] ),
    .B(_0530_),
    .C(_0521_),
    .D(_0523_),
    .X(_0579_));
 sky130_fd_sc_hd__a2111o_1 _3400_ (.A1(\core_1.execute.rf.reg_outputs[2][11] ),
    .A2(_0540_),
    .B1(_0578_),
    .C1(_0579_),
    .D1(_0565_),
    .X(_0580_));
 sky130_fd_sc_hd__or2_1 _3401_ (.A(net90),
    .B(_0516_),
    .X(_0581_));
 sky130_fd_sc_hd__o31ai_4 _3402_ (.A1(_0576_),
    .A2(_0577_),
    .A3(_0580_),
    .B1(_0581_),
    .Y(_0582_));
 sky130_fd_sc_hd__clkinv_2 _3403_ (.A(_0582_),
    .Y(net196));
 sky130_fd_sc_hd__a22o_1 _3404_ (.A1(\core_1.execute.rf.reg_outputs[5][10] ),
    .A2(_0526_),
    .B1(_0554_),
    .B2(\core_1.execute.rf.reg_outputs[4][10] ),
    .X(_0583_));
 sky130_fd_sc_hd__a22o_1 _3405_ (.A1(\core_1.execute.rf.reg_outputs[6][10] ),
    .A2(_0518_),
    .B1(_0531_),
    .B2(\core_1.execute.rf.reg_outputs[1][10] ),
    .X(_0584_));
 sky130_fd_sc_hd__and4b_1 _3406_ (.A_N(_0530_),
    .B(_0521_),
    .C(_0523_),
    .D(\core_1.execute.rf.reg_outputs[3][10] ),
    .X(_0585_));
 sky130_fd_sc_hd__and4_1 _3407_ (.A(\core_1.execute.rf.reg_outputs[7][10] ),
    .B(_0530_),
    .C(_0521_),
    .D(_0523_),
    .X(_0586_));
 sky130_fd_sc_hd__a2111o_1 _3408_ (.A1(\core_1.execute.rf.reg_outputs[2][10] ),
    .A2(_0540_),
    .B1(_0585_),
    .C1(_0586_),
    .D1(_0565_),
    .X(_0587_));
 sky130_fd_sc_hd__o32ai_4 _3409_ (.A1(_0583_),
    .A2(_0584_),
    .A3(_0587_),
    .B1(_0516_),
    .B2(net89),
    .Y(_0588_));
 sky130_fd_sc_hd__inv_2 _3410_ (.A(_0588_),
    .Y(net195));
 sky130_fd_sc_hd__and4b_1 _3411_ (.A_N(_0537_),
    .B(_0536_),
    .C(_0530_),
    .D(\core_1.execute.rf.reg_outputs[5][9] ),
    .X(_0589_));
 sky130_fd_sc_hd__and4b_1 _3412_ (.A_N(_0536_),
    .B(_0537_),
    .C(\core_1.execute.rf.reg_outputs[6][9] ),
    .D(_0533_),
    .X(_0590_));
 sky130_fd_sc_hd__and4bb_1 _3413_ (.A_N(_0533_),
    .B_N(_0537_),
    .C(_0536_),
    .D(\core_1.execute.rf.reg_outputs[1][9] ),
    .X(_0591_));
 sky130_fd_sc_hd__a2111o_1 _3414_ (.A1(\core_1.execute.rf.reg_outputs[4][9] ),
    .A2(_0554_),
    .B1(_0589_),
    .C1(_0590_),
    .D1(_0591_),
    .X(_0592_));
 sky130_fd_sc_hd__and4b_1 _3415_ (.A_N(_0533_),
    .B(_0536_),
    .C(_0537_),
    .D(\core_1.execute.rf.reg_outputs[3][9] ),
    .X(_0593_));
 sky130_fd_sc_hd__and4_1 _3416_ (.A(\core_1.execute.rf.reg_outputs[7][9] ),
    .B(_0533_),
    .C(_0536_),
    .D(_0537_),
    .X(_0594_));
 sky130_fd_sc_hd__a2111o_1 _3417_ (.A1(\core_1.execute.rf.reg_outputs[2][9] ),
    .A2(_0541_),
    .B1(_0593_),
    .C1(_0594_),
    .D1(_0566_),
    .X(_0595_));
 sky130_fd_sc_hd__o22ai_4 _3418_ (.A1(net103),
    .A2(_0516_),
    .B1(_0592_),
    .B2(_0595_),
    .Y(_0596_));
 sky130_fd_sc_hd__inv_2 _3419_ (.A(_0596_),
    .Y(net209));
 sky130_fd_sc_hd__a22o_1 _3420_ (.A1(\core_1.execute.rf.reg_outputs[5][8] ),
    .A2(_0527_),
    .B1(_0554_),
    .B2(\core_1.execute.rf.reg_outputs[4][8] ),
    .X(_0597_));
 sky130_fd_sc_hd__a22o_1 _3421_ (.A1(\core_1.execute.rf.reg_outputs[6][8] ),
    .A2(_0519_),
    .B1(_0531_),
    .B2(\core_1.execute.rf.reg_outputs[1][8] ),
    .X(_0598_));
 sky130_fd_sc_hd__and4b_1 _3422_ (.A_N(_0530_),
    .B(_0521_),
    .C(_0523_),
    .D(\core_1.execute.rf.reg_outputs[3][8] ),
    .X(_0599_));
 sky130_fd_sc_hd__and4_1 _3423_ (.A(\core_1.execute.rf.reg_outputs[7][8] ),
    .B(_0530_),
    .C(_0521_),
    .D(_0537_),
    .X(_0600_));
 sky130_fd_sc_hd__a2111o_1 _3424_ (.A1(\core_1.execute.rf.reg_outputs[2][8] ),
    .A2(_0540_),
    .B1(_0599_),
    .C1(_0600_),
    .D1(_0566_),
    .X(_0601_));
 sky130_fd_sc_hd__or2_1 _3425_ (.A(net102),
    .B(_0516_),
    .X(_0602_));
 sky130_fd_sc_hd__o31ai_4 _3426_ (.A1(_0597_),
    .A2(_0598_),
    .A3(_0601_),
    .B1(_0602_),
    .Y(_0603_));
 sky130_fd_sc_hd__inv_2 _3427_ (.A(_0603_),
    .Y(net208));
 sky130_fd_sc_hd__and4b_1 _3428_ (.A_N(_0522_),
    .B(_0524_),
    .C(\core_1.execute.rf.reg_outputs[6][7] ),
    .D(_0533_),
    .X(_0604_));
 sky130_fd_sc_hd__and4b_1 _3429_ (.A_N(_0524_),
    .B(_0522_),
    .C(_0520_),
    .D(\core_1.execute.rf.reg_outputs[5][7] ),
    .X(_0605_));
 sky130_fd_sc_hd__and4bb_1 _3430_ (.A_N(_0520_),
    .B_N(_0524_),
    .C(_0522_),
    .D(\core_1.execute.rf.reg_outputs[1][7] ),
    .X(_0606_));
 sky130_fd_sc_hd__a2111oi_1 _3431_ (.A1(\core_1.execute.rf.reg_outputs[4][7] ),
    .A2(_0554_),
    .B1(_0604_),
    .C1(_0605_),
    .D1(_0606_),
    .Y(_0607_));
 sky130_fd_sc_hd__and4b_1 _3432_ (.A_N(_0520_),
    .B(_0522_),
    .C(_0524_),
    .D(\core_1.execute.rf.reg_outputs[3][7] ),
    .X(_0608_));
 sky130_fd_sc_hd__and4_1 _3433_ (.A(\core_1.execute.rf.reg_outputs[7][7] ),
    .B(_0520_),
    .C(_0522_),
    .D(_0524_),
    .X(_0609_));
 sky130_fd_sc_hd__a2111oi_1 _3434_ (.A1(\core_1.execute.rf.reg_outputs[2][7] ),
    .A2(_0541_),
    .B1(_0608_),
    .C1(_0609_),
    .D1(_0566_),
    .Y(_0610_));
 sky130_fd_sc_hd__a2bb2o_4 _3435_ (.A1_N(net101),
    .A2_N(_0516_),
    .B1(_0607_),
    .B2(_0610_),
    .X(_0611_));
 sky130_fd_sc_hd__clkinv_4 _3436_ (.A(_0611_),
    .Y(net207));
 sky130_fd_sc_hd__and4_1 _3437_ (.A(\core_1.execute.rf.reg_outputs[7][6] ),
    .B(_0533_),
    .C(_0536_),
    .D(_0537_),
    .X(_0612_));
 sky130_fd_sc_hd__a221o_1 _3438_ (.A1(\core_1.execute.rf.reg_outputs[2][6] ),
    .A2(_0540_),
    .B1(_0542_),
    .B2(\core_1.execute.rf.reg_outputs[3][6] ),
    .C1(_0612_),
    .X(_0613_));
 sky130_fd_sc_hd__a22o_1 _3439_ (.A1(\core_1.execute.rf.reg_outputs[5][6] ),
    .A2(_0527_),
    .B1(_0532_),
    .B2(\core_1.execute.rf.reg_outputs[1][6] ),
    .X(_0614_));
 sky130_fd_sc_hd__a221o_1 _3440_ (.A1(\core_1.execute.rf.reg_outputs[4][6] ),
    .A2(_0538_),
    .B1(_0519_),
    .B2(\core_1.execute.rf.reg_outputs[6][6] ),
    .C1(_0566_),
    .X(_0615_));
 sky130_fd_sc_hd__or2_1 _3441_ (.A(net100),
    .B(_0516_),
    .X(_0616_));
 sky130_fd_sc_hd__o31ai_4 _3442_ (.A1(_0613_),
    .A2(_0614_),
    .A3(_0615_),
    .B1(_0616_),
    .Y(_0617_));
 sky130_fd_sc_hd__clkinv_4 _3443_ (.A(_0617_),
    .Y(net206));
 sky130_fd_sc_hd__a221o_1 _3444_ (.A1(\core_1.execute.rf.reg_outputs[4][5] ),
    .A2(_0538_),
    .B1(_0541_),
    .B2(\core_1.execute.rf.reg_outputs[2][5] ),
    .C1(_0566_),
    .X(_0618_));
 sky130_fd_sc_hd__a22o_1 _3445_ (.A1(\core_1.execute.rf.reg_outputs[5][5] ),
    .A2(_0527_),
    .B1(_0532_),
    .B2(\core_1.execute.rf.reg_outputs[1][5] ),
    .X(_0619_));
 sky130_fd_sc_hd__and4_1 _3446_ (.A(\core_1.execute.rf.reg_outputs[7][5] ),
    .B(_0548_),
    .C(_0556_),
    .D(_0562_),
    .X(_0620_));
 sky130_fd_sc_hd__a221o_1 _3447_ (.A1(\core_1.execute.rf.reg_outputs[6][5] ),
    .A2(_0519_),
    .B1(_0542_),
    .B2(\core_1.execute.rf.reg_outputs[3][5] ),
    .C1(_0620_),
    .X(_0621_));
 sky130_fd_sc_hd__or2_1 _3448_ (.A(net99),
    .B(_0516_),
    .X(_0622_));
 sky130_fd_sc_hd__o31ai_4 _3449_ (.A1(_0618_),
    .A2(_0619_),
    .A3(_0621_),
    .B1(_0622_),
    .Y(_0623_));
 sky130_fd_sc_hd__inv_2 _3450_ (.A(_0623_),
    .Y(net205));
 sky130_fd_sc_hd__a22o_1 _3451_ (.A1(\core_1.execute.rf.reg_outputs[5][4] ),
    .A2(_0527_),
    .B1(_0554_),
    .B2(\core_1.execute.rf.reg_outputs[4][4] ),
    .X(_0624_));
 sky130_fd_sc_hd__a22o_1 _3452_ (.A1(\core_1.execute.rf.reg_outputs[6][4] ),
    .A2(_0519_),
    .B1(_0532_),
    .B2(\core_1.execute.rf.reg_outputs[1][4] ),
    .X(_0625_));
 sky130_fd_sc_hd__and4b_1 _3453_ (.A_N(_0548_),
    .B(_0556_),
    .C(_0562_),
    .D(\core_1.execute.rf.reg_outputs[3][4] ),
    .X(_0626_));
 sky130_fd_sc_hd__and4_1 _3454_ (.A(\core_1.execute.rf.reg_outputs[7][4] ),
    .B(_0520_),
    .C(_0556_),
    .D(_0562_),
    .X(_0627_));
 sky130_fd_sc_hd__a2111o_1 _3455_ (.A1(\core_1.execute.rf.reg_outputs[2][4] ),
    .A2(_0541_),
    .B1(_0626_),
    .C1(_0627_),
    .D1(_0566_),
    .X(_0628_));
 sky130_fd_sc_hd__o32ai_4 _3456_ (.A1(_0624_),
    .A2(_0625_),
    .A3(_0628_),
    .B1(_0517_),
    .B2(net98),
    .Y(_0629_));
 sky130_fd_sc_hd__clkinv_4 _3457_ (.A(_0629_),
    .Y(net204));
 sky130_fd_sc_hd__a22o_1 _3458_ (.A1(\core_1.execute.rf.reg_outputs[5][3] ),
    .A2(_0527_),
    .B1(_0554_),
    .B2(\core_1.execute.rf.reg_outputs[4][3] ),
    .X(_0630_));
 sky130_fd_sc_hd__a22o_1 _3459_ (.A1(\core_1.execute.rf.reg_outputs[6][3] ),
    .A2(_0519_),
    .B1(_0532_),
    .B2(\core_1.execute.rf.reg_outputs[1][3] ),
    .X(_0631_));
 sky130_fd_sc_hd__and4b_1 _3460_ (.A_N(_0534_),
    .B(_0556_),
    .C(_0562_),
    .D(\core_1.execute.rf.reg_outputs[3][3] ),
    .X(_0632_));
 sky130_fd_sc_hd__and4_1 _3461_ (.A(\core_1.execute.rf.reg_outputs[7][3] ),
    .B(_0534_),
    .C(_0558_),
    .D(_0555_),
    .X(_0633_));
 sky130_fd_sc_hd__a2111o_1 _3462_ (.A1(\core_1.execute.rf.reg_outputs[2][3] ),
    .A2(_0541_),
    .B1(_0632_),
    .C1(_0633_),
    .D1(_0566_),
    .X(_0634_));
 sky130_fd_sc_hd__o32ai_4 _3463_ (.A1(_0630_),
    .A2(_0631_),
    .A3(_0634_),
    .B1(_0517_),
    .B2(net97),
    .Y(_0635_));
 sky130_fd_sc_hd__inv_2 _3464_ (.A(_0635_),
    .Y(net203));
 sky130_fd_sc_hd__and2_1 _3465_ (.A(\core_1.execute.rf.reg_outputs[7][2] ),
    .B(_0525_),
    .X(_0636_));
 sky130_fd_sc_hd__a22o_1 _3466_ (.A1(\core_1.execute.rf.reg_outputs[3][2] ),
    .A2(_0542_),
    .B1(_0532_),
    .B2(\core_1.execute.rf.reg_outputs[1][2] ),
    .X(_0637_));
 sky130_fd_sc_hd__or2b_1 _3467_ (.A(\core_1.execute.rf.reg_outputs[4][2] ),
    .B_N(_0520_),
    .X(_0638_));
 sky130_fd_sc_hd__and4b_1 _3468_ (.A_N(_0522_),
    .B(_0537_),
    .C(\core_1.execute.rf.reg_outputs[6][2] ),
    .D(_0533_),
    .X(_0639_));
 sky130_fd_sc_hd__and4b_1 _3469_ (.A_N(_0524_),
    .B(_0536_),
    .C(_0533_),
    .D(\core_1.execute.rf.reg_outputs[5][2] ),
    .X(_0640_));
 sky130_fd_sc_hd__and4bb_1 _3470_ (.A_N(_0520_),
    .B_N(_0522_),
    .C(_0524_),
    .D(\core_1.execute.rf.reg_outputs[2][2] ),
    .X(_0641_));
 sky130_fd_sc_hd__a2111o_1 _3471_ (.A1(_0538_),
    .A2(_0638_),
    .B1(_0639_),
    .C1(_0640_),
    .D1(_0641_),
    .X(_0642_));
 sky130_fd_sc_hd__o32ai_4 _3472_ (.A1(_0636_),
    .A2(_0637_),
    .A3(_0642_),
    .B1(_0517_),
    .B2(net96),
    .Y(_0643_));
 sky130_fd_sc_hd__inv_2 _3473_ (.A(_0643_),
    .Y(net202));
 sky130_fd_sc_hd__a22oi_4 _3474_ (.A1(\core_1.execute.rf.reg_outputs[5][1] ),
    .A2(_0527_),
    .B1(_0554_),
    .B2(\core_1.execute.rf.reg_outputs[4][1] ),
    .Y(_0644_));
 sky130_fd_sc_hd__a22oi_2 _3475_ (.A1(\core_1.execute.rf.reg_outputs[3][1] ),
    .A2(_0542_),
    .B1(_0532_),
    .B2(\core_1.execute.rf.reg_outputs[1][1] ),
    .Y(_0645_));
 sky130_fd_sc_hd__and4_1 _3476_ (.A(\core_1.execute.rf.reg_outputs[7][1] ),
    .B(_0520_),
    .C(_0522_),
    .D(_0524_),
    .X(_0646_));
 sky130_fd_sc_hd__and4b_1 _3477_ (.A_N(_0556_),
    .B(_0562_),
    .C(\core_1.execute.rf.reg_outputs[6][1] ),
    .D(_0520_),
    .X(_0647_));
 sky130_fd_sc_hd__a2111oi_4 _3478_ (.A1(\core_1.execute.rf.reg_outputs[2][1] ),
    .A2(_0541_),
    .B1(_0646_),
    .C1(_0647_),
    .D1(_0566_),
    .Y(_0648_));
 sky130_fd_sc_hd__nor2_1 _3479_ (.A(net95),
    .B(_0516_),
    .Y(_0649_));
 sky130_fd_sc_hd__a31o_4 _3480_ (.A1(_0644_),
    .A2(_0645_),
    .A3(_0648_),
    .B1(_0649_),
    .X(_0650_));
 sky130_fd_sc_hd__inv_2 _3481_ (.A(_0650_),
    .Y(net201));
 sky130_fd_sc_hd__and4_1 _3482_ (.A(\core_1.execute.rf.reg_outputs[7][0] ),
    .B(_0548_),
    .C(_0556_),
    .D(_0562_),
    .X(_0651_));
 sky130_fd_sc_hd__a221o_4 _3483_ (.A1(\core_1.execute.rf.reg_outputs[6][0] ),
    .A2(_0519_),
    .B1(_0532_),
    .B2(\core_1.execute.rf.reg_outputs[1][0] ),
    .C1(_0651_),
    .X(_0652_));
 sky130_fd_sc_hd__or2b_1 _3484_ (.A(\core_1.execute.rf.reg_outputs[4][0] ),
    .B_N(_0548_),
    .X(_0653_));
 sky130_fd_sc_hd__and4bb_1 _3485_ (.A_N(_0548_),
    .B_N(_0556_),
    .C(_0562_),
    .D(\core_1.execute.rf.reg_outputs[2][0] ),
    .X(_0654_));
 sky130_fd_sc_hd__and4b_1 _3486_ (.A_N(_0548_),
    .B(_0556_),
    .C(_0562_),
    .D(\core_1.execute.rf.reg_outputs[3][0] ),
    .X(_0655_));
 sky130_fd_sc_hd__and4b_1 _3487_ (.A_N(_0562_),
    .B(_0556_),
    .C(_0548_),
    .D(\core_1.execute.rf.reg_outputs[5][0] ),
    .X(_0656_));
 sky130_fd_sc_hd__a2111o_4 _3488_ (.A1(_0538_),
    .A2(_0653_),
    .B1(_0654_),
    .C1(_0655_),
    .D1(_0656_),
    .X(_0657_));
 sky130_fd_sc_hd__o22ai_4 _3489_ (.A1(net88),
    .A2(_0517_),
    .B1(_0652_),
    .B2(_0657_),
    .Y(_0658_));
 sky130_fd_sc_hd__clkinv_4 _3490_ (.A(_0658_),
    .Y(net194));
 sky130_fd_sc_hd__buf_6 _3491_ (.A(net71),
    .X(_0659_));
 sky130_fd_sc_hd__inv_2 _3492_ (.A(\core_1.fetch.pc_flush_override ),
    .Y(_0660_));
 sky130_fd_sc_hd__buf_4 _3493_ (.A(\core_1.fetch.out_buffer_valid ),
    .X(_0661_));
 sky130_fd_sc_hd__buf_6 _3494_ (.A(_0661_),
    .X(_0662_));
 sky130_fd_sc_hd__buf_6 _3495_ (.A(_0662_),
    .X(_0663_));
 sky130_fd_sc_hd__buf_4 _3496_ (.A(_0663_),
    .X(_0664_));
 sky130_fd_sc_hd__o21a_1 _3497_ (.A1(net19),
    .A2(net18),
    .B1(\core_1.execute.irq_en ),
    .X(_0665_));
 sky130_fd_sc_hd__or3_1 _3498_ (.A(net37),
    .B(\core_1.execute.sreg_irq_flags.i_d[2] ),
    .C(_0665_),
    .X(_0666_));
 sky130_fd_sc_hd__or2_4 _3499_ (.A(\core_1.execute.prev_sys ),
    .B(_0666_),
    .X(_0667_));
 sky130_fd_sc_hd__clkinv_4 _3500_ (.A(_0667_),
    .Y(_0668_));
 sky130_fd_sc_hd__nand2_2 _3501_ (.A(\core_1.execute.pc_high_out[3] ),
    .B(net105),
    .Y(_0669_));
 sky130_fd_sc_hd__clkbuf_4 _3502_ (.A(net105),
    .X(_0670_));
 sky130_fd_sc_hd__nand2_2 _3503_ (.A(\core_1.execute.pc_high_out[6] ),
    .B(_0670_),
    .Y(_0671_));
 sky130_fd_sc_hd__nand2_2 _3504_ (.A(\core_1.execute.pc_high_out[2] ),
    .B(net105),
    .Y(_0672_));
 sky130_fd_sc_hd__o22a_1 _3505_ (.A1(\core_1.execute.prev_pc_high[6] ),
    .A2(_0671_),
    .B1(_0672_),
    .B2(\core_1.execute.prev_pc_high[2] ),
    .X(_0673_));
 sky130_fd_sc_hd__nand2_2 _3506_ (.A(\core_1.execute.pc_high_out[1] ),
    .B(_0670_),
    .Y(_0674_));
 sky130_fd_sc_hd__nand2_1 _3507_ (.A(\core_1.execute.pc_high_out[7] ),
    .B(net105),
    .Y(_0675_));
 sky130_fd_sc_hd__a22o_1 _3508_ (.A1(\core_1.execute.prev_pc_high[7] ),
    .A2(_0675_),
    .B1(_0672_),
    .B2(\core_1.execute.prev_pc_high[2] ),
    .X(_0676_));
 sky130_fd_sc_hd__nand2_2 _3509_ (.A(\core_1.execute.pc_high_out[5] ),
    .B(_0670_),
    .Y(_0677_));
 sky130_fd_sc_hd__xnor2_1 _3510_ (.A(\core_1.execute.prev_pc_high[5] ),
    .B(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__a2bb2o_1 _3511_ (.A1_N(\core_1.execute.prev_pc_high[7] ),
    .A2_N(_0675_),
    .B1(_0669_),
    .B2(\core_1.execute.prev_pc_high[3] ),
    .X(_0679_));
 sky130_fd_sc_hd__nand2_2 _3512_ (.A(\core_1.execute.pc_high_out[4] ),
    .B(_0670_),
    .Y(_0680_));
 sky130_fd_sc_hd__a2bb2o_1 _3513_ (.A1_N(\core_1.execute.prev_pc_high[4] ),
    .A2_N(_0680_),
    .B1(_0671_),
    .B2(\core_1.execute.prev_pc_high[6] ),
    .X(_0681_));
 sky130_fd_sc_hd__or4_1 _3514_ (.A(_0676_),
    .B(_0678_),
    .C(_0679_),
    .D(_0681_),
    .X(_0682_));
 sky130_fd_sc_hd__a2bb2o_1 _3515_ (.A1_N(\core_1.execute.prev_pc_high[1] ),
    .A2_N(_0674_),
    .B1(_0680_),
    .B2(\core_1.execute.prev_pc_high[4] ),
    .X(_0683_));
 sky130_fd_sc_hd__nand2_2 _3516_ (.A(\core_1.execute.pc_high_out[0] ),
    .B(_0670_),
    .Y(_0684_));
 sky130_fd_sc_hd__xnor2_1 _3517_ (.A(\core_1.execute.prev_pc_high[0] ),
    .B(_0684_),
    .Y(_0685_));
 sky130_fd_sc_hd__a2111oi_1 _3518_ (.A1(\core_1.execute.prev_pc_high[1] ),
    .A2(_0674_),
    .B1(_0682_),
    .C1(_0683_),
    .D1(_0685_),
    .Y(_0686_));
 sky130_fd_sc_hd__o211a_2 _3519_ (.A1(\core_1.execute.prev_pc_high[3] ),
    .A2(_0669_),
    .B1(_0673_),
    .C1(_0686_),
    .X(_0687_));
 sky130_fd_sc_hd__nand2_1 _3520_ (.A(_0668_),
    .B(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hd__nor2_1 _3521_ (.A(\core_1.execute.hold_valid ),
    .B(\core_1.decode.o_submit ),
    .Y(_0689_));
 sky130_fd_sc_hd__or3_1 _3522_ (.A(\core_1.decode.i_flush ),
    .B(_0688_),
    .C(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__inv_2 _3523_ (.A(\core_1.execute.next_ready_delayed ),
    .Y(_0691_));
 sky130_fd_sc_hd__inv_2 _3524_ (.A(\core_1.dec_l_reg_sel[2] ),
    .Y(_0692_));
 sky130_fd_sc_hd__buf_4 _3525_ (.A(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__buf_4 _3526_ (.A(\core_1.dec_l_reg_sel[0] ),
    .X(_0694_));
 sky130_fd_sc_hd__clkbuf_4 _3527_ (.A(\core_1.dec_l_reg_sel[1] ),
    .X(_0695_));
 sky130_fd_sc_hd__nand2_4 _3528_ (.A(_0694_),
    .B(_0695_),
    .Y(_0696_));
 sky130_fd_sc_hd__inv_2 _3529_ (.A(\core_1.ew_reg_ie[2] ),
    .Y(_0697_));
 sky130_fd_sc_hd__buf_4 _3530_ (.A(\core_1.dec_l_reg_sel[1] ),
    .X(_0698_));
 sky130_fd_sc_hd__nand2b_4 _3531_ (.A_N(_0698_),
    .B(\core_1.dec_l_reg_sel[0] ),
    .Y(_0699_));
 sky130_fd_sc_hd__nor2_8 _3532_ (.A(\core_1.dec_l_reg_sel[0] ),
    .B(_0698_),
    .Y(_0700_));
 sky130_fd_sc_hd__clkbuf_4 _3533_ (.A(_0694_),
    .X(_0701_));
 sky130_fd_sc_hd__o21a_1 _3534_ (.A1(_0701_),
    .A2(\core_1.ew_reg_ie[3] ),
    .B1(_0695_),
    .X(_0702_));
 sky130_fd_sc_hd__a21oi_1 _3535_ (.A1(\core_1.ew_reg_ie[1] ),
    .A2(_0700_),
    .B1(_0702_),
    .Y(_0703_));
 sky130_fd_sc_hd__o211ai_1 _3536_ (.A1(_0697_),
    .A2(_0699_),
    .B1(_0703_),
    .C1(_0693_),
    .Y(_0704_));
 sky130_fd_sc_hd__and2_1 _3537_ (.A(_0693_),
    .B(_0696_),
    .X(_0705_));
 sky130_fd_sc_hd__mux4_1 _3538_ (.A0(\core_1.ew_reg_ie[5] ),
    .A1(\core_1.ew_reg_ie[6] ),
    .A2(\core_1.ew_reg_ie[7] ),
    .A3(\core_1.ew_reg_ie[4] ),
    .S0(_0701_),
    .S1(_0695_),
    .X(_0706_));
 sky130_fd_sc_hd__and2_2 _3539_ (.A(\core_1.execute.sreg_long_ptr_en ),
    .B(\core_1.dec_mem_long ),
    .X(_0707_));
 sky130_fd_sc_hd__o21a_1 _3540_ (.A1(_0705_),
    .A2(_0706_),
    .B1(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__o211a_1 _3541_ (.A1(_0693_),
    .A2(_0696_),
    .B1(_0704_),
    .C1(_0708_),
    .X(_0709_));
 sky130_fd_sc_hd__or2_1 _3542_ (.A(_0701_),
    .B(_0695_),
    .X(_0710_));
 sky130_fd_sc_hd__or3b_1 _3543_ (.A(_0701_),
    .B(\core_1.ew_reg_ie[2] ),
    .C_N(_0695_),
    .X(_0711_));
 sky130_fd_sc_hd__o221a_1 _3544_ (.A1(\core_1.ew_reg_ie[1] ),
    .A2(_0699_),
    .B1(_0710_),
    .B2(\core_1.ew_reg_ie[0] ),
    .C1(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__o211a_1 _3545_ (.A1(\core_1.ew_reg_ie[3] ),
    .A2(_0696_),
    .B1(_0712_),
    .C1(_0693_),
    .X(_0713_));
 sky130_fd_sc_hd__or3b_1 _3546_ (.A(_0701_),
    .B(\core_1.ew_reg_ie[6] ),
    .C_N(_0695_),
    .X(_0714_));
 sky130_fd_sc_hd__o221a_1 _3547_ (.A1(\core_1.ew_reg_ie[5] ),
    .A2(_0699_),
    .B1(_0710_),
    .B2(\core_1.ew_reg_ie[4] ),
    .C1(_0714_),
    .X(_0715_));
 sky130_fd_sc_hd__clkbuf_4 _3548_ (.A(\core_1.dec_l_reg_sel[2] ),
    .X(_0716_));
 sky130_fd_sc_hd__buf_4 _3549_ (.A(_0716_),
    .X(_0717_));
 sky130_fd_sc_hd__o211a_1 _3550_ (.A1(\core_1.ew_reg_ie[7] ),
    .A2(_0696_),
    .B1(_0715_),
    .C1(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__o31a_1 _3551_ (.A1(_0709_),
    .A2(_0713_),
    .A3(_0718_),
    .B1(\core_1.dec_used_operands[0] ),
    .X(_0719_));
 sky130_fd_sc_hd__mux4_1 _3552_ (.A0(\core_1.ew_reg_ie[0] ),
    .A1(\core_1.ew_reg_ie[1] ),
    .A2(\core_1.ew_reg_ie[2] ),
    .A3(\core_1.ew_reg_ie[3] ),
    .S0(_0558_),
    .S1(_0555_),
    .X(_0720_));
 sky130_fd_sc_hd__mux4_1 _3553_ (.A0(\core_1.ew_reg_ie[4] ),
    .A1(\core_1.ew_reg_ie[5] ),
    .A2(\core_1.ew_reg_ie[6] ),
    .A3(\core_1.ew_reg_ie[7] ),
    .S0(_0558_),
    .S1(_0555_),
    .X(_0721_));
 sky130_fd_sc_hd__or2_1 _3554_ (.A(_0535_),
    .B(_0721_),
    .X(_0722_));
 sky130_fd_sc_hd__o211a_1 _3555_ (.A1(_0534_),
    .A2(_0720_),
    .B1(_0722_),
    .C1(\core_1.dec_used_operands[1] ),
    .X(_0723_));
 sky130_fd_sc_hd__o22a_2 _3556_ (.A1(\core_1.ew_submit ),
    .A2(_0691_),
    .B1(_0719_),
    .B2(_0723_),
    .X(_0724_));
 sky130_fd_sc_hd__inv_2 _3557_ (.A(net20),
    .Y(_0725_));
 sky130_fd_sc_hd__a22o_4 _3558_ (.A1(net156),
    .A2(_0725_),
    .B1(\core_1.ew_mem_access ),
    .B2(\core_1.ew_submit ),
    .X(_0726_));
 sky130_fd_sc_hd__or2_2 _3559_ (.A(\core_1.execute.alu_mul_div.i_div ),
    .B(\core_1.execute.alu_mul_div.i_mod ),
    .X(_0727_));
 sky130_fd_sc_hd__nand2_1 _3560_ (.A(\core_1.decode.o_submit ),
    .B(_0727_),
    .Y(_0728_));
 sky130_fd_sc_hd__nand2_4 _3561_ (.A(\core_1.decode.o_submit ),
    .B(\core_1.execute.alu_mul_div.i_mul ),
    .Y(_0729_));
 sky130_fd_sc_hd__nand2_1 _3562_ (.A(_0728_),
    .B(_0729_),
    .Y(_0730_));
 sky130_fd_sc_hd__or2_2 _3563_ (.A(\core_1.execute.alu_mul_div.comp ),
    .B(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__or2_1 _3564_ (.A(_0726_),
    .B(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__or3_1 _3565_ (.A(_0690_),
    .B(_0724_),
    .C(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__inv_2 _3566_ (.A(_0733_),
    .Y(_0734_));
 sky130_fd_sc_hd__or2_4 _3567_ (.A(_0690_),
    .B(_0734_),
    .X(_0735_));
 sky130_fd_sc_hd__inv_2 _3568_ (.A(_0735_),
    .Y(_0736_));
 sky130_fd_sc_hd__nor2_2 _3569_ (.A(\core_1.decode.input_valid ),
    .B(_0736_),
    .Y(_0737_));
 sky130_fd_sc_hd__o21ai_1 _3570_ (.A1(_0664_),
    .A2(net70),
    .B1(_0737_),
    .Y(_0738_));
 sky130_fd_sc_hd__mux2_2 _3571_ (.A0(net38),
    .A1(\core_1.fetch.out_buffer_data_instr[0] ),
    .S(_0662_),
    .X(_0739_));
 sky130_fd_sc_hd__mux2_4 _3572_ (.A0(net49),
    .A1(\core_1.fetch.out_buffer_data_instr[1] ),
    .S(_0662_),
    .X(_0740_));
 sky130_fd_sc_hd__or2b_1 _3573_ (.A(_0739_),
    .B_N(_0740_),
    .X(_0741_));
 sky130_fd_sc_hd__mux2_2 _3574_ (.A0(net60),
    .A1(\core_1.fetch.out_buffer_data_instr[2] ),
    .S(_0663_),
    .X(_0742_));
 sky130_fd_sc_hd__mux2_2 _3575_ (.A0(net63),
    .A1(\core_1.fetch.out_buffer_data_instr[3] ),
    .S(_0663_),
    .X(_0743_));
 sky130_fd_sc_hd__nand2_1 _3576_ (.A(_0742_),
    .B(_0743_),
    .Y(_0744_));
 sky130_fd_sc_hd__nor2_1 _3577_ (.A(_0741_),
    .B(_0744_),
    .Y(_0745_));
 sky130_fd_sc_hd__mux2_4 _3578_ (.A0(net48),
    .A1(\core_1.fetch.out_buffer_data_instr[19] ),
    .S(\core_1.fetch.out_buffer_valid ),
    .X(_0746_));
 sky130_fd_sc_hd__mux2_4 _3579_ (.A0(net46),
    .A1(\core_1.fetch.out_buffer_data_instr[17] ),
    .S(\core_1.fetch.out_buffer_valid ),
    .X(_0747_));
 sky130_fd_sc_hd__mux2_4 _3580_ (.A0(net56),
    .A1(\core_1.fetch.out_buffer_data_instr[26] ),
    .S(_0661_),
    .X(_0748_));
 sky130_fd_sc_hd__mux2_4 _3581_ (.A0(net54),
    .A1(\core_1.fetch.out_buffer_data_instr[24] ),
    .S(_0661_),
    .X(_0749_));
 sky130_fd_sc_hd__or4b_1 _3582_ (.A(_0740_),
    .B(_0748_),
    .C(_0749_),
    .D_N(_0739_),
    .X(_0750_));
 sky130_fd_sc_hd__mux2_4 _3583_ (.A0(net61),
    .A1(\core_1.fetch.out_buffer_data_instr[30] ),
    .S(_0662_),
    .X(_0751_));
 sky130_fd_sc_hd__mux2_4 _3584_ (.A0(net50),
    .A1(\core_1.fetch.out_buffer_data_instr[20] ),
    .S(\core_1.fetch.out_buffer_valid ),
    .X(_0752_));
 sky130_fd_sc_hd__mux2_4 _3585_ (.A0(net47),
    .A1(\core_1.fetch.out_buffer_data_instr[18] ),
    .S(\core_1.fetch.out_buffer_valid ),
    .X(_0753_));
 sky130_fd_sc_hd__mux2_4 _3586_ (.A0(net53),
    .A1(\core_1.fetch.out_buffer_data_instr[23] ),
    .S(_0661_),
    .X(_0754_));
 sky130_fd_sc_hd__or4_1 _3587_ (.A(_0751_),
    .B(_0752_),
    .C(_0753_),
    .D(_0754_),
    .X(_0755_));
 sky130_fd_sc_hd__mux2_4 _3588_ (.A0(net58),
    .A1(\core_1.fetch.out_buffer_data_instr[28] ),
    .S(_0662_),
    .X(_0756_));
 sky130_fd_sc_hd__mux2_4 _3589_ (.A0(net45),
    .A1(\core_1.fetch.out_buffer_data_instr[16] ),
    .S(\core_1.fetch.out_buffer_valid ),
    .X(_0757_));
 sky130_fd_sc_hd__mux2_4 _3590_ (.A0(net51),
    .A1(\core_1.fetch.out_buffer_data_instr[21] ),
    .S(_0661_),
    .X(_0758_));
 sky130_fd_sc_hd__or2b_1 _3591_ (.A(\core_1.fetch.out_buffer_data_instr[31] ),
    .B_N(_0662_),
    .X(_0759_));
 sky130_fd_sc_hd__o21a_1 _3592_ (.A1(_0662_),
    .A2(net62),
    .B1(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__or4_1 _3593_ (.A(_0756_),
    .B(_0757_),
    .C(_0758_),
    .D(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__or2b_1 _3594_ (.A(\core_1.fetch.out_buffer_data_instr[25] ),
    .B_N(_0661_),
    .X(_0762_));
 sky130_fd_sc_hd__o21a_2 _3595_ (.A1(_0662_),
    .A2(net55),
    .B1(_0762_),
    .X(_0763_));
 sky130_fd_sc_hd__or2b_1 _3596_ (.A(\core_1.fetch.out_buffer_data_instr[27] ),
    .B_N(_0661_),
    .X(_0764_));
 sky130_fd_sc_hd__o21a_2 _3597_ (.A1(_0662_),
    .A2(net57),
    .B1(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__mux2_4 _3598_ (.A0(net52),
    .A1(\core_1.fetch.out_buffer_data_instr[22] ),
    .S(_0661_),
    .X(_0766_));
 sky130_fd_sc_hd__mux2_4 _3599_ (.A0(net59),
    .A1(\core_1.fetch.out_buffer_data_instr[29] ),
    .S(_0662_),
    .X(_0767_));
 sky130_fd_sc_hd__or4_1 _3600_ (.A(_0763_),
    .B(_0765_),
    .C(_0766_),
    .D(_0767_),
    .X(_0768_));
 sky130_fd_sc_hd__or3_2 _3601_ (.A(_0755_),
    .B(_0761_),
    .C(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__or4_1 _3602_ (.A(_0746_),
    .B(_0747_),
    .C(_0750_),
    .D(_0769_),
    .X(_0770_));
 sky130_fd_sc_hd__a211oi_1 _3603_ (.A1(_0741_),
    .A2(_0770_),
    .B1(_0742_),
    .C1(_0743_),
    .Y(_0771_));
 sky130_fd_sc_hd__mux2_2 _3604_ (.A0(net64),
    .A1(\core_1.fetch.out_buffer_data_instr[4] ),
    .S(_0663_),
    .X(_0772_));
 sky130_fd_sc_hd__mux2_1 _3605_ (.A0(net66),
    .A1(\core_1.fetch.out_buffer_data_instr[6] ),
    .S(_0663_),
    .X(_0773_));
 sky130_fd_sc_hd__mux2_2 _3606_ (.A0(net65),
    .A1(\core_1.fetch.out_buffer_data_instr[5] ),
    .S(_0663_),
    .X(_0774_));
 sky130_fd_sc_hd__nor2_1 _3607_ (.A(_0773_),
    .B(_0774_),
    .Y(_0775_));
 sky130_fd_sc_hd__o211a_1 _3608_ (.A1(_0745_),
    .A2(_0771_),
    .B1(_0772_),
    .C1(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__clkinv_4 _3609_ (.A(\core_1.fetch.pc_reset_override ),
    .Y(_0777_));
 sky130_fd_sc_hd__o221a_2 _3610_ (.A1(_0660_),
    .A2(\core_1.fetch.dbg_out ),
    .B1(_0738_),
    .B2(_0776_),
    .C1(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__nor2_8 _3611_ (.A(_0659_),
    .B(_0778_),
    .Y(_0779_));
 sky130_fd_sc_hd__clkbuf_8 _3612_ (.A(_0779_),
    .X(net177));
 sky130_fd_sc_hd__inv_2 _3613_ (.A(_0684_),
    .Y(net108));
 sky130_fd_sc_hd__inv_2 _3614_ (.A(_0674_),
    .Y(net109));
 sky130_fd_sc_hd__inv_2 _3615_ (.A(_0672_),
    .Y(net110));
 sky130_fd_sc_hd__inv_2 _3616_ (.A(_0669_),
    .Y(net111));
 sky130_fd_sc_hd__inv_2 _3617_ (.A(_0680_),
    .Y(net112));
 sky130_fd_sc_hd__clkinv_2 _3618_ (.A(_0677_),
    .Y(net113));
 sky130_fd_sc_hd__clkinv_2 _3619_ (.A(_0671_),
    .Y(net114));
 sky130_fd_sc_hd__inv_2 _3620_ (.A(_0675_),
    .Y(net115));
 sky130_fd_sc_hd__buf_4 _3621_ (.A(\core_1.decode.oc_alu_mode[4] ),
    .X(_0780_));
 sky130_fd_sc_hd__or2b_1 _3622_ (.A(\core_1.decode.i_instr_l[2] ),
    .B_N(\core_1.decode.i_instr_l[3] ),
    .X(_0781_));
 sky130_fd_sc_hd__inv_2 _3623_ (.A(\core_1.decode.i_instr_l[0] ),
    .Y(_0782_));
 sky130_fd_sc_hd__or2_1 _3624_ (.A(\core_1.decode.i_instr_l[1] ),
    .B(_0782_),
    .X(_0783_));
 sky130_fd_sc_hd__or2_1 _3625_ (.A(_0781_),
    .B(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__nand2_1 _3626_ (.A(\core_1.decode.i_instr_l[1] ),
    .B(\core_1.decode.i_instr_l[0] ),
    .Y(_0785_));
 sky130_fd_sc_hd__or2b_1 _3627_ (.A(\core_1.decode.i_instr_l[3] ),
    .B_N(\core_1.decode.i_instr_l[2] ),
    .X(_0786_));
 sky130_fd_sc_hd__buf_2 _3628_ (.A(_0786_),
    .X(_0787_));
 sky130_fd_sc_hd__or2_2 _3629_ (.A(\core_1.decode.i_instr_l[1] ),
    .B(\core_1.decode.i_instr_l[0] ),
    .X(_0788_));
 sky130_fd_sc_hd__or2_1 _3630_ (.A(_0781_),
    .B(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__o21a_1 _3631_ (.A1(_0785_),
    .A2(_0787_),
    .B1(_0789_),
    .X(_0790_));
 sky130_fd_sc_hd__or3_1 _3632_ (.A(\core_1.decode.i_instr_l[6] ),
    .B(\core_1.decode.i_instr_l[5] ),
    .C(\core_1.decode.i_instr_l[4] ),
    .X(_0791_));
 sky130_fd_sc_hd__a21oi_1 _3633_ (.A1(_0784_),
    .A2(_0790_),
    .B1(_0791_),
    .Y(_0792_));
 sky130_fd_sc_hd__or3b_1 _3634_ (.A(\core_1.decode.i_instr_l[6] ),
    .B(\core_1.decode.i_instr_l[4] ),
    .C_N(\core_1.decode.i_instr_l[5] ),
    .X(_0793_));
 sky130_fd_sc_hd__or3_1 _3635_ (.A(\core_1.decode.i_instr_l[3] ),
    .B(\core_1.decode.i_instr_l[2] ),
    .C(_0788_),
    .X(_0794_));
 sky130_fd_sc_hd__nor2_1 _3636_ (.A(_0793_),
    .B(_0794_),
    .Y(_0795_));
 sky130_fd_sc_hd__nor3_2 _3637_ (.A(\core_1.decode.i_instr_l[6] ),
    .B(\core_1.decode.i_instr_l[5] ),
    .C(\core_1.decode.i_instr_l[4] ),
    .Y(_0796_));
 sky130_fd_sc_hd__nand2_1 _3638_ (.A(\core_1.decode.i_instr_l[1] ),
    .B(_0782_),
    .Y(_0797_));
 sky130_fd_sc_hd__nor2_1 _3639_ (.A(_0787_),
    .B(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hd__clkbuf_4 _3640_ (.A(_0793_),
    .X(_0799_));
 sky130_fd_sc_hd__or3_2 _3641_ (.A(\core_1.decode.i_instr_l[3] ),
    .B(\core_1.decode.i_instr_l[2] ),
    .C(_0797_),
    .X(_0800_));
 sky130_fd_sc_hd__nor2_1 _3642_ (.A(_0799_),
    .B(_0800_),
    .Y(_0801_));
 sky130_fd_sc_hd__a21o_1 _3643_ (.A1(_0796_),
    .A2(_0798_),
    .B1(_0801_),
    .X(_0802_));
 sky130_fd_sc_hd__clkbuf_4 _3644_ (.A(_0791_),
    .X(_0803_));
 sky130_fd_sc_hd__or3_1 _3645_ (.A(\core_1.decode.i_instr_l[3] ),
    .B(\core_1.decode.i_instr_l[2] ),
    .C(_0785_),
    .X(_0804_));
 sky130_fd_sc_hd__clkbuf_2 _3646_ (.A(_0804_),
    .X(_0805_));
 sky130_fd_sc_hd__nor2_2 _3647_ (.A(_0799_),
    .B(_0781_),
    .Y(_0806_));
 sky130_fd_sc_hd__o21bai_1 _3648_ (.A1(_0803_),
    .A2(_0805_),
    .B1_N(_0806_),
    .Y(_0807_));
 sky130_fd_sc_hd__or4_1 _3649_ (.A(_0792_),
    .B(_0795_),
    .C(_0802_),
    .D(_0807_),
    .X(_0808_));
 sky130_fd_sc_hd__nor2_2 _3650_ (.A(\core_1.decode.i_flush ),
    .B(net71),
    .Y(_0809_));
 sky130_fd_sc_hd__o211ai_4 _3651_ (.A1(\core_1.decode.input_valid ),
    .A2(\core_1.decode.i_submit ),
    .B1(_0735_),
    .C1(_0809_),
    .Y(_0810_));
 sky130_fd_sc_hd__inv_4 _3652_ (.A(_0810_),
    .Y(_0811_));
 sky130_fd_sc_hd__buf_4 _3653_ (.A(_0811_),
    .X(_0812_));
 sky130_fd_sc_hd__mux2_1 _3654_ (.A0(_0780_),
    .A1(_0808_),
    .S(_0812_),
    .X(_0813_));
 sky130_fd_sc_hd__clkbuf_1 _3655_ (.A(_0813_),
    .X(_0007_));
 sky130_fd_sc_hd__buf_4 _3656_ (.A(\core_1.decode.oc_alu_mode[9] ),
    .X(_0814_));
 sky130_fd_sc_hd__clkbuf_4 _3657_ (.A(_0810_),
    .X(_0815_));
 sky130_fd_sc_hd__clkbuf_4 _3658_ (.A(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__or3b_1 _3659_ (.A(\core_1.decode.i_instr_l[6] ),
    .B(\core_1.decode.i_instr_l[5] ),
    .C_N(\core_1.decode.i_instr_l[4] ),
    .X(_0817_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _3660_ (.A(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__clkbuf_4 _3661_ (.A(_0818_),
    .X(_0819_));
 sky130_fd_sc_hd__nor2_2 _3662_ (.A(_0810_),
    .B(_0819_),
    .Y(_0820_));
 sky130_fd_sc_hd__a21oi_1 _3663_ (.A1(_0785_),
    .A2(_0788_),
    .B1(_0787_),
    .Y(_0821_));
 sky130_fd_sc_hd__a22o_1 _3664_ (.A1(_0814_),
    .A2(_0816_),
    .B1(_0820_),
    .B2(_0821_),
    .X(_0012_));
 sky130_fd_sc_hd__buf_6 _3665_ (.A(\core_1.decode.oc_alu_mode[12] ),
    .X(_0822_));
 sky130_fd_sc_hd__nor2_1 _3666_ (.A(_0783_),
    .B(_0787_),
    .Y(_0823_));
 sky130_fd_sc_hd__nor2_1 _3667_ (.A(_0798_),
    .B(_0823_),
    .Y(_0824_));
 sky130_fd_sc_hd__inv_2 _3668_ (.A(_0824_),
    .Y(_0825_));
 sky130_fd_sc_hd__nor2_1 _3669_ (.A(_0815_),
    .B(_0799_),
    .Y(_0826_));
 sky130_fd_sc_hd__a22o_1 _3670_ (.A1(_0822_),
    .A2(_0816_),
    .B1(_0825_),
    .B2(_0826_),
    .X(_0002_));
 sky130_fd_sc_hd__nand2_1 _3671_ (.A(\core_1.decode.i_instr_l[3] ),
    .B(\core_1.decode.i_instr_l[2] ),
    .Y(_0827_));
 sky130_fd_sc_hd__or2_2 _3672_ (.A(\core_1.decode.i_instr_l[1] ),
    .B(_0827_),
    .X(_0828_));
 sky130_fd_sc_hd__inv_2 _3673_ (.A(_0828_),
    .Y(_0829_));
 sky130_fd_sc_hd__clkbuf_4 _3674_ (.A(_0810_),
    .X(_0830_));
 sky130_fd_sc_hd__clkbuf_4 _3675_ (.A(\core_1.execute.alu_mul_div.i_div ),
    .X(_0831_));
 sky130_fd_sc_hd__a32o_1 _3676_ (.A1(\core_1.decode.i_instr_l[0] ),
    .A2(_0820_),
    .A3(_0829_),
    .B1(_0830_),
    .B2(_0831_),
    .X(_0008_));
 sky130_fd_sc_hd__buf_4 _3677_ (.A(\core_1.decode.oc_alu_mode[6] ),
    .X(_0832_));
 sky130_fd_sc_hd__or2_1 _3678_ (.A(_0783_),
    .B(_0787_),
    .X(_0833_));
 sky130_fd_sc_hd__nand2_1 _3679_ (.A(_0789_),
    .B(_0833_),
    .Y(_0834_));
 sky130_fd_sc_hd__a22o_1 _3680_ (.A1(_0832_),
    .A2(_0816_),
    .B1(_0820_),
    .B2(_0834_),
    .X(_0009_));
 sky130_fd_sc_hd__buf_4 _3681_ (.A(\core_1.execute.alu_mul_div.i_mod ),
    .X(_0835_));
 sky130_fd_sc_hd__or2_1 _3682_ (.A(_0788_),
    .B(_0827_),
    .X(_0836_));
 sky130_fd_sc_hd__nor2_1 _3683_ (.A(_0799_),
    .B(_0836_),
    .Y(_0837_));
 sky130_fd_sc_hd__mux2_1 _3684_ (.A0(_0835_),
    .A1(_0837_),
    .S(_0812_),
    .X(_0838_));
 sky130_fd_sc_hd__clkbuf_1 _3685_ (.A(_0838_),
    .X(_0000_));
 sky130_fd_sc_hd__buf_4 _3686_ (.A(\core_1.decode.oc_alu_mode[2] ),
    .X(_0839_));
 sky130_fd_sc_hd__and2b_1 _3687_ (.A_N(\core_1.decode.i_instr_l[2] ),
    .B(\core_1.decode.i_instr_l[3] ),
    .X(_0840_));
 sky130_fd_sc_hd__nand2_1 _3688_ (.A(\core_1.decode.i_instr_l[1] ),
    .B(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__o22a_1 _3689_ (.A1(_0787_),
    .A2(_0797_),
    .B1(_0841_),
    .B2(_0782_),
    .X(_0842_));
 sky130_fd_sc_hd__nand2_1 _3690_ (.A(_0805_),
    .B(_0842_),
    .Y(_0843_));
 sky130_fd_sc_hd__a22o_1 _3691_ (.A1(_0839_),
    .A2(_0816_),
    .B1(_0820_),
    .B2(_0843_),
    .X(_0005_));
 sky130_fd_sc_hd__o22ai_2 _3692_ (.A1(_0805_),
    .A2(_0799_),
    .B1(_0784_),
    .B2(_0818_),
    .Y(_0844_));
 sky130_fd_sc_hd__mux2_1 _3693_ (.A0(\core_1.decode.oc_alu_mode[13] ),
    .A1(_0844_),
    .S(_0812_),
    .X(_0845_));
 sky130_fd_sc_hd__clkbuf_1 _3694_ (.A(_0845_),
    .X(_0003_));
 sky130_fd_sc_hd__buf_4 _3695_ (.A(\core_1.decode.oc_alu_mode[7] ),
    .X(_0846_));
 sky130_fd_sc_hd__or2_2 _3696_ (.A(_0785_),
    .B(_0827_),
    .X(_0847_));
 sky130_fd_sc_hd__nor2_1 _3697_ (.A(_0819_),
    .B(_0847_),
    .Y(_0848_));
 sky130_fd_sc_hd__or2_1 _3698_ (.A(_0788_),
    .B(_0787_),
    .X(_0849_));
 sky130_fd_sc_hd__and3_1 _3699_ (.A(_0800_),
    .B(_0849_),
    .C(_0847_),
    .X(_0850_));
 sky130_fd_sc_hd__nor2_1 _3700_ (.A(_0803_),
    .B(_0850_),
    .Y(_0851_));
 sky130_fd_sc_hd__or2_2 _3701_ (.A(_0797_),
    .B(_0827_),
    .X(_0852_));
 sky130_fd_sc_hd__nor2_1 _3702_ (.A(_0803_),
    .B(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__or3_1 _3703_ (.A(\core_1.decode.i_instr_l[3] ),
    .B(\core_1.decode.i_instr_l[2] ),
    .C(_0783_),
    .X(_0854_));
 sky130_fd_sc_hd__nor2_1 _3704_ (.A(_0799_),
    .B(_0854_),
    .Y(_0855_));
 sky130_fd_sc_hd__a21o_1 _3705_ (.A1(_0796_),
    .A2(_0823_),
    .B1(_0855_),
    .X(_0856_));
 sky130_fd_sc_hd__or4_1 _3706_ (.A(_0848_),
    .B(_0851_),
    .C(_0853_),
    .D(_0856_),
    .X(_0857_));
 sky130_fd_sc_hd__mux2_1 _3707_ (.A0(_0846_),
    .A1(_0857_),
    .S(_0812_),
    .X(_0858_));
 sky130_fd_sc_hd__clkbuf_1 _3708_ (.A(_0858_),
    .X(_0010_));
 sky130_fd_sc_hd__buf_2 _3709_ (.A(\core_1.execute.alu_mul_div.i_mul ),
    .X(_0859_));
 sky130_fd_sc_hd__clkbuf_4 _3710_ (.A(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__nor2_1 _3711_ (.A(_0788_),
    .B(_0827_),
    .Y(_0861_));
 sky130_fd_sc_hd__a22o_1 _3712_ (.A1(_0860_),
    .A2(_0816_),
    .B1(_0820_),
    .B2(_0861_),
    .X(_0011_));
 sky130_fd_sc_hd__buf_4 _3713_ (.A(\core_1.decode.oc_alu_mode[11] ),
    .X(_0862_));
 sky130_fd_sc_hd__buf_4 _3714_ (.A(_0862_),
    .X(_0863_));
 sky130_fd_sc_hd__a21oi_1 _3715_ (.A1(_0828_),
    .A2(_0841_),
    .B1(_0803_),
    .Y(_0864_));
 sky130_fd_sc_hd__mux2_1 _3716_ (.A0(_0863_),
    .A1(_0864_),
    .S(_0812_),
    .X(_0865_));
 sky130_fd_sc_hd__clkbuf_1 _3717_ (.A(_0865_),
    .X(_0001_));
 sky130_fd_sc_hd__nor2_1 _3718_ (.A(_0785_),
    .B(_0787_),
    .Y(_0866_));
 sky130_fd_sc_hd__a22o_1 _3719_ (.A1(\core_1.decode.oc_alu_mode[3] ),
    .A2(_0816_),
    .B1(_0866_),
    .B2(_0826_),
    .X(_0006_));
 sky130_fd_sc_hd__o32a_1 _3720_ (.A1(\core_1.decode.i_instr_l[0] ),
    .A2(_0819_),
    .A3(_0841_),
    .B1(_0849_),
    .B2(_0799_),
    .X(_0867_));
 sky130_fd_sc_hd__inv_2 _3721_ (.A(_0867_),
    .Y(_0868_));
 sky130_fd_sc_hd__mux2_1 _3722_ (.A0(\core_1.decode.oc_alu_mode[1] ),
    .A1(_0868_),
    .S(_0812_),
    .X(_0869_));
 sky130_fd_sc_hd__clkbuf_1 _3723_ (.A(_0869_),
    .X(_0004_));
 sky130_fd_sc_hd__nor2_4 _3724_ (.A(\core_1.fetch.pc_flush_override ),
    .B(\core_1.decode.i_flush ),
    .Y(_0870_));
 sky130_fd_sc_hd__buf_4 _3725_ (.A(_0870_),
    .X(_0871_));
 sky130_fd_sc_hd__inv_2 _3726_ (.A(\core_1.fetch.prev_request_pc[14] ),
    .Y(_0872_));
 sky130_fd_sc_hd__o21ai_1 _3727_ (.A1(_0663_),
    .A2(net62),
    .B1(_0759_),
    .Y(_0873_));
 sky130_fd_sc_hd__o2bb2a_1 _3728_ (.A1_N(_0872_),
    .A2_N(_0751_),
    .B1(_0873_),
    .B2(\core_1.fetch.prev_request_pc[15] ),
    .X(_0874_));
 sky130_fd_sc_hd__inv_2 _3729_ (.A(\core_1.fetch.prev_request_pc[12] ),
    .Y(_0875_));
 sky130_fd_sc_hd__inv_2 _3730_ (.A(\core_1.fetch.prev_request_pc[13] ),
    .Y(_0876_));
 sky130_fd_sc_hd__inv_2 _3731_ (.A(\core_1.fetch.prev_request_pc[6] ),
    .Y(_0877_));
 sky130_fd_sc_hd__inv_2 _3732_ (.A(\core_1.fetch.prev_request_pc[7] ),
    .Y(_0878_));
 sky130_fd_sc_hd__inv_2 _3733_ (.A(\core_1.fetch.prev_request_pc[5] ),
    .Y(_0879_));
 sky130_fd_sc_hd__inv_2 _3734_ (.A(\core_1.fetch.prev_request_pc[4] ),
    .Y(_0880_));
 sky130_fd_sc_hd__inv_2 _3735_ (.A(\core_1.fetch.prev_request_pc[3] ),
    .Y(_0881_));
 sky130_fd_sc_hd__inv_2 _3736_ (.A(\core_1.fetch.prev_request_pc[2] ),
    .Y(_0882_));
 sky130_fd_sc_hd__inv_2 _3737_ (.A(\core_1.fetch.prev_request_pc[1] ),
    .Y(_0883_));
 sky130_fd_sc_hd__inv_2 _3738_ (.A(\core_1.fetch.prev_request_pc[0] ),
    .Y(_0884_));
 sky130_fd_sc_hd__a211o_1 _3739_ (.A1(_0883_),
    .A2(_0747_),
    .B1(_0757_),
    .C1(_0884_),
    .X(_0885_));
 sky130_fd_sc_hd__o221a_1 _3740_ (.A1(_0882_),
    .A2(_0753_),
    .B1(_0747_),
    .B2(_0883_),
    .C1(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__a221o_1 _3741_ (.A1(_0881_),
    .A2(_0746_),
    .B1(_0753_),
    .B2(_0882_),
    .C1(_0886_),
    .X(_0887_));
 sky130_fd_sc_hd__o221a_1 _3742_ (.A1(_0881_),
    .A2(_0746_),
    .B1(_0752_),
    .B2(_0880_),
    .C1(_0887_),
    .X(_0888_));
 sky130_fd_sc_hd__a221o_1 _3743_ (.A1(_0880_),
    .A2(_0752_),
    .B1(_0758_),
    .B2(_0879_),
    .C1(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__o221a_1 _3744_ (.A1(_0877_),
    .A2(_0766_),
    .B1(_0758_),
    .B2(_0879_),
    .C1(_0889_),
    .X(_0890_));
 sky130_fd_sc_hd__a221o_1 _3745_ (.A1(_0877_),
    .A2(_0766_),
    .B1(_0754_),
    .B2(_0878_),
    .C1(_0890_),
    .X(_0891_));
 sky130_fd_sc_hd__inv_2 _3746_ (.A(\core_1.fetch.prev_request_pc[8] ),
    .Y(_0892_));
 sky130_fd_sc_hd__o21ai_4 _3747_ (.A1(_0661_),
    .A2(net57),
    .B1(_0764_),
    .Y(_0893_));
 sky130_fd_sc_hd__inv_2 _3748_ (.A(\core_1.fetch.prev_request_pc[10] ),
    .Y(_0894_));
 sky130_fd_sc_hd__a2bb2o_1 _3749_ (.A1_N(\core_1.fetch.prev_request_pc[11] ),
    .A2_N(_0893_),
    .B1(_0748_),
    .B2(_0894_),
    .X(_0895_));
 sky130_fd_sc_hd__nand2_1 _3750_ (.A(\core_1.fetch.prev_request_pc[11] ),
    .B(_0893_),
    .Y(_0896_));
 sky130_fd_sc_hd__o21ai_1 _3751_ (.A1(_0894_),
    .A2(_0748_),
    .B1(_0896_),
    .Y(_0897_));
 sky130_fd_sc_hd__nor2_1 _3752_ (.A(_0895_),
    .B(_0897_),
    .Y(_0898_));
 sky130_fd_sc_hd__o21ai_4 _3753_ (.A1(_0661_),
    .A2(net55),
    .B1(_0762_),
    .Y(_0899_));
 sky130_fd_sc_hd__o2bb2a_1 _3754_ (.A1_N(_0749_),
    .A2_N(_0892_),
    .B1(\core_1.fetch.prev_request_pc[9] ),
    .B2(_0899_),
    .X(_0900_));
 sky130_fd_sc_hd__o2bb2a_1 _3755_ (.A1_N(\core_1.fetch.prev_request_pc[9] ),
    .A2_N(_0899_),
    .B1(_0754_),
    .B2(_0878_),
    .X(_0901_));
 sky130_fd_sc_hd__o2111a_1 _3756_ (.A1(_0892_),
    .A2(_0749_),
    .B1(_0898_),
    .C1(_0900_),
    .D1(_0901_),
    .X(_0902_));
 sky130_fd_sc_hd__a21oi_1 _3757_ (.A1(\core_1.fetch.prev_request_pc[9] ),
    .A2(_0899_),
    .B1(_0900_),
    .Y(_0903_));
 sky130_fd_sc_hd__a22o_1 _3758_ (.A1(_0895_),
    .A2(_0896_),
    .B1(_0898_),
    .B2(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__a21o_1 _3759_ (.A1(_0891_),
    .A2(_0902_),
    .B1(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__o21a_1 _3760_ (.A1(_0875_),
    .A2(_0756_),
    .B1(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__a221o_1 _3761_ (.A1(_0875_),
    .A2(_0756_),
    .B1(_0767_),
    .B2(_0876_),
    .C1(_0906_),
    .X(_0907_));
 sky130_fd_sc_hd__nand2_1 _3762_ (.A(\core_1.fetch.prev_request_pc[15] ),
    .B(_0873_),
    .Y(_0908_));
 sky130_fd_sc_hd__o221a_1 _3763_ (.A1(_0872_),
    .A2(_0751_),
    .B1(_0767_),
    .B2(_0876_),
    .C1(_0908_),
    .X(_0909_));
 sky130_fd_sc_hd__and2b_1 _3764_ (.A_N(_0874_),
    .B(_0908_),
    .X(_0910_));
 sky130_fd_sc_hd__a31o_1 _3765_ (.A1(_0874_),
    .A2(_0907_),
    .A3(_0909_),
    .B1(_0910_),
    .X(_0911_));
 sky130_fd_sc_hd__mux2_1 _3766_ (.A0(net69),
    .A1(\core_1.fetch.out_buffer_data_instr[9] ),
    .S(_0663_),
    .X(_0912_));
 sky130_fd_sc_hd__mux2_2 _3767_ (.A0(net67),
    .A1(\core_1.fetch.out_buffer_data_instr[7] ),
    .S(_0663_),
    .X(_0913_));
 sky130_fd_sc_hd__mux2_2 _3768_ (.A0(net39),
    .A1(\core_1.fetch.out_buffer_data_instr[10] ),
    .S(_0663_),
    .X(_0914_));
 sky130_fd_sc_hd__mux2_1 _3769_ (.A0(net68),
    .A1(\core_1.fetch.out_buffer_data_instr[8] ),
    .S(_0664_),
    .X(_0915_));
 sky130_fd_sc_hd__o41a_2 _3770_ (.A1(_0912_),
    .A2(_0913_),
    .A3(_0914_),
    .A4(_0915_),
    .B1(_0745_),
    .X(_0916_));
 sky130_fd_sc_hd__or3_1 _3771_ (.A(\core_1.fetch.pc_reset_override ),
    .B(_0773_),
    .C(_0774_),
    .X(_0917_));
 sky130_fd_sc_hd__or4b_4 _3772_ (.A(_0772_),
    .B(_0744_),
    .C(_0917_),
    .D_N(_0740_),
    .X(_0918_));
 sky130_fd_sc_hd__a21oi_4 _3773_ (.A1(_0911_),
    .A2(_0916_),
    .B1(_0918_),
    .Y(_0919_));
 sky130_fd_sc_hd__clkbuf_4 _3774_ (.A(_0919_),
    .X(_0920_));
 sky130_fd_sc_hd__or2_4 _3775_ (.A(\core_1.fetch.pc_flush_override ),
    .B(\core_1.decode.i_flush ),
    .X(_0921_));
 sky130_fd_sc_hd__a21o_1 _3776_ (.A1(_0757_),
    .A2(_0920_),
    .B1(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__buf_4 _3777_ (.A(_0920_),
    .X(_0923_));
 sky130_fd_sc_hd__nor2_1 _3778_ (.A(\core_1.fetch.prev_request_pc[0] ),
    .B(_0923_),
    .Y(_0924_));
 sky130_fd_sc_hd__buf_4 _3779_ (.A(_0777_),
    .X(_0925_));
 sky130_fd_sc_hd__o221a_1 _3780_ (.A1(net72),
    .A2(_0871_),
    .B1(_0922_),
    .B2(_0924_),
    .C1(_0925_),
    .X(net161));
 sky130_fd_sc_hd__clkbuf_4 _3781_ (.A(_0921_),
    .X(_0926_));
 sky130_fd_sc_hd__xor2_1 _3782_ (.A(\core_1.fetch.prev_request_pc[1] ),
    .B(\core_1.fetch.prev_request_pc[0] ),
    .X(_0927_));
 sky130_fd_sc_hd__mux2_1 _3783_ (.A0(_0927_),
    .A1(_0747_),
    .S(_0920_),
    .X(_0928_));
 sky130_fd_sc_hd__or2_1 _3784_ (.A(net79),
    .B(_0870_),
    .X(_0929_));
 sky130_fd_sc_hd__o211a_1 _3785_ (.A1(_0926_),
    .A2(_0928_),
    .B1(_0929_),
    .C1(_0925_),
    .X(net168));
 sky130_fd_sc_hd__a21oi_1 _3786_ (.A1(\core_1.fetch.prev_request_pc[1] ),
    .A2(\core_1.fetch.prev_request_pc[0] ),
    .B1(\core_1.fetch.prev_request_pc[2] ),
    .Y(_0930_));
 sky130_fd_sc_hd__and3_1 _3787_ (.A(\core_1.fetch.prev_request_pc[2] ),
    .B(\core_1.fetch.prev_request_pc[1] ),
    .C(\core_1.fetch.prev_request_pc[0] ),
    .X(_0931_));
 sky130_fd_sc_hd__nor3_1 _3788_ (.A(_0923_),
    .B(_0930_),
    .C(_0931_),
    .Y(_0932_));
 sky130_fd_sc_hd__clkbuf_4 _3789_ (.A(_0920_),
    .X(_0933_));
 sky130_fd_sc_hd__a21o_1 _3790_ (.A1(_0753_),
    .A2(_0933_),
    .B1(_0926_),
    .X(_0934_));
 sky130_fd_sc_hd__o221a_1 _3791_ (.A1(net80),
    .A2(_0871_),
    .B1(_0932_),
    .B2(_0934_),
    .C1(_0925_),
    .X(net169));
 sky130_fd_sc_hd__and2_1 _3792_ (.A(\core_1.fetch.prev_request_pc[3] ),
    .B(_0931_),
    .X(_0935_));
 sky130_fd_sc_hd__or2_1 _3793_ (.A(\core_1.fetch.prev_request_pc[3] ),
    .B(_0931_),
    .X(_0936_));
 sky130_fd_sc_hd__nor3b_1 _3794_ (.A(_0923_),
    .B(_0935_),
    .C_N(_0936_),
    .Y(_0937_));
 sky130_fd_sc_hd__a21o_1 _3795_ (.A1(_0746_),
    .A2(_0933_),
    .B1(_0926_),
    .X(_0938_));
 sky130_fd_sc_hd__o221a_1 _3796_ (.A1(net81),
    .A2(_0871_),
    .B1(_0937_),
    .B2(_0938_),
    .C1(_0925_),
    .X(net170));
 sky130_fd_sc_hd__xnor2_1 _3797_ (.A(\core_1.fetch.prev_request_pc[4] ),
    .B(_0935_),
    .Y(_0939_));
 sky130_fd_sc_hd__nor2_1 _3798_ (.A(_0923_),
    .B(_0939_),
    .Y(_0940_));
 sky130_fd_sc_hd__a21o_1 _3799_ (.A1(_0752_),
    .A2(_0933_),
    .B1(_0926_),
    .X(_0941_));
 sky130_fd_sc_hd__o221a_1 _3800_ (.A1(net82),
    .A2(_0871_),
    .B1(_0940_),
    .B2(_0941_),
    .C1(_0925_),
    .X(net171));
 sky130_fd_sc_hd__and3_1 _3801_ (.A(\core_1.fetch.prev_request_pc[5] ),
    .B(\core_1.fetch.prev_request_pc[4] ),
    .C(_0935_),
    .X(_0942_));
 sky130_fd_sc_hd__a21oi_1 _3802_ (.A1(\core_1.fetch.prev_request_pc[4] ),
    .A2(_0935_),
    .B1(\core_1.fetch.prev_request_pc[5] ),
    .Y(_0943_));
 sky130_fd_sc_hd__nor3_1 _3803_ (.A(_0923_),
    .B(_0942_),
    .C(_0943_),
    .Y(_0944_));
 sky130_fd_sc_hd__a21o_1 _3804_ (.A1(_0758_),
    .A2(_0933_),
    .B1(_0926_),
    .X(_0945_));
 sky130_fd_sc_hd__o221a_1 _3805_ (.A1(net83),
    .A2(_0871_),
    .B1(_0944_),
    .B2(_0945_),
    .C1(_0777_),
    .X(net172));
 sky130_fd_sc_hd__and2_1 _3806_ (.A(\core_1.fetch.prev_request_pc[6] ),
    .B(_0942_),
    .X(_0946_));
 sky130_fd_sc_hd__nor2_1 _3807_ (.A(\core_1.fetch.prev_request_pc[6] ),
    .B(_0942_),
    .Y(_0947_));
 sky130_fd_sc_hd__nor3_1 _3808_ (.A(_0923_),
    .B(_0946_),
    .C(_0947_),
    .Y(_0948_));
 sky130_fd_sc_hd__a21o_1 _3809_ (.A1(_0766_),
    .A2(_0933_),
    .B1(_0926_),
    .X(_0949_));
 sky130_fd_sc_hd__o221a_1 _3810_ (.A1(net84),
    .A2(_0871_),
    .B1(_0948_),
    .B2(_0949_),
    .C1(_0777_),
    .X(net173));
 sky130_fd_sc_hd__xnor2_1 _3811_ (.A(\core_1.fetch.prev_request_pc[7] ),
    .B(_0946_),
    .Y(_0950_));
 sky130_fd_sc_hd__nor2_1 _3812_ (.A(_0923_),
    .B(_0950_),
    .Y(_0951_));
 sky130_fd_sc_hd__a21o_1 _3813_ (.A1(_0754_),
    .A2(_0933_),
    .B1(_0926_),
    .X(_0952_));
 sky130_fd_sc_hd__o221a_1 _3814_ (.A1(net85),
    .A2(_0870_),
    .B1(_0951_),
    .B2(_0952_),
    .C1(_0777_),
    .X(net174));
 sky130_fd_sc_hd__and3_1 _3815_ (.A(\core_1.fetch.prev_request_pc[8] ),
    .B(\core_1.fetch.prev_request_pc[7] ),
    .C(_0946_),
    .X(_0953_));
 sky130_fd_sc_hd__a21oi_1 _3816_ (.A1(\core_1.fetch.prev_request_pc[7] ),
    .A2(_0946_),
    .B1(\core_1.fetch.prev_request_pc[8] ),
    .Y(_0954_));
 sky130_fd_sc_hd__o31a_1 _3817_ (.A1(_0919_),
    .A2(_0953_),
    .A3(_0954_),
    .B1(_0870_),
    .X(_0955_));
 sky130_fd_sc_hd__a21bo_1 _3818_ (.A1(_0749_),
    .A2(_0933_),
    .B1_N(_0955_),
    .X(_0956_));
 sky130_fd_sc_hd__o211a_1 _3819_ (.A1(net86),
    .A2(_0871_),
    .B1(_0956_),
    .C1(_0925_),
    .X(net175));
 sky130_fd_sc_hd__and2_1 _3820_ (.A(\core_1.fetch.prev_request_pc[9] ),
    .B(_0953_),
    .X(_0957_));
 sky130_fd_sc_hd__nor2_1 _3821_ (.A(\core_1.fetch.prev_request_pc[9] ),
    .B(_0953_),
    .Y(_0958_));
 sky130_fd_sc_hd__o31a_1 _3822_ (.A1(_0919_),
    .A2(_0957_),
    .A3(_0958_),
    .B1(_0870_),
    .X(_0959_));
 sky130_fd_sc_hd__a21bo_1 _3823_ (.A1(_0763_),
    .A2(_0933_),
    .B1_N(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__o211a_1 _3824_ (.A1(net87),
    .A2(_0871_),
    .B1(_0960_),
    .C1(_0925_),
    .X(net176));
 sky130_fd_sc_hd__xnor2_1 _3825_ (.A(\core_1.fetch.prev_request_pc[10] ),
    .B(_0957_),
    .Y(_0961_));
 sky130_fd_sc_hd__nor2_1 _3826_ (.A(_0920_),
    .B(_0961_),
    .Y(_0962_));
 sky130_fd_sc_hd__a211o_1 _3827_ (.A1(_0748_),
    .A2(_0920_),
    .B1(_0921_),
    .C1(_0962_),
    .X(_0963_));
 sky130_fd_sc_hd__o211a_1 _3828_ (.A1(net73),
    .A2(_0871_),
    .B1(_0963_),
    .C1(_0925_),
    .X(net162));
 sky130_fd_sc_hd__and3_1 _3829_ (.A(\core_1.fetch.prev_request_pc[11] ),
    .B(\core_1.fetch.prev_request_pc[10] ),
    .C(_0957_),
    .X(_0964_));
 sky130_fd_sc_hd__a21oi_1 _3830_ (.A1(\core_1.fetch.prev_request_pc[10] ),
    .A2(_0957_),
    .B1(\core_1.fetch.prev_request_pc[11] ),
    .Y(_0965_));
 sky130_fd_sc_hd__nor3_1 _3831_ (.A(_0923_),
    .B(_0964_),
    .C(_0965_),
    .Y(_0966_));
 sky130_fd_sc_hd__a21o_1 _3832_ (.A1(_0765_),
    .A2(_0933_),
    .B1(_0926_),
    .X(_0967_));
 sky130_fd_sc_hd__o221a_1 _3833_ (.A1(net74),
    .A2(_0870_),
    .B1(_0966_),
    .B2(_0967_),
    .C1(_0777_),
    .X(net163));
 sky130_fd_sc_hd__xnor2_1 _3834_ (.A(_0875_),
    .B(_0964_),
    .Y(_0968_));
 sky130_fd_sc_hd__mux2_1 _3835_ (.A0(_0968_),
    .A1(_0756_),
    .S(_0920_),
    .X(_0969_));
 sky130_fd_sc_hd__or2_1 _3836_ (.A(net75),
    .B(_0870_),
    .X(_0970_));
 sky130_fd_sc_hd__o211a_1 _3837_ (.A1(_0926_),
    .A2(_0969_),
    .B1(_0970_),
    .C1(_0925_),
    .X(net164));
 sky130_fd_sc_hd__and3_1 _3838_ (.A(\core_1.fetch.prev_request_pc[13] ),
    .B(\core_1.fetch.prev_request_pc[12] ),
    .C(_0964_),
    .X(_0971_));
 sky130_fd_sc_hd__a21oi_1 _3839_ (.A1(\core_1.fetch.prev_request_pc[12] ),
    .A2(_0964_),
    .B1(\core_1.fetch.prev_request_pc[13] ),
    .Y(_0972_));
 sky130_fd_sc_hd__nor3_1 _3840_ (.A(_0923_),
    .B(_0971_),
    .C(_0972_),
    .Y(_0973_));
 sky130_fd_sc_hd__a21o_1 _3841_ (.A1(_0767_),
    .A2(_0933_),
    .B1(_0921_),
    .X(_0974_));
 sky130_fd_sc_hd__o221a_1 _3842_ (.A1(net76),
    .A2(_0870_),
    .B1(_0973_),
    .B2(_0974_),
    .C1(_0777_),
    .X(net165));
 sky130_fd_sc_hd__nand2_1 _3843_ (.A(\core_1.fetch.prev_request_pc[14] ),
    .B(_0971_),
    .Y(_0975_));
 sky130_fd_sc_hd__o21ba_1 _3844_ (.A1(\core_1.fetch.prev_request_pc[14] ),
    .A2(_0971_),
    .B1_N(_0919_),
    .X(_0976_));
 sky130_fd_sc_hd__a221o_1 _3845_ (.A1(_0751_),
    .A2(_0920_),
    .B1(_0975_),
    .B2(_0976_),
    .C1(_0921_),
    .X(_0977_));
 sky130_fd_sc_hd__o211a_1 _3846_ (.A1(net77),
    .A2(_0871_),
    .B1(_0977_),
    .C1(_0925_),
    .X(net166));
 sky130_fd_sc_hd__xor2_1 _3847_ (.A(\core_1.fetch.prev_request_pc[15] ),
    .B(_0975_),
    .X(_0978_));
 sky130_fd_sc_hd__nor2_1 _3848_ (.A(_0923_),
    .B(_0978_),
    .Y(_0979_));
 sky130_fd_sc_hd__a21o_1 _3849_ (.A1(_0760_),
    .A2(_0920_),
    .B1(_0921_),
    .X(_0980_));
 sky130_fd_sc_hd__o221a_1 _3850_ (.A1(net78),
    .A2(_0870_),
    .B1(_0979_),
    .B2(_0980_),
    .C1(_0777_),
    .X(net167));
 sky130_fd_sc_hd__mux2_1 _3851_ (.A0(\core_1.fetch.prev_req_branch_pred ),
    .A1(_0920_),
    .S(net70),
    .X(_0981_));
 sky130_fd_sc_hd__clkbuf_1 _3852_ (.A(_0981_),
    .X(\core_1.fetch.current_req_branch_pred ));
 sky130_fd_sc_hd__nand2_4 _3853_ (.A(\core_1.ew_addr[0] ),
    .B(\core_1.ew_mem_width ),
    .Y(_0982_));
 sky130_fd_sc_hd__clkbuf_4 _3854_ (.A(_0982_),
    .X(_0983_));
 sky130_fd_sc_hd__buf_4 _3855_ (.A(_0983_),
    .X(net157));
 sky130_fd_sc_hd__and2_1 _3856_ (.A(\core_1.ew_data[0] ),
    .B(net157),
    .X(_0984_));
 sky130_fd_sc_hd__clkbuf_1 _3857_ (.A(_0984_),
    .X(net139));
 sky130_fd_sc_hd__and2_1 _3858_ (.A(\core_1.ew_data[1] ),
    .B(net157),
    .X(_0985_));
 sky130_fd_sc_hd__clkbuf_1 _3859_ (.A(_0985_),
    .X(net146));
 sky130_fd_sc_hd__and2_1 _3860_ (.A(\core_1.ew_data[2] ),
    .B(net157),
    .X(_0986_));
 sky130_fd_sc_hd__clkbuf_1 _3861_ (.A(_0986_),
    .X(net147));
 sky130_fd_sc_hd__and2_1 _3862_ (.A(\core_1.ew_data[3] ),
    .B(net157),
    .X(_0987_));
 sky130_fd_sc_hd__clkbuf_1 _3863_ (.A(_0987_),
    .X(net148));
 sky130_fd_sc_hd__and2_1 _3864_ (.A(\core_1.ew_data[4] ),
    .B(net157),
    .X(_0988_));
 sky130_fd_sc_hd__clkbuf_1 _3865_ (.A(_0988_),
    .X(net149));
 sky130_fd_sc_hd__and2_1 _3866_ (.A(\core_1.ew_data[5] ),
    .B(net157),
    .X(_0989_));
 sky130_fd_sc_hd__clkbuf_1 _3867_ (.A(_0989_),
    .X(net150));
 sky130_fd_sc_hd__and2_1 _3868_ (.A(\core_1.ew_data[6] ),
    .B(net157),
    .X(_0990_));
 sky130_fd_sc_hd__clkbuf_1 _3869_ (.A(_0990_),
    .X(net151));
 sky130_fd_sc_hd__and2_1 _3870_ (.A(\core_1.ew_data[7] ),
    .B(net157),
    .X(_0991_));
 sky130_fd_sc_hd__clkbuf_1 _3871_ (.A(_0991_),
    .X(net152));
 sky130_fd_sc_hd__mux2_1 _3872_ (.A0(\core_1.ew_data[0] ),
    .A1(\core_1.ew_data[8] ),
    .S(net157),
    .X(_0992_));
 sky130_fd_sc_hd__clkbuf_1 _3873_ (.A(_0992_),
    .X(net153));
 sky130_fd_sc_hd__mux2_1 _3874_ (.A0(\core_1.ew_data[1] ),
    .A1(\core_1.ew_data[9] ),
    .S(_0983_),
    .X(_0993_));
 sky130_fd_sc_hd__clkbuf_1 _3875_ (.A(_0993_),
    .X(net154));
 sky130_fd_sc_hd__mux2_1 _3876_ (.A0(\core_1.ew_data[2] ),
    .A1(\core_1.ew_data[10] ),
    .S(_0983_),
    .X(_0994_));
 sky130_fd_sc_hd__clkbuf_1 _3877_ (.A(_0994_),
    .X(net140));
 sky130_fd_sc_hd__mux2_1 _3878_ (.A0(\core_1.ew_data[3] ),
    .A1(\core_1.ew_data[11] ),
    .S(_0983_),
    .X(_0995_));
 sky130_fd_sc_hd__clkbuf_1 _3879_ (.A(_0995_),
    .X(net141));
 sky130_fd_sc_hd__mux2_1 _3880_ (.A0(\core_1.ew_data[4] ),
    .A1(\core_1.ew_data[12] ),
    .S(_0983_),
    .X(_0996_));
 sky130_fd_sc_hd__clkbuf_1 _3881_ (.A(_0996_),
    .X(net142));
 sky130_fd_sc_hd__mux2_1 _3882_ (.A0(\core_1.ew_data[5] ),
    .A1(\core_1.ew_data[13] ),
    .S(_0983_),
    .X(_0997_));
 sky130_fd_sc_hd__clkbuf_1 _3883_ (.A(_0997_),
    .X(net143));
 sky130_fd_sc_hd__mux2_1 _3884_ (.A0(\core_1.ew_data[6] ),
    .A1(\core_1.ew_data[14] ),
    .S(_0983_),
    .X(_0998_));
 sky130_fd_sc_hd__clkbuf_1 _3885_ (.A(_0998_),
    .X(net144));
 sky130_fd_sc_hd__mux2_1 _3886_ (.A0(\core_1.ew_data[7] ),
    .A1(\core_1.ew_data[15] ),
    .S(_0983_),
    .X(_0999_));
 sky130_fd_sc_hd__clkbuf_1 _3887_ (.A(_0999_),
    .X(net145));
 sky130_fd_sc_hd__or2b_2 _3888_ (.A(\core_1.ew_addr[0] ),
    .B_N(\core_1.ew_mem_width ),
    .X(_1000_));
 sky130_fd_sc_hd__clkbuf_1 _3889_ (.A(_1000_),
    .X(net158));
 sky130_fd_sc_hd__inv_2 _3890_ (.A(net17),
    .Y(net160));
 sky130_fd_sc_hd__nor2_2 _3891_ (.A(\core_1.decode.i_flush ),
    .B(\core_1.fetch.flush_event_invalidate ),
    .Y(_1001_));
 sky130_fd_sc_hd__o211ai_4 _3892_ (.A1(_0664_),
    .A2(net70),
    .B1(_0737_),
    .C1(_1001_),
    .Y(_1002_));
 sky130_fd_sc_hd__inv_2 _3893_ (.A(_1002_),
    .Y(\core_1.fetch.submitable ));
 sky130_fd_sc_hd__and2_1 _3894_ (.A(net155),
    .B(\core_1.ew_addr_high[0] ),
    .X(_1003_));
 sky130_fd_sc_hd__clkbuf_1 _3895_ (.A(_1003_),
    .X(net122));
 sky130_fd_sc_hd__nor3_1 _3896_ (.A(\core_1.decode.i_flush ),
    .B(_0688_),
    .C(_0689_),
    .Y(_1004_));
 sky130_fd_sc_hd__nor3b_2 _3897_ (.A(_0724_),
    .B(_0732_),
    .C_N(_1004_),
    .Y(_1005_));
 sky130_fd_sc_hd__clkbuf_4 _3898_ (.A(_1005_),
    .X(_1006_));
 sky130_fd_sc_hd__clkbuf_4 _3899_ (.A(_1006_),
    .X(_1007_));
 sky130_fd_sc_hd__inv_2 _3900_ (.A(net211),
    .Y(_1008_));
 sky130_fd_sc_hd__clkbuf_4 _3901_ (.A(_1008_),
    .X(_1009_));
 sky130_fd_sc_hd__inv_2 _3902_ (.A(net186),
    .Y(_1010_));
 sky130_fd_sc_hd__nor4_4 _3903_ (.A(net189),
    .B(net188),
    .C(net191),
    .D(net190),
    .Y(_1011_));
 sky130_fd_sc_hd__and3b_1 _3904_ (.A_N(net187),
    .B(_1010_),
    .C(_1011_),
    .X(_1012_));
 sky130_fd_sc_hd__nor3_4 _3905_ (.A(net193),
    .B(net180),
    .C(net179),
    .Y(_1013_));
 sky130_fd_sc_hd__nor4_4 _3906_ (.A(net182),
    .B(net181),
    .C(net184),
    .D(net183),
    .Y(_1014_));
 sky130_fd_sc_hd__and4bb_1 _3907_ (.A_N(net185),
    .B_N(net192),
    .C(_1013_),
    .D(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__clkbuf_2 _3908_ (.A(_1015_),
    .X(_1016_));
 sky130_fd_sc_hd__and3_2 _3909_ (.A(_1009_),
    .B(_1012_),
    .C(_1016_),
    .X(_1017_));
 sky130_fd_sc_hd__clkbuf_4 _3910_ (.A(\core_1.dec_sreg_irt ),
    .X(_1018_));
 sky130_fd_sc_hd__buf_4 _3911_ (.A(_1018_),
    .X(_1019_));
 sky130_fd_sc_hd__a21o_1 _3912_ (.A1(\core_1.dec_sreg_store ),
    .A2(_1017_),
    .B1(_1019_),
    .X(_1020_));
 sky130_fd_sc_hd__inv_2 _3913_ (.A(\core_1.dec_jump_cond_code[1] ),
    .Y(_1021_));
 sky130_fd_sc_hd__inv_2 _3914_ (.A(\core_1.dec_jump_cond_code[0] ),
    .Y(_1022_));
 sky130_fd_sc_hd__a211oi_1 _3915_ (.A1(\core_1.execute.alu_flag_reg.o_d[0] ),
    .A2(_1022_),
    .B1(_1021_),
    .C1(\core_1.execute.alu_flag_reg.o_d[1] ),
    .Y(_1023_));
 sky130_fd_sc_hd__a31o_1 _3916_ (.A1(\core_1.execute.alu_flag_reg.o_d[4] ),
    .A2(\core_1.dec_jump_cond_code[0] ),
    .A3(_1021_),
    .B1(_1023_),
    .X(_1024_));
 sky130_fd_sc_hd__nor2_1 _3917_ (.A(\core_1.dec_jump_cond_code[0] ),
    .B(\core_1.dec_jump_cond_code[1] ),
    .Y(_1025_));
 sky130_fd_sc_hd__o21a_1 _3918_ (.A1(\core_1.execute.alu_flag_reg.o_d[1] ),
    .A2(\core_1.execute.alu_flag_reg.o_d[0] ),
    .B1(_1025_),
    .X(_1026_));
 sky130_fd_sc_hd__mux2_1 _3919_ (.A0(_1024_),
    .A1(_1026_),
    .S(\core_1.dec_jump_cond_code[2] ),
    .X(_1027_));
 sky130_fd_sc_hd__nand2_1 _3920_ (.A(\core_1.dec_jump_cond_code[3] ),
    .B(_1027_),
    .Y(_1028_));
 sky130_fd_sc_hd__mux2_1 _3921_ (.A0(\core_1.execute.alu_flag_reg.o_d[1] ),
    .A1(\core_1.execute.alu_flag_reg.o_d[2] ),
    .S(\core_1.dec_jump_cond_code[1] ),
    .X(_1029_));
 sky130_fd_sc_hd__a31o_1 _3922_ (.A1(\core_1.execute.alu_flag_reg.o_d[0] ),
    .A2(_1022_),
    .A3(\core_1.dec_jump_cond_code[1] ),
    .B1(\core_1.dec_jump_cond_code[2] ),
    .X(_1030_));
 sky130_fd_sc_hd__a21oi_1 _3923_ (.A1(\core_1.dec_jump_cond_code[0] ),
    .A2(_1029_),
    .B1(_1030_),
    .Y(_1031_));
 sky130_fd_sc_hd__mux2_1 _3924_ (.A0(\core_1.execute.alu_flag_reg.o_d[2] ),
    .A1(\core_1.execute.alu_flag_reg.o_d[0] ),
    .S(\core_1.dec_jump_cond_code[0] ),
    .X(_1032_));
 sky130_fd_sc_hd__o21ai_1 _3925_ (.A1(\core_1.execute.alu_flag_reg.o_d[2] ),
    .A2(\core_1.execute.alu_flag_reg.o_d[0] ),
    .B1(_1021_),
    .Y(_1033_));
 sky130_fd_sc_hd__o221a_1 _3926_ (.A1(_1021_),
    .A2(_1032_),
    .B1(_1033_),
    .B2(_1022_),
    .C1(\core_1.dec_jump_cond_code[2] ),
    .X(_1034_));
 sky130_fd_sc_hd__inv_2 _3927_ (.A(\core_1.execute.alu_flag_reg.o_d[3] ),
    .Y(_1035_));
 sky130_fd_sc_hd__o21a_1 _3928_ (.A1(_1035_),
    .A2(\core_1.dec_jump_cond_code[2] ),
    .B1(\core_1.dec_jump_cond_code[3] ),
    .X(_1036_));
 sky130_fd_sc_hd__o21ai_1 _3929_ (.A1(\core_1.execute.alu_flag_reg.o_d[2] ),
    .A2(\core_1.execute.alu_flag_reg.o_d[0] ),
    .B1(\core_1.dec_jump_cond_code[2] ),
    .Y(_1037_));
 sky130_fd_sc_hd__nand2_1 _3930_ (.A(_1025_),
    .B(_1037_),
    .Y(_1038_));
 sky130_fd_sc_hd__o32a_1 _3931_ (.A1(\core_1.dec_jump_cond_code[3] ),
    .A2(_1031_),
    .A3(_1034_),
    .B1(_1036_),
    .B2(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__a21boi_1 _3932_ (.A1(_1028_),
    .A2(_1039_),
    .B1_N(\core_1.dec_jump_cond_code[4] ),
    .Y(_1040_));
 sky130_fd_sc_hd__and3_1 _3933_ (.A(\core_1.dec_jump_cond_code[4] ),
    .B(_1028_),
    .C(_1039_),
    .X(_1041_));
 sky130_fd_sc_hd__mux2_1 _3934_ (.A0(_1040_),
    .A1(_1041_),
    .S(\core_1.de_jmp_pred ),
    .X(_1042_));
 sky130_fd_sc_hd__or4b_4 _3935_ (.A(_0724_),
    .B(_0726_),
    .C(_0731_),
    .D_N(_1004_),
    .X(_1043_));
 sky130_fd_sc_hd__nor2_1 _3936_ (.A(\core_1.dec_jump_cond_code[4] ),
    .B(_1020_),
    .Y(_1044_));
 sky130_fd_sc_hd__nor2_2 _3937_ (.A(_1043_),
    .B(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__nand2_1 _3938_ (.A(\core_1.execute.sreg_jtr_buff.o_d[0] ),
    .B(_1045_),
    .Y(_1046_));
 sky130_fd_sc_hd__and2b_2 _3939_ (.A_N(_1044_),
    .B(_1005_),
    .X(_1047_));
 sky130_fd_sc_hd__nor2_1 _3940_ (.A(_0667_),
    .B(_1047_),
    .Y(_1048_));
 sky130_fd_sc_hd__a21oi_1 _3941_ (.A1(\core_1.execute.sreg_jtr_buff.o_d[0] ),
    .A2(_0668_),
    .B1(_1048_),
    .Y(_1049_));
 sky130_fd_sc_hd__and3_1 _3942_ (.A(net192),
    .B(\core_1.dec_sreg_store ),
    .C(_1013_),
    .X(_1050_));
 sky130_fd_sc_hd__and4_1 _3943_ (.A(_1005_),
    .B(_1011_),
    .C(_1014_),
    .D(_1050_),
    .X(_1051_));
 sky130_fd_sc_hd__o21ai_1 _3944_ (.A1(_1049_),
    .A2(_1051_),
    .B1(net106),
    .Y(_1052_));
 sky130_fd_sc_hd__o211a_2 _3945_ (.A1(net106),
    .A2(_1046_),
    .B1(_1052_),
    .C1(_0687_),
    .X(_1053_));
 sky130_fd_sc_hd__or3b_1 _3946_ (.A(_1020_),
    .B(_1042_),
    .C_N(_1053_),
    .X(_1054_));
 sky130_fd_sc_hd__a21o_1 _3947_ (.A1(_1007_),
    .A2(_1054_),
    .B1(_0688_),
    .X(_0013_));
 sky130_fd_sc_hd__clkbuf_4 _3948_ (.A(_0659_),
    .X(_1055_));
 sky130_fd_sc_hd__buf_6 _3949_ (.A(_1055_),
    .X(_1056_));
 sky130_fd_sc_hd__nor2_1 _3950_ (.A(_1056_),
    .B(_1053_),
    .Y(_0014_));
 sky130_fd_sc_hd__buf_6 _3951_ (.A(\core_1.dec_sreg_store ),
    .X(_1057_));
 sky130_fd_sc_hd__and3_1 _3952_ (.A(\core_1.execute.sreg_priv_control.o_d[0] ),
    .B(_1057_),
    .C(_0734_),
    .X(_1058_));
 sky130_fd_sc_hd__clkbuf_1 _3953_ (.A(_1058_),
    .X(net210));
 sky130_fd_sc_hd__buf_4 _3954_ (.A(_0812_),
    .X(_0015_));
 sky130_fd_sc_hd__buf_4 _3955_ (.A(_0811_),
    .X(_1059_));
 sky130_fd_sc_hd__mux2_1 _3956_ (.A0(net178),
    .A1(\core_1.decode.i_imm_pass[0] ),
    .S(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__clkbuf_1 _3957_ (.A(_1060_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _3958_ (.A0(net185),
    .A1(\core_1.decode.i_imm_pass[1] ),
    .S(_1059_),
    .X(_1061_));
 sky130_fd_sc_hd__clkbuf_1 _3959_ (.A(_1061_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _3960_ (.A0(net186),
    .A1(\core_1.decode.i_imm_pass[2] ),
    .S(_1059_),
    .X(_1062_));
 sky130_fd_sc_hd__clkbuf_1 _3961_ (.A(_1062_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _3962_ (.A0(net187),
    .A1(\core_1.decode.i_imm_pass[3] ),
    .S(_1059_),
    .X(_1063_));
 sky130_fd_sc_hd__clkbuf_1 _3963_ (.A(_1063_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _3964_ (.A0(net188),
    .A1(\core_1.decode.i_imm_pass[4] ),
    .S(_1059_),
    .X(_1064_));
 sky130_fd_sc_hd__clkbuf_1 _3965_ (.A(_1064_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _3966_ (.A0(net189),
    .A1(\core_1.decode.i_imm_pass[5] ),
    .S(_1059_),
    .X(_1065_));
 sky130_fd_sc_hd__clkbuf_1 _3967_ (.A(_1065_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _3968_ (.A0(net190),
    .A1(\core_1.decode.i_imm_pass[6] ),
    .S(_1059_),
    .X(_1066_));
 sky130_fd_sc_hd__clkbuf_1 _3969_ (.A(_1066_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _3970_ (.A0(net191),
    .A1(\core_1.decode.i_imm_pass[7] ),
    .S(_1059_),
    .X(_1067_));
 sky130_fd_sc_hd__clkbuf_1 _3971_ (.A(_1067_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _3972_ (.A0(net192),
    .A1(\core_1.decode.i_imm_pass[8] ),
    .S(_1059_),
    .X(_1068_));
 sky130_fd_sc_hd__clkbuf_1 _3973_ (.A(_1068_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _3974_ (.A0(net193),
    .A1(\core_1.decode.i_imm_pass[9] ),
    .S(_1059_),
    .X(_1069_));
 sky130_fd_sc_hd__clkbuf_1 _3975_ (.A(_1069_),
    .X(_0025_));
 sky130_fd_sc_hd__buf_8 _3976_ (.A(_0811_),
    .X(_1070_));
 sky130_fd_sc_hd__mux2_1 _3977_ (.A0(net179),
    .A1(\core_1.decode.i_imm_pass[10] ),
    .S(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__clkbuf_1 _3978_ (.A(_1071_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _3979_ (.A0(net180),
    .A1(\core_1.decode.i_imm_pass[11] ),
    .S(_1070_),
    .X(_1072_));
 sky130_fd_sc_hd__clkbuf_1 _3980_ (.A(_1072_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _3981_ (.A0(net181),
    .A1(\core_1.decode.i_imm_pass[12] ),
    .S(_1070_),
    .X(_1073_));
 sky130_fd_sc_hd__clkbuf_1 _3982_ (.A(_1073_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _3983_ (.A0(net182),
    .A1(\core_1.decode.i_imm_pass[13] ),
    .S(_1070_),
    .X(_1074_));
 sky130_fd_sc_hd__clkbuf_1 _3984_ (.A(_1074_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _3985_ (.A0(net183),
    .A1(\core_1.decode.i_imm_pass[14] ),
    .S(_1070_),
    .X(_1075_));
 sky130_fd_sc_hd__clkbuf_1 _3986_ (.A(_1075_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _3987_ (.A0(net184),
    .A1(\core_1.decode.i_imm_pass[15] ),
    .S(_1070_),
    .X(_1076_));
 sky130_fd_sc_hd__clkbuf_1 _3988_ (.A(_1076_),
    .X(_0031_));
 sky130_fd_sc_hd__or3_1 _3989_ (.A(_0810_),
    .B(_0819_),
    .C(_0852_),
    .X(_1077_));
 sky130_fd_sc_hd__a211o_1 _3990_ (.A1(_0847_),
    .A2(_0852_),
    .B1(_0803_),
    .C1(_0810_),
    .X(_1078_));
 sky130_fd_sc_hd__o211a_1 _3991_ (.A1(\core_1.dec_pc_inc ),
    .A2(_0812_),
    .B1(_1077_),
    .C1(_1078_),
    .X(_0032_));
 sky130_fd_sc_hd__buf_4 _3992_ (.A(\core_1.dec_r_bus_imm ),
    .X(_1079_));
 sky130_fd_sc_hd__o21bai_1 _3993_ (.A1(_0818_),
    .A2(_0847_),
    .B1_N(_0795_),
    .Y(_1080_));
 sky130_fd_sc_hd__or3_1 _3994_ (.A(_0801_),
    .B(_0855_),
    .C(_1080_),
    .X(_1081_));
 sky130_fd_sc_hd__a21oi_1 _3995_ (.A1(_0800_),
    .A2(_0824_),
    .B1(_0803_),
    .Y(_1082_));
 sky130_fd_sc_hd__or3_1 _3996_ (.A(_0807_),
    .B(_1081_),
    .C(_1082_),
    .X(_1083_));
 sky130_fd_sc_hd__a21oi_1 _3997_ (.A1(_0790_),
    .A2(_0842_),
    .B1(_0819_),
    .Y(_1084_));
 sky130_fd_sc_hd__o21a_1 _3998_ (.A1(\core_1.decode.i_instr_l[0] ),
    .A2(_0787_),
    .B1(_0805_),
    .X(_1085_));
 sky130_fd_sc_hd__nor2_1 _3999_ (.A(_0799_),
    .B(_1085_),
    .Y(_1086_));
 sky130_fd_sc_hd__o211a_1 _4000_ (.A1(_0782_),
    .A2(_0828_),
    .B1(_0842_),
    .C1(_0789_),
    .X(_1087_));
 sky130_fd_sc_hd__a31o_1 _4001_ (.A1(_0850_),
    .A2(_0852_),
    .A3(_1087_),
    .B1(_0803_),
    .X(_1088_));
 sky130_fd_sc_hd__or4b_1 _4002_ (.A(_1083_),
    .B(_1084_),
    .C(_1086_),
    .D_N(_1088_),
    .X(_1089_));
 sky130_fd_sc_hd__mux2_1 _4003_ (.A0(_1079_),
    .A1(_1089_),
    .S(_1070_),
    .X(_1090_));
 sky130_fd_sc_hd__clkbuf_1 _4004_ (.A(_1090_),
    .X(_0033_));
 sky130_fd_sc_hd__o21bai_1 _4005_ (.A1(_0819_),
    .A2(_0841_),
    .B1_N(_0844_),
    .Y(_1091_));
 sky130_fd_sc_hd__a21oi_1 _4006_ (.A1(_0805_),
    .A2(_0787_),
    .B1(_0799_),
    .Y(_1092_));
 sky130_fd_sc_hd__or2_1 _4007_ (.A(_0792_),
    .B(_1092_),
    .X(_1093_));
 sky130_fd_sc_hd__and2_1 _4008_ (.A(_0805_),
    .B(_0849_),
    .X(_1094_));
 sky130_fd_sc_hd__a31o_1 _4009_ (.A1(_0790_),
    .A2(_0824_),
    .A3(_1094_),
    .B1(_0818_),
    .X(_1095_));
 sky130_fd_sc_hd__or4b_1 _4010_ (.A(_0864_),
    .B(_1091_),
    .C(_1093_),
    .D_N(_1095_),
    .X(_1096_));
 sky130_fd_sc_hd__mux2_1 _4011_ (.A0(\core_1.dec_alu_flags_ie ),
    .A1(_1096_),
    .S(_1070_),
    .X(_1097_));
 sky130_fd_sc_hd__clkbuf_1 _4012_ (.A(_1097_),
    .X(_0034_));
 sky130_fd_sc_hd__and3_1 _4013_ (.A(\core_1.decode.i_instr_l[0] ),
    .B(_0796_),
    .C(_0840_),
    .X(_1098_));
 sky130_fd_sc_hd__mux2_1 _4014_ (.A0(\core_1.dec_alu_carry_en ),
    .A1(_1098_),
    .S(_1070_),
    .X(_1099_));
 sky130_fd_sc_hd__clkbuf_1 _4015_ (.A(_1099_),
    .X(_0035_));
 sky130_fd_sc_hd__nor2_1 _4016_ (.A(\core_1.decode.i_instr_l[3] ),
    .B(\core_1.decode.i_instr_l[2] ),
    .Y(_1100_));
 sky130_fd_sc_hd__a311o_1 _4017_ (.A1(\core_1.decode.i_instr_l[0] ),
    .A2(_0796_),
    .A3(_1100_),
    .B1(_0795_),
    .C1(_0837_),
    .X(_1101_));
 sky130_fd_sc_hd__a211o_1 _4018_ (.A1(_0782_),
    .A2(_0806_),
    .B1(_1093_),
    .C1(_1101_),
    .X(_1102_));
 sky130_fd_sc_hd__a21oi_1 _4019_ (.A1(_0790_),
    .A2(_0828_),
    .B1(_0819_),
    .Y(_1103_));
 sky130_fd_sc_hd__or4_4 _4020_ (.A(_1091_),
    .B(_1096_),
    .C(_1102_),
    .D(_1103_),
    .X(_1104_));
 sky130_fd_sc_hd__a21o_2 _4021_ (.A1(\core_1.decode.i_instr_l[0] ),
    .A2(_0806_),
    .B1(_0802_),
    .X(_1105_));
 sky130_fd_sc_hd__a221o_1 _4022_ (.A1(\core_1.decode.i_instr_l[10] ),
    .A2(_1104_),
    .B1(_1105_),
    .B2(\core_1.decode.i_instr_l[13] ),
    .C1(_0815_),
    .X(_1106_));
 sky130_fd_sc_hd__o21a_1 _4023_ (.A1(_0701_),
    .A2(_0015_),
    .B1(_1106_),
    .X(_0036_));
 sky130_fd_sc_hd__a221o_1 _4024_ (.A1(\core_1.decode.i_instr_l[11] ),
    .A2(_1104_),
    .B1(_1105_),
    .B2(\core_1.decode.i_instr_l[14] ),
    .C1(_0815_),
    .X(_1107_));
 sky130_fd_sc_hd__o21a_1 _4025_ (.A1(_0695_),
    .A2(_0015_),
    .B1(_1107_),
    .X(_0037_));
 sky130_fd_sc_hd__a221o_1 _4026_ (.A1(\core_1.decode.i_instr_l[12] ),
    .A2(_1104_),
    .B1(_1105_),
    .B2(\core_1.decode.i_instr_l[15] ),
    .C1(_0815_),
    .X(_1108_));
 sky130_fd_sc_hd__o21a_1 _4027_ (.A1(_0717_),
    .A2(_0015_),
    .B1(_1108_),
    .X(_0038_));
 sky130_fd_sc_hd__nor2_1 _4028_ (.A(_0794_),
    .B(_0818_),
    .Y(_1109_));
 sky130_fd_sc_hd__a21o_1 _4029_ (.A1(_0783_),
    .A2(_0797_),
    .B1(_0781_),
    .X(_1110_));
 sky130_fd_sc_hd__o21ai_1 _4030_ (.A1(_0803_),
    .A2(_1110_),
    .B1(_1095_),
    .Y(_1111_));
 sky130_fd_sc_hd__or4_1 _4031_ (.A(_0851_),
    .B(_1080_),
    .C(_1109_),
    .D(_1111_),
    .X(_1112_));
 sky130_fd_sc_hd__a32o_1 _4032_ (.A1(_0828_),
    .A2(_1094_),
    .A3(_1110_),
    .B1(_0836_),
    .B2(_0819_),
    .X(_1113_));
 sky130_fd_sc_hd__a22oi_2 _4033_ (.A1(_0799_),
    .A2(_0819_),
    .B1(_0833_),
    .B2(_1113_),
    .Y(_1114_));
 sky130_fd_sc_hd__o31a_1 _4034_ (.A1(_1102_),
    .A2(_1112_),
    .A3(_1114_),
    .B1(_0811_),
    .X(_1115_));
 sky130_fd_sc_hd__and2b_1 _4035_ (.A_N(\core_1.decode.i_instr_l[9] ),
    .B(_1115_),
    .X(_1116_));
 sky130_fd_sc_hd__and2b_1 _4036_ (.A_N(\core_1.decode.i_instr_l[7] ),
    .B(_1116_),
    .X(_1117_));
 sky130_fd_sc_hd__inv_2 _4037_ (.A(\core_1.decode.i_instr_l[8] ),
    .Y(_1118_));
 sky130_fd_sc_hd__a22o_1 _4038_ (.A1(\core_1.dec_rf_ie[0] ),
    .A2(_0816_),
    .B1(_1117_),
    .B2(_1118_),
    .X(_0039_));
 sky130_fd_sc_hd__a32o_1 _4039_ (.A1(_1118_),
    .A2(\core_1.decode.i_instr_l[7] ),
    .A3(_1116_),
    .B1(_0830_),
    .B2(\core_1.dec_rf_ie[1] ),
    .X(_0040_));
 sky130_fd_sc_hd__a22o_1 _4040_ (.A1(\core_1.dec_rf_ie[2] ),
    .A2(_0830_),
    .B1(_1117_),
    .B2(\core_1.decode.i_instr_l[8] ),
    .X(_0041_));
 sky130_fd_sc_hd__a32o_1 _4041_ (.A1(\core_1.decode.i_instr_l[8] ),
    .A2(\core_1.decode.i_instr_l[7] ),
    .A3(_1116_),
    .B1(_0830_),
    .B2(\core_1.dec_rf_ie[3] ),
    .X(_0042_));
 sky130_fd_sc_hd__and2_1 _4042_ (.A(\core_1.decode.i_instr_l[9] ),
    .B(_1115_),
    .X(_1119_));
 sky130_fd_sc_hd__or2b_1 _4043_ (.A(\core_1.decode.i_instr_l[7] ),
    .B_N(_1119_),
    .X(_1120_));
 sky130_fd_sc_hd__a2bb2o_1 _4044_ (.A1_N(\core_1.decode.i_instr_l[8] ),
    .A2_N(_1120_),
    .B1(_0816_),
    .B2(\core_1.dec_rf_ie[4] ),
    .X(_0043_));
 sky130_fd_sc_hd__a32o_1 _4045_ (.A1(_1118_),
    .A2(\core_1.decode.i_instr_l[7] ),
    .A3(_1119_),
    .B1(_0830_),
    .B2(\core_1.dec_rf_ie[5] ),
    .X(_0044_));
 sky130_fd_sc_hd__a2bb2o_1 _4046_ (.A1_N(_1118_),
    .A2_N(_1120_),
    .B1(_0816_),
    .B2(\core_1.dec_rf_ie[6] ),
    .X(_0045_));
 sky130_fd_sc_hd__a32o_1 _4047_ (.A1(\core_1.decode.i_instr_l[8] ),
    .A2(\core_1.decode.i_instr_l[7] ),
    .A3(_1119_),
    .B1(_0815_),
    .B2(\core_1.dec_rf_ie[7] ),
    .X(_0046_));
 sky130_fd_sc_hd__a211o_1 _4048_ (.A1(_0840_),
    .A2(_0788_),
    .B1(_0866_),
    .C1(_0861_),
    .X(_1121_));
 sky130_fd_sc_hd__a21o_2 _4049_ (.A1(_0796_),
    .A2(_1121_),
    .B1(_1114_),
    .X(_1122_));
 sky130_fd_sc_hd__or2_1 _4050_ (.A(_0856_),
    .B(_1105_),
    .X(_1123_));
 sky130_fd_sc_hd__nor2_1 _4051_ (.A(_0819_),
    .B(_0854_),
    .Y(_1124_));
 sky130_fd_sc_hd__or2_2 _4052_ (.A(_1123_),
    .B(_1124_),
    .X(_1125_));
 sky130_fd_sc_hd__a221o_1 _4053_ (.A1(\core_1.decode.i_instr_l[13] ),
    .A2(_1122_),
    .B1(_1125_),
    .B2(\core_1.decode.i_instr_l[10] ),
    .C1(_0815_),
    .X(_1126_));
 sky130_fd_sc_hd__o21a_1 _4054_ (.A1(_0558_),
    .A2(_0015_),
    .B1(_1126_),
    .X(_0047_));
 sky130_fd_sc_hd__a221o_1 _4055_ (.A1(\core_1.decode.i_instr_l[14] ),
    .A2(_1122_),
    .B1(_1125_),
    .B2(\core_1.decode.i_instr_l[11] ),
    .C1(_0815_),
    .X(_1127_));
 sky130_fd_sc_hd__o21a_1 _4056_ (.A1(_0555_),
    .A2(_0015_),
    .B1(_1127_),
    .X(_0048_));
 sky130_fd_sc_hd__a221o_1 _4057_ (.A1(\core_1.decode.i_instr_l[15] ),
    .A2(_1122_),
    .B1(_1125_),
    .B2(\core_1.decode.i_instr_l[12] ),
    .C1(_0815_),
    .X(_1128_));
 sky130_fd_sc_hd__o21a_1 _4058_ (.A1(_0534_),
    .A2(_0015_),
    .B1(_1128_),
    .X(_0049_));
 sky130_fd_sc_hd__nor3_2 _4059_ (.A(_0803_),
    .B(_0810_),
    .C(_0852_),
    .Y(_1129_));
 sky130_fd_sc_hd__a22o_1 _4060_ (.A1(\core_1.dec_jump_cond_code[0] ),
    .A2(_0830_),
    .B1(_1129_),
    .B2(\core_1.decode.i_instr_l[7] ),
    .X(_0050_));
 sky130_fd_sc_hd__a22o_1 _4061_ (.A1(\core_1.dec_jump_cond_code[1] ),
    .A2(_0830_),
    .B1(_1129_),
    .B2(\core_1.decode.i_instr_l[8] ),
    .X(_0051_));
 sky130_fd_sc_hd__a22o_1 _4062_ (.A1(\core_1.dec_jump_cond_code[2] ),
    .A2(_0830_),
    .B1(_1129_),
    .B2(\core_1.decode.i_instr_l[9] ),
    .X(_0052_));
 sky130_fd_sc_hd__a22o_1 _4063_ (.A1(\core_1.dec_jump_cond_code[3] ),
    .A2(_0830_),
    .B1(_1129_),
    .B2(\core_1.decode.i_instr_l[10] ),
    .X(_0053_));
 sky130_fd_sc_hd__a21bo_1 _4064_ (.A1(\core_1.dec_jump_cond_code[4] ),
    .A2(_0816_),
    .B1_N(_1078_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _4065_ (.A0(\core_1.de_jmp_pred ),
    .A1(\core_1.decode.i_jmp_pred_pass ),
    .S(_1070_),
    .X(_1130_));
 sky130_fd_sc_hd__clkbuf_1 _4066_ (.A(_1130_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _4067_ (.A0(\core_1.dec_mem_access ),
    .A1(_1083_),
    .S(_0811_),
    .X(_1131_));
 sky130_fd_sc_hd__clkbuf_1 _4068_ (.A(_1131_),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _4069_ (.A0(\core_1.dec_mem_we ),
    .A1(_1123_),
    .S(_0811_),
    .X(_1132_));
 sky130_fd_sc_hd__clkbuf_1 _4070_ (.A(_1132_),
    .X(_0057_));
 sky130_fd_sc_hd__or3_1 _4071_ (.A(_0810_),
    .B(_1104_),
    .C(_1105_),
    .X(_1133_));
 sky130_fd_sc_hd__o21a_1 _4072_ (.A1(\core_1.dec_used_operands[0] ),
    .A2(_0015_),
    .B1(_1133_),
    .X(_0058_));
 sky130_fd_sc_hd__or3_1 _4073_ (.A(_0810_),
    .B(_1122_),
    .C(_1125_),
    .X(_1134_));
 sky130_fd_sc_hd__o21a_1 _4074_ (.A1(\core_1.dec_used_operands[1] ),
    .A2(_0015_),
    .B1(_1134_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _4075_ (.A0(\core_1.dec_sreg_load ),
    .A1(_1109_),
    .S(_0811_),
    .X(_1135_));
 sky130_fd_sc_hd__clkbuf_1 _4076_ (.A(_1135_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _4077_ (.A0(_1057_),
    .A1(_1124_),
    .S(_0811_),
    .X(_1136_));
 sky130_fd_sc_hd__clkbuf_1 _4078_ (.A(_1136_),
    .X(_0061_));
 sky130_fd_sc_hd__clkinv_2 _4079_ (.A(\core_1.dec_sreg_jal_over ),
    .Y(_1137_));
 sky130_fd_sc_hd__buf_4 _4080_ (.A(_1137_),
    .X(_1138_));
 sky130_fd_sc_hd__or3_1 _4081_ (.A(_0803_),
    .B(_0810_),
    .C(_0847_),
    .X(_1139_));
 sky130_fd_sc_hd__o21ai_1 _4082_ (.A1(_1138_),
    .A2(_0812_),
    .B1(_1139_),
    .Y(_0062_));
 sky130_fd_sc_hd__clkinv_2 _4083_ (.A(\core_1.dec_sreg_irt ),
    .Y(_1140_));
 sky130_fd_sc_hd__buf_4 _4084_ (.A(_1140_),
    .X(_1141_));
 sky130_fd_sc_hd__o21ai_1 _4085_ (.A1(_1141_),
    .A2(_0812_),
    .B1(_1077_),
    .Y(_0063_));
 sky130_fd_sc_hd__inv_2 _4086_ (.A(_0800_),
    .Y(_1142_));
 sky130_fd_sc_hd__a22o_1 _4087_ (.A1(\core_1.dec_sys ),
    .A2(_0830_),
    .B1(_1142_),
    .B2(_0820_),
    .X(_0064_));
 sky130_fd_sc_hd__a211o_1 _4088_ (.A1(\core_1.decode.i_instr_l[1] ),
    .A2(_0806_),
    .B1(_1081_),
    .C1(_0815_),
    .X(_1143_));
 sky130_fd_sc_hd__o21a_1 _4089_ (.A1(\core_1.dec_mem_width ),
    .A2(_0015_),
    .B1(_1143_),
    .X(_0065_));
 sky130_fd_sc_hd__o211a_1 _4090_ (.A1(\core_1.decode.input_valid ),
    .A2(\core_1.decode.i_submit ),
    .B1(_0736_),
    .C1(_0809_),
    .X(_0066_));
 sky130_fd_sc_hd__and3_2 _4091_ (.A(net211),
    .B(_1012_),
    .C(_1016_),
    .X(_1144_));
 sky130_fd_sc_hd__buf_4 _4092_ (.A(_1144_),
    .X(_1145_));
 sky130_fd_sc_hd__clkbuf_4 _4093_ (.A(_1019_),
    .X(_1146_));
 sky130_fd_sc_hd__a31o_1 _4094_ (.A1(\core_1.execute.sreg_priv_control.o_d[0] ),
    .A2(\core_1.dec_sreg_store ),
    .A3(_1145_),
    .B1(_1146_),
    .X(_1147_));
 sky130_fd_sc_hd__nand3_2 _4095_ (.A(_1141_),
    .B(_1005_),
    .C(_1147_),
    .Y(_1148_));
 sky130_fd_sc_hd__and2_1 _4096_ (.A(_0668_),
    .B(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__clkbuf_4 _4097_ (.A(_1149_),
    .X(_1150_));
 sky130_fd_sc_hd__or2_1 _4098_ (.A(_0659_),
    .B(_0667_),
    .X(_1151_));
 sky130_fd_sc_hd__clkbuf_4 _4099_ (.A(_1148_),
    .X(_1152_));
 sky130_fd_sc_hd__nor2_1 _4100_ (.A(_0658_),
    .B(_1152_),
    .Y(_1153_));
 sky130_fd_sc_hd__a211o_1 _4101_ (.A1(\core_1.execute.sreg_priv_control.o_d[0] ),
    .A2(_1150_),
    .B1(_1151_),
    .C1(_1153_),
    .X(_0067_));
 sky130_fd_sc_hd__inv_2 _4102_ (.A(net71),
    .Y(_1154_));
 sky130_fd_sc_hd__buf_6 _4103_ (.A(_1154_),
    .X(_1155_));
 sky130_fd_sc_hd__clkbuf_4 _4104_ (.A(_1155_),
    .X(_1156_));
 sky130_fd_sc_hd__a2bb2o_1 _4105_ (.A1_N(_0650_),
    .A2_N(_1152_),
    .B1(_1150_),
    .B2(\core_1.execute.sreg_data_page ),
    .X(_1157_));
 sky130_fd_sc_hd__and2_1 _4106_ (.A(_1156_),
    .B(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__clkbuf_1 _4107_ (.A(_1158_),
    .X(_0068_));
 sky130_fd_sc_hd__a2bb2o_1 _4108_ (.A1_N(_0635_),
    .A2_N(_1152_),
    .B1(_1150_),
    .B2(\core_1.execute.sreg_long_ptr_en ),
    .X(_1159_));
 sky130_fd_sc_hd__and2_1 _4109_ (.A(_1156_),
    .B(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__clkbuf_1 _4110_ (.A(_1160_),
    .X(_0069_));
 sky130_fd_sc_hd__a2bb2o_1 _4111_ (.A1_N(_0629_),
    .A2_N(_1152_),
    .B1(_1150_),
    .B2(\core_1.execute.sreg_priv_control.o_d[4] ),
    .X(_1161_));
 sky130_fd_sc_hd__and2_1 _4112_ (.A(_1156_),
    .B(_1161_),
    .X(_1162_));
 sky130_fd_sc_hd__clkbuf_1 _4113_ (.A(_1162_),
    .X(_0070_));
 sky130_fd_sc_hd__nand2_1 _4114_ (.A(\core_1.execute.sreg_priv_control.o_d[5] ),
    .B(_1150_),
    .Y(_1163_));
 sky130_fd_sc_hd__or3_1 _4115_ (.A(_1146_),
    .B(_0623_),
    .C(_1152_),
    .X(_1164_));
 sky130_fd_sc_hd__buf_4 _4116_ (.A(_0659_),
    .X(_1165_));
 sky130_fd_sc_hd__a21oi_1 _4117_ (.A1(_1163_),
    .A2(_1164_),
    .B1(_1165_),
    .Y(_0071_));
 sky130_fd_sc_hd__a2bb2o_1 _4118_ (.A1_N(_0617_),
    .A2_N(_1152_),
    .B1(_1150_),
    .B2(\core_1.execute.sreg_priv_control.o_d[6] ),
    .X(_1166_));
 sky130_fd_sc_hd__and2_1 _4119_ (.A(_1156_),
    .B(_1166_),
    .X(_1167_));
 sky130_fd_sc_hd__clkbuf_1 _4120_ (.A(_1167_),
    .X(_0072_));
 sky130_fd_sc_hd__a2bb2o_1 _4121_ (.A1_N(_0611_),
    .A2_N(_1152_),
    .B1(_1150_),
    .B2(\core_1.execute.sreg_priv_control.o_d[7] ),
    .X(_1168_));
 sky130_fd_sc_hd__and2_1 _4122_ (.A(_1156_),
    .B(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__clkbuf_1 _4123_ (.A(_1169_),
    .X(_0073_));
 sky130_fd_sc_hd__a2bb2o_1 _4124_ (.A1_N(_0603_),
    .A2_N(_1152_),
    .B1(_1150_),
    .B2(\core_1.execute.sreg_priv_control.o_d[8] ),
    .X(_1170_));
 sky130_fd_sc_hd__and2_1 _4125_ (.A(_1156_),
    .B(_1170_),
    .X(_1171_));
 sky130_fd_sc_hd__clkbuf_1 _4126_ (.A(_1171_),
    .X(_0074_));
 sky130_fd_sc_hd__a2bb2o_1 _4127_ (.A1_N(_0596_),
    .A2_N(_1148_),
    .B1(_1149_),
    .B2(\core_1.execute.sreg_priv_control.o_d[9] ),
    .X(_1172_));
 sky130_fd_sc_hd__and2_1 _4128_ (.A(_1156_),
    .B(_1172_),
    .X(_1173_));
 sky130_fd_sc_hd__clkbuf_1 _4129_ (.A(_1173_),
    .X(_0075_));
 sky130_fd_sc_hd__a2bb2o_1 _4130_ (.A1_N(_0588_),
    .A2_N(_1148_),
    .B1(_1149_),
    .B2(\core_1.execute.sreg_priv_control.o_d[10] ),
    .X(_1174_));
 sky130_fd_sc_hd__and2_1 _4131_ (.A(_1156_),
    .B(_1174_),
    .X(_1175_));
 sky130_fd_sc_hd__clkbuf_1 _4132_ (.A(_1175_),
    .X(_0076_));
 sky130_fd_sc_hd__a2bb2o_1 _4133_ (.A1_N(_0582_),
    .A2_N(_1148_),
    .B1(_1149_),
    .B2(\core_1.execute.sreg_priv_control.o_d[11] ),
    .X(_1176_));
 sky130_fd_sc_hd__and2_1 _4134_ (.A(_1156_),
    .B(_1176_),
    .X(_1177_));
 sky130_fd_sc_hd__clkbuf_1 _4135_ (.A(_1177_),
    .X(_0077_));
 sky130_fd_sc_hd__buf_4 _4136_ (.A(_1154_),
    .X(_1178_));
 sky130_fd_sc_hd__a2bb2o_1 _4137_ (.A1_N(_0575_),
    .A2_N(_1148_),
    .B1(_1149_),
    .B2(\core_1.execute.sreg_priv_control.o_d[12] ),
    .X(_1179_));
 sky130_fd_sc_hd__and2_1 _4138_ (.A(_1178_),
    .B(_1179_),
    .X(_1180_));
 sky130_fd_sc_hd__clkbuf_1 _4139_ (.A(_1180_),
    .X(_0078_));
 sky130_fd_sc_hd__nand2_1 _4140_ (.A(\core_1.execute.sreg_priv_control.o_d[13] ),
    .B(_1150_),
    .Y(_1181_));
 sky130_fd_sc_hd__or3_1 _4141_ (.A(_1146_),
    .B(_0568_),
    .C(_1152_),
    .X(_1182_));
 sky130_fd_sc_hd__a21oi_1 _4142_ (.A1(_1181_),
    .A2(_1182_),
    .B1(_1165_),
    .Y(_0079_));
 sky130_fd_sc_hd__a2bb2o_1 _4143_ (.A1_N(_0553_),
    .A2_N(_1148_),
    .B1(_1149_),
    .B2(\core_1.execute.sreg_priv_control.o_d[14] ),
    .X(_1183_));
 sky130_fd_sc_hd__and2_1 _4144_ (.A(_1178_),
    .B(_1183_),
    .X(_1184_));
 sky130_fd_sc_hd__clkbuf_1 _4145_ (.A(_1184_),
    .X(_0080_));
 sky130_fd_sc_hd__nand2_1 _4146_ (.A(\core_1.execute.sreg_priv_control.o_d[15] ),
    .B(_1150_),
    .Y(_1185_));
 sky130_fd_sc_hd__or3_1 _4147_ (.A(_1146_),
    .B(_0545_),
    .C(_1152_),
    .X(_1186_));
 sky130_fd_sc_hd__a21oi_1 _4148_ (.A1(_1185_),
    .A2(_1186_),
    .B1(_1165_),
    .Y(_0081_));
 sky130_fd_sc_hd__clkbuf_4 _4149_ (.A(\core_1.execute.alu_mul_div.cbit[3] ),
    .X(_1187_));
 sky130_fd_sc_hd__clkbuf_4 _4150_ (.A(_1187_),
    .X(_1188_));
 sky130_fd_sc_hd__inv_2 _4151_ (.A(\core_1.execute.alu_mul_div.cbit[2] ),
    .Y(_1189_));
 sky130_fd_sc_hd__clkbuf_4 _4152_ (.A(_1189_),
    .X(_1190_));
 sky130_fd_sc_hd__buf_4 _4153_ (.A(_1190_),
    .X(_1191_));
 sky130_fd_sc_hd__buf_4 _4154_ (.A(\core_1.execute.alu_mul_div.cbit[0] ),
    .X(_1192_));
 sky130_fd_sc_hd__buf_4 _4155_ (.A(\core_1.execute.alu_mul_div.cbit[1] ),
    .X(_1193_));
 sky130_fd_sc_hd__nand2_4 _4156_ (.A(_1192_),
    .B(_1193_),
    .Y(_1194_));
 sky130_fd_sc_hd__nor2_2 _4157_ (.A(_1191_),
    .B(_1194_),
    .Y(_1195_));
 sky130_fd_sc_hd__nand2_2 _4158_ (.A(_1188_),
    .B(_1195_),
    .Y(_1196_));
 sky130_fd_sc_hd__clkbuf_4 _4159_ (.A(_1196_),
    .X(_1197_));
 sky130_fd_sc_hd__or4b_2 _4160_ (.A(\core_1.decode.i_flush ),
    .B(_0659_),
    .C(_0688_),
    .D_N(_0731_),
    .X(_1198_));
 sky130_fd_sc_hd__o21ba_1 _4161_ (.A1(_0730_),
    .A2(_1197_),
    .B1_N(_1198_),
    .X(_0082_));
 sky130_fd_sc_hd__inv_2 _4162_ (.A(_1001_),
    .Y(_1199_));
 sky130_fd_sc_hd__or4b_1 _4163_ (.A(_0659_),
    .B(_0737_),
    .C(_1199_),
    .D_N(net70),
    .X(_1200_));
 sky130_fd_sc_hd__clkbuf_4 _4164_ (.A(_1200_),
    .X(_1201_));
 sky130_fd_sc_hd__buf_4 _4165_ (.A(_1201_),
    .X(_1202_));
 sky130_fd_sc_hd__mux2_1 _4166_ (.A0(net38),
    .A1(\core_1.fetch.out_buffer_data_instr[0] ),
    .S(_1202_),
    .X(_1203_));
 sky130_fd_sc_hd__clkbuf_1 _4167_ (.A(_1203_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _4168_ (.A0(net49),
    .A1(\core_1.fetch.out_buffer_data_instr[1] ),
    .S(_1202_),
    .X(_1204_));
 sky130_fd_sc_hd__clkbuf_1 _4169_ (.A(_1204_),
    .X(_0084_));
 sky130_fd_sc_hd__mux2_1 _4170_ (.A0(net60),
    .A1(\core_1.fetch.out_buffer_data_instr[2] ),
    .S(_1202_),
    .X(_1205_));
 sky130_fd_sc_hd__clkbuf_1 _4171_ (.A(_1205_),
    .X(_0085_));
 sky130_fd_sc_hd__mux2_1 _4172_ (.A0(net63),
    .A1(\core_1.fetch.out_buffer_data_instr[3] ),
    .S(_1202_),
    .X(_1206_));
 sky130_fd_sc_hd__clkbuf_1 _4173_ (.A(_1206_),
    .X(_0086_));
 sky130_fd_sc_hd__mux2_1 _4174_ (.A0(net64),
    .A1(\core_1.fetch.out_buffer_data_instr[4] ),
    .S(_1202_),
    .X(_1207_));
 sky130_fd_sc_hd__clkbuf_1 _4175_ (.A(_1207_),
    .X(_0087_));
 sky130_fd_sc_hd__mux2_1 _4176_ (.A0(net65),
    .A1(\core_1.fetch.out_buffer_data_instr[5] ),
    .S(_1202_),
    .X(_1208_));
 sky130_fd_sc_hd__clkbuf_1 _4177_ (.A(_1208_),
    .X(_0088_));
 sky130_fd_sc_hd__mux2_1 _4178_ (.A0(net66),
    .A1(\core_1.fetch.out_buffer_data_instr[6] ),
    .S(_1202_),
    .X(_1209_));
 sky130_fd_sc_hd__clkbuf_1 _4179_ (.A(_1209_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _4180_ (.A0(net67),
    .A1(\core_1.fetch.out_buffer_data_instr[7] ),
    .S(_1202_),
    .X(_1210_));
 sky130_fd_sc_hd__clkbuf_1 _4181_ (.A(_1210_),
    .X(_0090_));
 sky130_fd_sc_hd__mux2_1 _4182_ (.A0(net68),
    .A1(\core_1.fetch.out_buffer_data_instr[8] ),
    .S(_1202_),
    .X(_1211_));
 sky130_fd_sc_hd__clkbuf_1 _4183_ (.A(_1211_),
    .X(_0091_));
 sky130_fd_sc_hd__mux2_1 _4184_ (.A0(net69),
    .A1(\core_1.fetch.out_buffer_data_instr[9] ),
    .S(_1202_),
    .X(_1212_));
 sky130_fd_sc_hd__clkbuf_1 _4185_ (.A(_1212_),
    .X(_0092_));
 sky130_fd_sc_hd__buf_4 _4186_ (.A(_1201_),
    .X(_1213_));
 sky130_fd_sc_hd__mux2_1 _4187_ (.A0(net39),
    .A1(\core_1.fetch.out_buffer_data_instr[10] ),
    .S(_1213_),
    .X(_1214_));
 sky130_fd_sc_hd__clkbuf_1 _4188_ (.A(_1214_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _4189_ (.A0(net40),
    .A1(\core_1.fetch.out_buffer_data_instr[11] ),
    .S(_1213_),
    .X(_1215_));
 sky130_fd_sc_hd__clkbuf_1 _4190_ (.A(_1215_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _4191_ (.A0(net41),
    .A1(\core_1.fetch.out_buffer_data_instr[12] ),
    .S(_1213_),
    .X(_1216_));
 sky130_fd_sc_hd__clkbuf_1 _4192_ (.A(_1216_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _4193_ (.A0(net42),
    .A1(\core_1.fetch.out_buffer_data_instr[13] ),
    .S(_1213_),
    .X(_1217_));
 sky130_fd_sc_hd__clkbuf_1 _4194_ (.A(_1217_),
    .X(_0096_));
 sky130_fd_sc_hd__mux2_1 _4195_ (.A0(net43),
    .A1(\core_1.fetch.out_buffer_data_instr[14] ),
    .S(_1213_),
    .X(_1218_));
 sky130_fd_sc_hd__clkbuf_1 _4196_ (.A(_1218_),
    .X(_0097_));
 sky130_fd_sc_hd__mux2_1 _4197_ (.A0(net44),
    .A1(\core_1.fetch.out_buffer_data_instr[15] ),
    .S(_1213_),
    .X(_1219_));
 sky130_fd_sc_hd__clkbuf_1 _4198_ (.A(_1219_),
    .X(_0098_));
 sky130_fd_sc_hd__mux2_1 _4199_ (.A0(net45),
    .A1(\core_1.fetch.out_buffer_data_instr[16] ),
    .S(_1213_),
    .X(_1220_));
 sky130_fd_sc_hd__clkbuf_1 _4200_ (.A(_1220_),
    .X(_0099_));
 sky130_fd_sc_hd__mux2_1 _4201_ (.A0(net46),
    .A1(\core_1.fetch.out_buffer_data_instr[17] ),
    .S(_1213_),
    .X(_1221_));
 sky130_fd_sc_hd__clkbuf_1 _4202_ (.A(_1221_),
    .X(_0100_));
 sky130_fd_sc_hd__mux2_1 _4203_ (.A0(net47),
    .A1(\core_1.fetch.out_buffer_data_instr[18] ),
    .S(_1213_),
    .X(_1222_));
 sky130_fd_sc_hd__clkbuf_1 _4204_ (.A(_1222_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _4205_ (.A0(net48),
    .A1(\core_1.fetch.out_buffer_data_instr[19] ),
    .S(_1213_),
    .X(_1223_));
 sky130_fd_sc_hd__clkbuf_1 _4206_ (.A(_1223_),
    .X(_0102_));
 sky130_fd_sc_hd__buf_4 _4207_ (.A(_1201_),
    .X(_1224_));
 sky130_fd_sc_hd__mux2_1 _4208_ (.A0(net50),
    .A1(\core_1.fetch.out_buffer_data_instr[20] ),
    .S(_1224_),
    .X(_1225_));
 sky130_fd_sc_hd__clkbuf_1 _4209_ (.A(_1225_),
    .X(_0103_));
 sky130_fd_sc_hd__mux2_1 _4210_ (.A0(net51),
    .A1(\core_1.fetch.out_buffer_data_instr[21] ),
    .S(_1224_),
    .X(_1226_));
 sky130_fd_sc_hd__clkbuf_1 _4211_ (.A(_1226_),
    .X(_0104_));
 sky130_fd_sc_hd__mux2_1 _4212_ (.A0(net52),
    .A1(\core_1.fetch.out_buffer_data_instr[22] ),
    .S(_1224_),
    .X(_1227_));
 sky130_fd_sc_hd__clkbuf_1 _4213_ (.A(_1227_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _4214_ (.A0(net53),
    .A1(\core_1.fetch.out_buffer_data_instr[23] ),
    .S(_1224_),
    .X(_1228_));
 sky130_fd_sc_hd__clkbuf_1 _4215_ (.A(_1228_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _4216_ (.A0(net54),
    .A1(\core_1.fetch.out_buffer_data_instr[24] ),
    .S(_1224_),
    .X(_1229_));
 sky130_fd_sc_hd__clkbuf_1 _4217_ (.A(_1229_),
    .X(_0107_));
 sky130_fd_sc_hd__mux2_1 _4218_ (.A0(net55),
    .A1(\core_1.fetch.out_buffer_data_instr[25] ),
    .S(_1224_),
    .X(_1230_));
 sky130_fd_sc_hd__clkbuf_1 _4219_ (.A(_1230_),
    .X(_0108_));
 sky130_fd_sc_hd__mux2_1 _4220_ (.A0(net56),
    .A1(\core_1.fetch.out_buffer_data_instr[26] ),
    .S(_1224_),
    .X(_1231_));
 sky130_fd_sc_hd__clkbuf_1 _4221_ (.A(_1231_),
    .X(_0109_));
 sky130_fd_sc_hd__mux2_1 _4222_ (.A0(net57),
    .A1(\core_1.fetch.out_buffer_data_instr[27] ),
    .S(_1224_),
    .X(_1232_));
 sky130_fd_sc_hd__clkbuf_1 _4223_ (.A(_1232_),
    .X(_0110_));
 sky130_fd_sc_hd__mux2_1 _4224_ (.A0(net58),
    .A1(\core_1.fetch.out_buffer_data_instr[28] ),
    .S(_1224_),
    .X(_1233_));
 sky130_fd_sc_hd__clkbuf_1 _4225_ (.A(_1233_),
    .X(_0111_));
 sky130_fd_sc_hd__mux2_1 _4226_ (.A0(net59),
    .A1(\core_1.fetch.out_buffer_data_instr[29] ),
    .S(_1224_),
    .X(_1234_));
 sky130_fd_sc_hd__clkbuf_1 _4227_ (.A(_1234_),
    .X(_0112_));
 sky130_fd_sc_hd__mux2_1 _4228_ (.A0(net61),
    .A1(\core_1.fetch.out_buffer_data_instr[30] ),
    .S(_1201_),
    .X(_1235_));
 sky130_fd_sc_hd__clkbuf_1 _4229_ (.A(_1235_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_1 _4230_ (.A0(net62),
    .A1(\core_1.fetch.out_buffer_data_instr[31] ),
    .S(_1201_),
    .X(_1236_));
 sky130_fd_sc_hd__clkbuf_1 _4231_ (.A(_1236_),
    .X(_0114_));
 sky130_fd_sc_hd__a21o_1 _4232_ (.A1(net70),
    .A2(_1001_),
    .B1(_0664_),
    .X(_1237_));
 sky130_fd_sc_hd__o211a_1 _4233_ (.A1(\core_1.decode.input_valid ),
    .A2(_0736_),
    .B1(_0809_),
    .C1(_1237_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_1 _4234_ (.A0(\core_1.fetch.current_req_branch_pred ),
    .A1(\core_1.fetch.out_buffer_data_pred ),
    .S(_1201_),
    .X(_1238_));
 sky130_fd_sc_hd__clkbuf_1 _4235_ (.A(_1238_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_1 _4236_ (.A0(\core_1.fetch.prev_request_pc[0] ),
    .A1(net161),
    .S(net177),
    .X(_1239_));
 sky130_fd_sc_hd__clkbuf_1 _4237_ (.A(_1239_),
    .X(_0117_));
 sky130_fd_sc_hd__mux2_1 _4238_ (.A0(\core_1.fetch.prev_request_pc[1] ),
    .A1(net168),
    .S(net177),
    .X(_1240_));
 sky130_fd_sc_hd__clkbuf_1 _4239_ (.A(_1240_),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _4240_ (.A0(\core_1.fetch.prev_request_pc[2] ),
    .A1(net169),
    .S(net177),
    .X(_1241_));
 sky130_fd_sc_hd__clkbuf_1 _4241_ (.A(_1241_),
    .X(_0119_));
 sky130_fd_sc_hd__mux2_1 _4242_ (.A0(\core_1.fetch.prev_request_pc[3] ),
    .A1(net170),
    .S(net177),
    .X(_1242_));
 sky130_fd_sc_hd__clkbuf_1 _4243_ (.A(_1242_),
    .X(_0120_));
 sky130_fd_sc_hd__mux2_1 _4244_ (.A0(\core_1.fetch.prev_request_pc[4] ),
    .A1(net171),
    .S(net177),
    .X(_1243_));
 sky130_fd_sc_hd__clkbuf_1 _4245_ (.A(_1243_),
    .X(_0121_));
 sky130_fd_sc_hd__mux2_1 _4246_ (.A0(\core_1.fetch.prev_request_pc[5] ),
    .A1(net172),
    .S(net177),
    .X(_1244_));
 sky130_fd_sc_hd__clkbuf_1 _4247_ (.A(_1244_),
    .X(_0122_));
 sky130_fd_sc_hd__mux2_1 _4248_ (.A0(\core_1.fetch.prev_request_pc[6] ),
    .A1(net173),
    .S(net177),
    .X(_1245_));
 sky130_fd_sc_hd__clkbuf_1 _4249_ (.A(_1245_),
    .X(_0123_));
 sky130_fd_sc_hd__mux2_1 _4250_ (.A0(\core_1.fetch.prev_request_pc[7] ),
    .A1(net174),
    .S(net177),
    .X(_1246_));
 sky130_fd_sc_hd__clkbuf_1 _4251_ (.A(_1246_),
    .X(_0124_));
 sky130_fd_sc_hd__mux2_1 _4252_ (.A0(\core_1.fetch.prev_request_pc[8] ),
    .A1(net175),
    .S(_0779_),
    .X(_1247_));
 sky130_fd_sc_hd__clkbuf_1 _4253_ (.A(_1247_),
    .X(_0125_));
 sky130_fd_sc_hd__mux2_1 _4254_ (.A0(\core_1.fetch.prev_request_pc[9] ),
    .A1(net176),
    .S(_0779_),
    .X(_1248_));
 sky130_fd_sc_hd__clkbuf_1 _4255_ (.A(_1248_),
    .X(_0126_));
 sky130_fd_sc_hd__mux2_1 _4256_ (.A0(\core_1.fetch.prev_request_pc[10] ),
    .A1(net162),
    .S(_0779_),
    .X(_1249_));
 sky130_fd_sc_hd__clkbuf_1 _4257_ (.A(_1249_),
    .X(_0127_));
 sky130_fd_sc_hd__mux2_1 _4258_ (.A0(\core_1.fetch.prev_request_pc[11] ),
    .A1(net163),
    .S(_0779_),
    .X(_1250_));
 sky130_fd_sc_hd__clkbuf_1 _4259_ (.A(_1250_),
    .X(_0128_));
 sky130_fd_sc_hd__mux2_1 _4260_ (.A0(\core_1.fetch.prev_request_pc[12] ),
    .A1(net164),
    .S(_0779_),
    .X(_1251_));
 sky130_fd_sc_hd__clkbuf_1 _4261_ (.A(_1251_),
    .X(_0129_));
 sky130_fd_sc_hd__mux2_1 _4262_ (.A0(\core_1.fetch.prev_request_pc[13] ),
    .A1(net165),
    .S(_0779_),
    .X(_1252_));
 sky130_fd_sc_hd__clkbuf_1 _4263_ (.A(_1252_),
    .X(_0130_));
 sky130_fd_sc_hd__mux2_1 _4264_ (.A0(\core_1.fetch.prev_request_pc[14] ),
    .A1(net166),
    .S(_0779_),
    .X(_1253_));
 sky130_fd_sc_hd__clkbuf_1 _4265_ (.A(_1253_),
    .X(_0131_));
 sky130_fd_sc_hd__mux2_1 _4266_ (.A0(\core_1.fetch.prev_request_pc[15] ),
    .A1(net167),
    .S(_0779_),
    .X(_1254_));
 sky130_fd_sc_hd__clkbuf_1 _4267_ (.A(_1254_),
    .X(_0132_));
 sky130_fd_sc_hd__buf_4 _4268_ (.A(_1002_),
    .X(_1255_));
 sky130_fd_sc_hd__mux2_1 _4269_ (.A0(_0739_),
    .A1(\core_1.decode.i_instr_l[0] ),
    .S(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__clkbuf_1 _4270_ (.A(_1256_),
    .X(_0133_));
 sky130_fd_sc_hd__mux2_1 _4271_ (.A0(_0740_),
    .A1(\core_1.decode.i_instr_l[1] ),
    .S(_1255_),
    .X(_1257_));
 sky130_fd_sc_hd__clkbuf_1 _4272_ (.A(_1257_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _4273_ (.A0(_0742_),
    .A1(\core_1.decode.i_instr_l[2] ),
    .S(_1255_),
    .X(_1258_));
 sky130_fd_sc_hd__clkbuf_1 _4274_ (.A(_1258_),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _4275_ (.A0(_0743_),
    .A1(\core_1.decode.i_instr_l[3] ),
    .S(_1255_),
    .X(_1259_));
 sky130_fd_sc_hd__clkbuf_1 _4276_ (.A(_1259_),
    .X(_0136_));
 sky130_fd_sc_hd__mux2_1 _4277_ (.A0(_0772_),
    .A1(\core_1.decode.i_instr_l[4] ),
    .S(_1255_),
    .X(_1260_));
 sky130_fd_sc_hd__clkbuf_1 _4278_ (.A(_1260_),
    .X(_0137_));
 sky130_fd_sc_hd__mux2_1 _4279_ (.A0(_0774_),
    .A1(\core_1.decode.i_instr_l[5] ),
    .S(_1255_),
    .X(_1261_));
 sky130_fd_sc_hd__clkbuf_1 _4280_ (.A(_1261_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_1 _4281_ (.A0(_0773_),
    .A1(\core_1.decode.i_instr_l[6] ),
    .S(_1255_),
    .X(_1262_));
 sky130_fd_sc_hd__clkbuf_1 _4282_ (.A(_1262_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_1 _4283_ (.A0(_0913_),
    .A1(\core_1.decode.i_instr_l[7] ),
    .S(_1255_),
    .X(_1263_));
 sky130_fd_sc_hd__clkbuf_1 _4284_ (.A(_1263_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_1 _4285_ (.A0(_0915_),
    .A1(\core_1.decode.i_instr_l[8] ),
    .S(_1255_),
    .X(_1264_));
 sky130_fd_sc_hd__clkbuf_1 _4286_ (.A(_1264_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_1 _4287_ (.A0(_0912_),
    .A1(\core_1.decode.i_instr_l[9] ),
    .S(_1255_),
    .X(_1265_));
 sky130_fd_sc_hd__clkbuf_1 _4288_ (.A(_1265_),
    .X(_0142_));
 sky130_fd_sc_hd__buf_4 _4289_ (.A(_1002_),
    .X(_1266_));
 sky130_fd_sc_hd__mux2_1 _4290_ (.A0(_0914_),
    .A1(\core_1.decode.i_instr_l[10] ),
    .S(_1266_),
    .X(_1267_));
 sky130_fd_sc_hd__clkbuf_1 _4291_ (.A(_1267_),
    .X(_0143_));
 sky130_fd_sc_hd__mux2_1 _4292_ (.A0(net40),
    .A1(\core_1.fetch.out_buffer_data_instr[11] ),
    .S(_0664_),
    .X(_1268_));
 sky130_fd_sc_hd__mux2_1 _4293_ (.A0(_1268_),
    .A1(\core_1.decode.i_instr_l[11] ),
    .S(_1266_),
    .X(_1269_));
 sky130_fd_sc_hd__clkbuf_1 _4294_ (.A(_1269_),
    .X(_0144_));
 sky130_fd_sc_hd__mux2_1 _4295_ (.A0(net41),
    .A1(\core_1.fetch.out_buffer_data_instr[12] ),
    .S(_0664_),
    .X(_1270_));
 sky130_fd_sc_hd__mux2_1 _4296_ (.A0(_1270_),
    .A1(\core_1.decode.i_instr_l[12] ),
    .S(_1266_),
    .X(_1271_));
 sky130_fd_sc_hd__clkbuf_1 _4297_ (.A(_1271_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_1 _4298_ (.A0(net42),
    .A1(\core_1.fetch.out_buffer_data_instr[13] ),
    .S(_0664_),
    .X(_1272_));
 sky130_fd_sc_hd__mux2_1 _4299_ (.A0(_1272_),
    .A1(\core_1.decode.i_instr_l[13] ),
    .S(_1266_),
    .X(_1273_));
 sky130_fd_sc_hd__clkbuf_1 _4300_ (.A(_1273_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_1 _4301_ (.A0(net43),
    .A1(\core_1.fetch.out_buffer_data_instr[14] ),
    .S(_0664_),
    .X(_1274_));
 sky130_fd_sc_hd__mux2_1 _4302_ (.A0(_1274_),
    .A1(\core_1.decode.i_instr_l[14] ),
    .S(_1266_),
    .X(_1275_));
 sky130_fd_sc_hd__clkbuf_1 _4303_ (.A(_1275_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_1 _4304_ (.A0(net44),
    .A1(\core_1.fetch.out_buffer_data_instr[15] ),
    .S(_0664_),
    .X(_1276_));
 sky130_fd_sc_hd__mux2_1 _4305_ (.A0(_1276_),
    .A1(\core_1.decode.i_instr_l[15] ),
    .S(_1266_),
    .X(_1277_));
 sky130_fd_sc_hd__clkbuf_1 _4306_ (.A(_1277_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_1 _4307_ (.A0(_0757_),
    .A1(\core_1.decode.i_imm_pass[0] ),
    .S(_1266_),
    .X(_1278_));
 sky130_fd_sc_hd__clkbuf_1 _4308_ (.A(_1278_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_1 _4309_ (.A0(_0747_),
    .A1(\core_1.decode.i_imm_pass[1] ),
    .S(_1266_),
    .X(_1279_));
 sky130_fd_sc_hd__clkbuf_1 _4310_ (.A(_1279_),
    .X(_0150_));
 sky130_fd_sc_hd__mux2_1 _4311_ (.A0(_0753_),
    .A1(\core_1.decode.i_imm_pass[2] ),
    .S(_1266_),
    .X(_1280_));
 sky130_fd_sc_hd__clkbuf_1 _4312_ (.A(_1280_),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _4313_ (.A0(_0746_),
    .A1(\core_1.decode.i_imm_pass[3] ),
    .S(_1266_),
    .X(_1281_));
 sky130_fd_sc_hd__clkbuf_1 _4314_ (.A(_1281_),
    .X(_0152_));
 sky130_fd_sc_hd__buf_4 _4315_ (.A(_1002_),
    .X(_1282_));
 sky130_fd_sc_hd__mux2_1 _4316_ (.A0(_0752_),
    .A1(\core_1.decode.i_imm_pass[4] ),
    .S(_1282_),
    .X(_1283_));
 sky130_fd_sc_hd__clkbuf_1 _4317_ (.A(_1283_),
    .X(_0153_));
 sky130_fd_sc_hd__mux2_1 _4318_ (.A0(_0758_),
    .A1(\core_1.decode.i_imm_pass[5] ),
    .S(_1282_),
    .X(_1284_));
 sky130_fd_sc_hd__clkbuf_1 _4319_ (.A(_1284_),
    .X(_0154_));
 sky130_fd_sc_hd__mux2_1 _4320_ (.A0(_0766_),
    .A1(\core_1.decode.i_imm_pass[6] ),
    .S(_1282_),
    .X(_1285_));
 sky130_fd_sc_hd__clkbuf_1 _4321_ (.A(_1285_),
    .X(_0155_));
 sky130_fd_sc_hd__mux2_1 _4322_ (.A0(_0754_),
    .A1(\core_1.decode.i_imm_pass[7] ),
    .S(_1282_),
    .X(_1286_));
 sky130_fd_sc_hd__clkbuf_1 _4323_ (.A(_1286_),
    .X(_0156_));
 sky130_fd_sc_hd__mux2_1 _4324_ (.A0(_0749_),
    .A1(\core_1.decode.i_imm_pass[8] ),
    .S(_1282_),
    .X(_1287_));
 sky130_fd_sc_hd__clkbuf_1 _4325_ (.A(_1287_),
    .X(_0157_));
 sky130_fd_sc_hd__mux2_1 _4326_ (.A0(_0763_),
    .A1(\core_1.decode.i_imm_pass[9] ),
    .S(_1282_),
    .X(_1288_));
 sky130_fd_sc_hd__clkbuf_1 _4327_ (.A(_1288_),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _4328_ (.A0(_0748_),
    .A1(\core_1.decode.i_imm_pass[10] ),
    .S(_1282_),
    .X(_1289_));
 sky130_fd_sc_hd__clkbuf_1 _4329_ (.A(_1289_),
    .X(_0159_));
 sky130_fd_sc_hd__mux2_1 _4330_ (.A0(_0765_),
    .A1(\core_1.decode.i_imm_pass[11] ),
    .S(_1282_),
    .X(_1290_));
 sky130_fd_sc_hd__clkbuf_1 _4331_ (.A(_1290_),
    .X(_0160_));
 sky130_fd_sc_hd__mux2_1 _4332_ (.A0(_0756_),
    .A1(\core_1.decode.i_imm_pass[12] ),
    .S(_1282_),
    .X(_1291_));
 sky130_fd_sc_hd__clkbuf_1 _4333_ (.A(_1291_),
    .X(_0161_));
 sky130_fd_sc_hd__mux2_1 _4334_ (.A0(_0767_),
    .A1(\core_1.decode.i_imm_pass[13] ),
    .S(_1282_),
    .X(_1292_));
 sky130_fd_sc_hd__clkbuf_1 _4335_ (.A(_1292_),
    .X(_0162_));
 sky130_fd_sc_hd__mux2_1 _4336_ (.A0(_0751_),
    .A1(\core_1.decode.i_imm_pass[14] ),
    .S(_1002_),
    .X(_1293_));
 sky130_fd_sc_hd__clkbuf_1 _4337_ (.A(_1293_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_1 _4338_ (.A0(_0760_),
    .A1(\core_1.decode.i_imm_pass[15] ),
    .S(_1002_),
    .X(_1294_));
 sky130_fd_sc_hd__clkbuf_1 _4339_ (.A(_1294_),
    .X(_0164_));
 sky130_fd_sc_hd__nor2_1 _4340_ (.A(_1055_),
    .B(net70),
    .Y(_1295_));
 sky130_fd_sc_hd__a21o_1 _4341_ (.A1(\core_1.fetch.dbg_out ),
    .A2(_1295_),
    .B1(net177),
    .X(_0165_));
 sky130_fd_sc_hd__o211a_1 _4342_ (.A1(\core_1.fetch.flush_event_invalidate ),
    .A2(\core_1.fetch.dbg_out ),
    .B1(_1199_),
    .C1(_1295_),
    .X(_0166_));
 sky130_fd_sc_hd__and3_1 _4343_ (.A(_1178_),
    .B(_0778_),
    .C(_0926_),
    .X(_1296_));
 sky130_fd_sc_hd__clkbuf_1 _4344_ (.A(_1296_),
    .X(_0167_));
 sky130_fd_sc_hd__clkbuf_1 _4345_ (.A(_1055_),
    .X(_1297_));
 sky130_fd_sc_hd__clkbuf_1 _4346_ (.A(_1297_),
    .X(_0168_));
 sky130_fd_sc_hd__inv_2 _4347_ (.A(net37),
    .Y(_1298_));
 sky130_fd_sc_hd__buf_4 _4348_ (.A(\core_1.ew_mem_access ),
    .X(_1299_));
 sky130_fd_sc_hd__buf_4 _4349_ (.A(_1299_),
    .X(_1300_));
 sky130_fd_sc_hd__mux2_1 _4350_ (.A0(_1298_),
    .A1(_1300_),
    .S(\core_1.ew_submit ),
    .X(_1301_));
 sky130_fd_sc_hd__and3_1 _4351_ (.A(_1178_),
    .B(_0726_),
    .C(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__clkbuf_1 _4352_ (.A(_1302_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_1 _4353_ (.A0(\core_1.fetch.current_req_branch_pred ),
    .A1(\core_1.fetch.out_buffer_data_pred ),
    .S(_0664_),
    .X(_1303_));
 sky130_fd_sc_hd__mux2_1 _4354_ (.A0(\core_1.decode.i_jmp_pred_pass ),
    .A1(_1303_),
    .S(\core_1.fetch.submitable ),
    .X(_1304_));
 sky130_fd_sc_hd__clkbuf_1 _4355_ (.A(_1304_),
    .X(_0170_));
 sky130_fd_sc_hd__nor2_2 _4356_ (.A(_1020_),
    .B(_1040_),
    .Y(_1305_));
 sky130_fd_sc_hd__or2_4 _4357_ (.A(_0733_),
    .B(_1305_),
    .X(_1306_));
 sky130_fd_sc_hd__clkbuf_4 _4358_ (.A(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__nand2_2 _4359_ (.A(_1141_),
    .B(\core_1.dec_sreg_store ),
    .Y(_1308_));
 sky130_fd_sc_hd__clkbuf_4 _4360_ (.A(_1308_),
    .X(_1309_));
 sky130_fd_sc_hd__nand2_1 _4361_ (.A(\core_1.execute.sreg_irq_pc.o_d[1] ),
    .B(\core_1.dec_sreg_irt ),
    .Y(_1310_));
 sky130_fd_sc_hd__nor2_2 _4362_ (.A(_1146_),
    .B(_1057_),
    .Y(_1311_));
 sky130_fd_sc_hd__clkinv_2 _4363_ (.A(\core_1.execute.alu_mul_div.i_mod ),
    .Y(_1312_));
 sky130_fd_sc_hd__clkbuf_4 _4364_ (.A(_1312_),
    .X(_1313_));
 sky130_fd_sc_hd__buf_2 _4365_ (.A(_0727_),
    .X(_1314_));
 sky130_fd_sc_hd__a21bo_1 _4366_ (.A1(\core_1.execute.alu_mul_div.div_res[1] ),
    .A2(_1313_),
    .B1_N(_1314_),
    .X(_1315_));
 sky130_fd_sc_hd__inv_2 _4367_ (.A(\core_1.execute.alu_mul_div.i_mul ),
    .Y(_1316_));
 sky130_fd_sc_hd__nand2_4 _4368_ (.A(net185),
    .B(\core_1.dec_r_bus_imm ),
    .Y(_1317_));
 sky130_fd_sc_hd__a311o_4 _4369_ (.A1(_0644_),
    .A2(_0645_),
    .A3(_0648_),
    .B1(_0649_),
    .C1(\core_1.dec_r_bus_imm ),
    .X(_1318_));
 sky130_fd_sc_hd__nand2_4 _4370_ (.A(_1317_),
    .B(_1318_),
    .Y(_1319_));
 sky130_fd_sc_hd__inv_2 _4371_ (.A(\core_1.dec_r_bus_imm ),
    .Y(_1320_));
 sky130_fd_sc_hd__buf_8 _4372_ (.A(_1320_),
    .X(_1321_));
 sky130_fd_sc_hd__nor2_2 _4373_ (.A(_1009_),
    .B(_1321_),
    .Y(_1322_));
 sky130_fd_sc_hd__o221a_2 _4374_ (.A1(net88),
    .A2(_0517_),
    .B1(_0652_),
    .B2(_0657_),
    .C1(_1320_),
    .X(_1323_));
 sky130_fd_sc_hd__nor2_2 _4375_ (.A(_1322_),
    .B(_1323_),
    .Y(_1324_));
 sky130_fd_sc_hd__nor2_1 _4376_ (.A(_1319_),
    .B(_1324_),
    .Y(_1325_));
 sky130_fd_sc_hd__nand2_4 _4377_ (.A(net211),
    .B(_1079_),
    .Y(_1326_));
 sky130_fd_sc_hd__o221ai_4 _4378_ (.A1(net88),
    .A2(_0517_),
    .B1(_0652_),
    .B2(_0657_),
    .C1(_1321_),
    .Y(_1327_));
 sky130_fd_sc_hd__nand2_4 _4379_ (.A(_1326_),
    .B(_1327_),
    .Y(_1328_));
 sky130_fd_sc_hd__nand2_1 _4380_ (.A(\core_1.decode.oc_alu_mode[12] ),
    .B(_1328_),
    .Y(_1329_));
 sky130_fd_sc_hd__a22o_4 _4381_ (.A1(\core_1.decode.oc_alu_mode[12] ),
    .A2(_1325_),
    .B1(_1329_),
    .B2(_1319_),
    .X(_1330_));
 sky130_fd_sc_hd__clkbuf_4 _4382_ (.A(\core_1.decode.oc_alu_mode[12] ),
    .X(_1331_));
 sky130_fd_sc_hd__and3_1 _4383_ (.A(\core_1.execute.rf.reg_outputs[7][0] ),
    .B(\core_1.dec_l_reg_sel[2] ),
    .C(\core_1.dec_l_reg_sel[1] ),
    .X(_1332_));
 sky130_fd_sc_hd__and3b_1 _4384_ (.A_N(_0698_),
    .B(\core_1.dec_l_reg_sel[2] ),
    .C(\core_1.execute.rf.reg_outputs[5][0] ),
    .X(_1333_));
 sky130_fd_sc_hd__and3b_1 _4385_ (.A_N(_0716_),
    .B(_0698_),
    .C(\core_1.execute.rf.reg_outputs[3][0] ),
    .X(_1334_));
 sky130_fd_sc_hd__o31a_1 _4386_ (.A1(_1332_),
    .A2(_1333_),
    .A3(_1334_),
    .B1(_0694_),
    .X(_1335_));
 sky130_fd_sc_hd__nor3b_4 _4387_ (.A(_0716_),
    .B(\core_1.dec_l_reg_sel[0] ),
    .C_N(\core_1.dec_l_reg_sel[1] ),
    .Y(_1336_));
 sky130_fd_sc_hd__nor3b_4 _4388_ (.A(\core_1.dec_l_reg_sel[0] ),
    .B(_0698_),
    .C_N(_0716_),
    .Y(_1337_));
 sky130_fd_sc_hd__a22o_1 _4389_ (.A1(\core_1.execute.rf.reg_outputs[2][0] ),
    .A2(_1336_),
    .B1(_1337_),
    .B2(\core_1.execute.rf.reg_outputs[4][0] ),
    .X(_1338_));
 sky130_fd_sc_hd__nor2_1 _4390_ (.A(\core_1.dec_l_reg_sel[2] ),
    .B(\core_1.dec_l_reg_sel[1] ),
    .Y(_1339_));
 sky130_fd_sc_hd__and3b_4 _4391_ (.A_N(\core_1.dec_l_reg_sel[0] ),
    .B(\core_1.dec_l_reg_sel[1] ),
    .C(\core_1.dec_l_reg_sel[2] ),
    .X(_1340_));
 sky130_fd_sc_hd__nor3_4 _4392_ (.A(\core_1.dec_l_reg_sel[2] ),
    .B(\core_1.dec_l_reg_sel[0] ),
    .C(\core_1.dec_l_reg_sel[1] ),
    .Y(_1341_));
 sky130_fd_sc_hd__a221o_1 _4393_ (.A1(\core_1.execute.rf.reg_outputs[1][0] ),
    .A2(_1339_),
    .B1(_1340_),
    .B2(\core_1.execute.rf.reg_outputs[6][0] ),
    .C1(_1341_),
    .X(_1342_));
 sky130_fd_sc_hd__or3_4 _4394_ (.A(_1335_),
    .B(_1338_),
    .C(_1342_),
    .X(_1343_));
 sky130_fd_sc_hd__nand2_2 _4395_ (.A(_0692_),
    .B(_0700_),
    .Y(_1344_));
 sky130_fd_sc_hd__or2_4 _4396_ (.A(net88),
    .B(_1344_),
    .X(_1345_));
 sky130_fd_sc_hd__and2_4 _4397_ (.A(_1343_),
    .B(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__mux2_8 _4398_ (.A0(net191),
    .A1(net207),
    .S(_1321_),
    .X(_1347_));
 sky130_fd_sc_hd__mux2_2 _4399_ (.A0(net190),
    .A1(net206),
    .S(_1321_),
    .X(_1348_));
 sky130_fd_sc_hd__or2_1 _4400_ (.A(_1347_),
    .B(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__buf_8 _4401_ (.A(_1321_),
    .X(_1350_));
 sky130_fd_sc_hd__mux2_8 _4402_ (.A0(net183),
    .A1(net199),
    .S(_1350_),
    .X(_1351_));
 sky130_fd_sc_hd__mux2_4 _4403_ (.A0(net179),
    .A1(net195),
    .S(_1321_),
    .X(_1352_));
 sky130_fd_sc_hd__mux2_2 _4404_ (.A0(net180),
    .A1(net196),
    .S(_1321_),
    .X(_1353_));
 sky130_fd_sc_hd__mux2_8 _4405_ (.A0(net193),
    .A1(net209),
    .S(_1321_),
    .X(_1354_));
 sky130_fd_sc_hd__mux2_8 _4406_ (.A0(net192),
    .A1(net208),
    .S(_1321_),
    .X(_1355_));
 sky130_fd_sc_hd__or4_1 _4407_ (.A(_1352_),
    .B(_1353_),
    .C(_1354_),
    .D(_1355_),
    .X(_1356_));
 sky130_fd_sc_hd__inv_2 _4408_ (.A(net184),
    .Y(_1357_));
 sky130_fd_sc_hd__mux2_8 _4409_ (.A0(_1357_),
    .A1(_0545_),
    .S(_1350_),
    .X(_1358_));
 sky130_fd_sc_hd__or4b_4 _4410_ (.A(_1349_),
    .B(_1351_),
    .C(_1356_),
    .D_N(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__inv_2 _4411_ (.A(\core_1.decode.oc_alu_mode[12] ),
    .Y(_1360_));
 sky130_fd_sc_hd__nand2_1 _4412_ (.A(net189),
    .B(_1079_),
    .Y(_1361_));
 sky130_fd_sc_hd__o21a_2 _4413_ (.A1(_1079_),
    .A2(_0623_),
    .B1(_1361_),
    .X(_1362_));
 sky130_fd_sc_hd__buf_4 _4414_ (.A(_1362_),
    .X(_1363_));
 sky130_fd_sc_hd__and4_2 _4415_ (.A(_1317_),
    .B(_1318_),
    .C(_1326_),
    .D(_1327_),
    .X(_1364_));
 sky130_fd_sc_hd__nand2_1 _4416_ (.A(net187),
    .B(_1079_),
    .Y(_1365_));
 sky130_fd_sc_hd__o21a_4 _4417_ (.A1(_1079_),
    .A2(_0635_),
    .B1(_1365_),
    .X(_1366_));
 sky130_fd_sc_hd__mux2_2 _4418_ (.A0(_1010_),
    .A1(_0643_),
    .S(_1350_),
    .X(_1367_));
 sky130_fd_sc_hd__nor2_2 _4419_ (.A(net188),
    .B(_1321_),
    .Y(_1368_));
 sky130_fd_sc_hd__a211o_1 _4420_ (.A1(_1350_),
    .A2(_0629_),
    .B1(_1368_),
    .C1(_1360_),
    .X(_1369_));
 sky130_fd_sc_hd__a31o_1 _4421_ (.A1(_1364_),
    .A2(_1366_),
    .A3(_1367_),
    .B1(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__mux2_8 _4422_ (.A0(net182),
    .A1(net198),
    .S(_1350_),
    .X(_1371_));
 sky130_fd_sc_hd__nand2_1 _4423_ (.A(net181),
    .B(_1079_),
    .Y(_1372_));
 sky130_fd_sc_hd__o21ai_4 _4424_ (.A1(_1079_),
    .A2(_0575_),
    .B1(_1372_),
    .Y(_1373_));
 sky130_fd_sc_hd__nor2_1 _4425_ (.A(_1371_),
    .B(_1373_),
    .Y(_1374_));
 sky130_fd_sc_hd__o211a_1 _4426_ (.A1(_1360_),
    .A2(_1363_),
    .B1(_1370_),
    .C1(_1374_),
    .X(_1375_));
 sky130_fd_sc_hd__buf_6 _4427_ (.A(_1344_),
    .X(_1376_));
 sky130_fd_sc_hd__buf_6 _4428_ (.A(_1376_),
    .X(_1377_));
 sky130_fd_sc_hd__nor2_2 _4429_ (.A(_0717_),
    .B(_0699_),
    .Y(_1378_));
 sky130_fd_sc_hd__nor2_4 _4430_ (.A(_0693_),
    .B(_0699_),
    .Y(_1379_));
 sky130_fd_sc_hd__clkbuf_4 _4431_ (.A(_1336_),
    .X(_1380_));
 sky130_fd_sc_hd__a22o_1 _4432_ (.A1(\core_1.execute.rf.reg_outputs[5][15] ),
    .A2(_1379_),
    .B1(_1380_),
    .B2(\core_1.execute.rf.reg_outputs[2][15] ),
    .X(_1381_));
 sky130_fd_sc_hd__nor2_4 _4433_ (.A(_0693_),
    .B(_0696_),
    .Y(_1382_));
 sky130_fd_sc_hd__nor2_4 _4434_ (.A(_0717_),
    .B(_0696_),
    .Y(_1383_));
 sky130_fd_sc_hd__buf_4 _4435_ (.A(_1340_),
    .X(_1384_));
 sky130_fd_sc_hd__or2b_1 _4436_ (.A(\core_1.execute.rf.reg_outputs[4][15] ),
    .B_N(_0717_),
    .X(_1385_));
 sky130_fd_sc_hd__a22o_1 _4437_ (.A1(\core_1.execute.rf.reg_outputs[6][15] ),
    .A2(_1384_),
    .B1(_1385_),
    .B2(_0700_),
    .X(_1386_));
 sky130_fd_sc_hd__a221o_1 _4438_ (.A1(\core_1.execute.rf.reg_outputs[7][15] ),
    .A2(_1382_),
    .B1(_1383_),
    .B2(\core_1.execute.rf.reg_outputs[3][15] ),
    .C1(_1386_),
    .X(_1387_));
 sky130_fd_sc_hd__a211o_2 _4439_ (.A1(\core_1.execute.rf.reg_outputs[1][15] ),
    .A2(_1378_),
    .B1(_1381_),
    .C1(_1387_),
    .X(_1388_));
 sky130_fd_sc_hd__o21ai_4 _4440_ (.A1(net94),
    .A2(_1377_),
    .B1(_1388_),
    .Y(_1389_));
 sky130_fd_sc_hd__nand2_1 _4441_ (.A(\core_1.decode.oc_alu_mode[12] ),
    .B(_1389_),
    .Y(_1390_));
 sky130_fd_sc_hd__and3b_1 _4442_ (.A_N(_1359_),
    .B(_1375_),
    .C(_1390_),
    .X(_1391_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _4443_ (.A(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__buf_2 _4444_ (.A(_1392_),
    .X(_1393_));
 sky130_fd_sc_hd__o21ai_4 _4445_ (.A1(_1331_),
    .A2(_1346_),
    .B1(_1393_),
    .Y(_1394_));
 sky130_fd_sc_hd__a22o_1 _4446_ (.A1(\core_1.execute.rf.reg_outputs[2][1] ),
    .A2(_1336_),
    .B1(_1337_),
    .B2(\core_1.execute.rf.reg_outputs[4][1] ),
    .X(_1395_));
 sky130_fd_sc_hd__and3_1 _4447_ (.A(\core_1.execute.rf.reg_outputs[7][1] ),
    .B(_0716_),
    .C(_0698_),
    .X(_1396_));
 sky130_fd_sc_hd__and3b_1 _4448_ (.A_N(_0698_),
    .B(_0716_),
    .C(\core_1.execute.rf.reg_outputs[5][1] ),
    .X(_1397_));
 sky130_fd_sc_hd__and3b_1 _4449_ (.A_N(_0716_),
    .B(_0698_),
    .C(\core_1.execute.rf.reg_outputs[3][1] ),
    .X(_1398_));
 sky130_fd_sc_hd__o31a_1 _4450_ (.A1(_1396_),
    .A2(_1397_),
    .A3(_1398_),
    .B1(_0694_),
    .X(_1399_));
 sky130_fd_sc_hd__clkbuf_4 _4451_ (.A(_1339_),
    .X(_1400_));
 sky130_fd_sc_hd__a221o_1 _4452_ (.A1(\core_1.execute.rf.reg_outputs[1][1] ),
    .A2(_1400_),
    .B1(_1340_),
    .B2(\core_1.execute.rf.reg_outputs[6][1] ),
    .C1(_1341_),
    .X(_1401_));
 sky130_fd_sc_hd__or3_2 _4453_ (.A(_1395_),
    .B(_1399_),
    .C(_1401_),
    .X(_1402_));
 sky130_fd_sc_hd__o21ai_4 _4454_ (.A1(net95),
    .A2(_1376_),
    .B1(_1402_),
    .Y(_1403_));
 sky130_fd_sc_hd__clkinv_2 _4455_ (.A(_1403_),
    .Y(_1404_));
 sky130_fd_sc_hd__o21ai_1 _4456_ (.A1(_0822_),
    .A2(_1404_),
    .B1(_1393_),
    .Y(_1405_));
 sky130_fd_sc_hd__buf_4 _4457_ (.A(_1324_),
    .X(_1406_));
 sky130_fd_sc_hd__buf_4 _4458_ (.A(_1406_),
    .X(_1407_));
 sky130_fd_sc_hd__mux2_1 _4459_ (.A0(_1394_),
    .A1(_1405_),
    .S(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__or2_2 _4460_ (.A(_1330_),
    .B(_1408_),
    .X(_1409_));
 sky130_fd_sc_hd__a21oi_4 _4461_ (.A1(_1350_),
    .A2(_0629_),
    .B1(_1368_),
    .Y(_1410_));
 sky130_fd_sc_hd__o21ai_4 _4462_ (.A1(_1079_),
    .A2(_0635_),
    .B1(_1365_),
    .Y(_1411_));
 sky130_fd_sc_hd__mux2_2 _4463_ (.A0(net186),
    .A1(net202),
    .S(_1350_),
    .X(_1412_));
 sky130_fd_sc_hd__buf_4 _4464_ (.A(_1412_),
    .X(_1413_));
 sky130_fd_sc_hd__nor2_2 _4465_ (.A(_1411_),
    .B(_1413_),
    .Y(_1414_));
 sky130_fd_sc_hd__and3_1 _4466_ (.A(\core_1.decode.oc_alu_mode[12] ),
    .B(_1364_),
    .C(_1414_),
    .X(_1415_));
 sky130_fd_sc_hd__xnor2_2 _4467_ (.A(_1410_),
    .B(_1415_),
    .Y(_1416_));
 sky130_fd_sc_hd__o211ai_4 _4468_ (.A1(_0822_),
    .A2(\core_1.decode.oc_alu_mode[13] ),
    .B1(_1363_),
    .C1(_1416_),
    .Y(_1417_));
 sky130_fd_sc_hd__buf_4 _4469_ (.A(_1367_),
    .X(_1418_));
 sky130_fd_sc_hd__nand2_2 _4470_ (.A(_1364_),
    .B(_1418_),
    .Y(_1419_));
 sky130_fd_sc_hd__nand2_4 _4471_ (.A(_0822_),
    .B(_1419_),
    .Y(_1420_));
 sky130_fd_sc_hd__xnor2_4 _4472_ (.A(_1411_),
    .B(_1420_),
    .Y(_1421_));
 sky130_fd_sc_hd__nor2_2 _4473_ (.A(_1417_),
    .B(_1421_),
    .Y(_1422_));
 sky130_fd_sc_hd__nor2_4 _4474_ (.A(_1360_),
    .B(_1364_),
    .Y(_1423_));
 sky130_fd_sc_hd__xnor2_4 _4475_ (.A(_1413_),
    .B(_1423_),
    .Y(_1424_));
 sky130_fd_sc_hd__nand2_2 _4476_ (.A(_1422_),
    .B(_1424_),
    .Y(_1425_));
 sky130_fd_sc_hd__and2_1 _4477_ (.A(_1317_),
    .B(_1318_),
    .X(_1426_));
 sky130_fd_sc_hd__buf_2 _4478_ (.A(_1426_),
    .X(_1427_));
 sky130_fd_sc_hd__a22o_1 _4479_ (.A1(_1326_),
    .A2(_1327_),
    .B1(_1343_),
    .B2(_1345_),
    .X(_1428_));
 sky130_fd_sc_hd__nand2_1 _4480_ (.A(\core_1.execute.alu_flag_reg.o_d[1] ),
    .B(\core_1.dec_alu_carry_en ),
    .Y(_1429_));
 sky130_fd_sc_hd__a41o_1 _4481_ (.A1(_1326_),
    .A2(_1327_),
    .A3(_1343_),
    .A4(_1345_),
    .B1(_1429_),
    .X(_1430_));
 sky130_fd_sc_hd__and3_1 _4482_ (.A(_1427_),
    .B(_1428_),
    .C(_1430_),
    .X(_1431_));
 sky130_fd_sc_hd__a21oi_1 _4483_ (.A1(_1428_),
    .A2(_1430_),
    .B1(_1427_),
    .Y(_1432_));
 sky130_fd_sc_hd__o21ai_1 _4484_ (.A1(_1431_),
    .A2(_1432_),
    .B1(_1403_),
    .Y(_1433_));
 sky130_fd_sc_hd__o31a_1 _4485_ (.A1(_1403_),
    .A2(_1431_),
    .A3(_1432_),
    .B1(_0862_),
    .X(_1434_));
 sky130_fd_sc_hd__nor2_1 _4486_ (.A(_1427_),
    .B(_1403_),
    .Y(_1435_));
 sky130_fd_sc_hd__nand2_2 _4487_ (.A(_1427_),
    .B(_1403_),
    .Y(_1436_));
 sky130_fd_sc_hd__and2b_1 _4488_ (.A_N(_1435_),
    .B(_1436_),
    .X(_1437_));
 sky130_fd_sc_hd__inv_2 _4489_ (.A(_1429_),
    .Y(_1438_));
 sky130_fd_sc_hd__a211o_1 _4490_ (.A1(_1343_),
    .A2(_1345_),
    .B1(_1322_),
    .C1(_1323_),
    .X(_1439_));
 sky130_fd_sc_hd__o211a_1 _4491_ (.A1(_1322_),
    .A2(_1323_),
    .B1(_1343_),
    .C1(_1345_),
    .X(_1440_));
 sky130_fd_sc_hd__a21o_1 _4492_ (.A1(_1438_),
    .A2(_1439_),
    .B1(_1440_),
    .X(_1441_));
 sky130_fd_sc_hd__xor2_1 _4493_ (.A(_1437_),
    .B(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__or4_1 _4494_ (.A(\core_1.decode.oc_alu_mode[7] ),
    .B(\core_1.decode.oc_alu_mode[11] ),
    .C(\core_1.decode.oc_alu_mode[3] ),
    .D(\core_1.decode.oc_alu_mode[1] ),
    .X(_1443_));
 sky130_fd_sc_hd__or4_1 _4495_ (.A(\core_1.decode.oc_alu_mode[4] ),
    .B(\core_1.decode.oc_alu_mode[12] ),
    .C(\core_1.decode.oc_alu_mode[2] ),
    .D(\core_1.decode.oc_alu_mode[13] ),
    .X(_1444_));
 sky130_fd_sc_hd__nor4_4 _4496_ (.A(\core_1.decode.oc_alu_mode[9] ),
    .B(\core_1.decode.oc_alu_mode[6] ),
    .C(_1443_),
    .D(_1444_),
    .Y(_1445_));
 sky130_fd_sc_hd__or2_2 _4497_ (.A(\core_1.decode.oc_alu_mode[3] ),
    .B(_1445_),
    .X(_1446_));
 sky130_fd_sc_hd__a22o_1 _4498_ (.A1(\core_1.decode.oc_alu_mode[7] ),
    .A2(_1319_),
    .B1(_1404_),
    .B2(_1446_),
    .X(_1447_));
 sky130_fd_sc_hd__a221o_1 _4499_ (.A1(_0814_),
    .A2(_1436_),
    .B1(_1437_),
    .B2(\core_1.decode.oc_alu_mode[6] ),
    .C1(_1447_),
    .X(_1448_));
 sky130_fd_sc_hd__a221o_1 _4500_ (.A1(_0839_),
    .A2(_1435_),
    .B1(_1442_),
    .B2(\core_1.decode.oc_alu_mode[4] ),
    .C1(_1448_),
    .X(_1449_));
 sky130_fd_sc_hd__a21oi_2 _4501_ (.A1(_1433_),
    .A2(_1434_),
    .B1(_1449_),
    .Y(_1450_));
 sky130_fd_sc_hd__buf_4 _4502_ (.A(_1411_),
    .X(_1451_));
 sky130_fd_sc_hd__a22o_1 _4503_ (.A1(\core_1.execute.rf.reg_outputs[5][10] ),
    .A2(_1379_),
    .B1(_1383_),
    .B2(\core_1.execute.rf.reg_outputs[3][10] ),
    .X(_1452_));
 sky130_fd_sc_hd__o21a_1 _4504_ (.A1(\core_1.execute.rf.reg_outputs[4][10] ),
    .A2(_0693_),
    .B1(_0700_),
    .X(_1453_));
 sky130_fd_sc_hd__a221o_1 _4505_ (.A1(\core_1.execute.rf.reg_outputs[1][10] ),
    .A2(_1378_),
    .B1(_1380_),
    .B2(\core_1.execute.rf.reg_outputs[2][10] ),
    .C1(_1453_),
    .X(_1454_));
 sky130_fd_sc_hd__a221o_1 _4506_ (.A1(\core_1.execute.rf.reg_outputs[7][10] ),
    .A2(_1382_),
    .B1(_1384_),
    .B2(\core_1.execute.rf.reg_outputs[6][10] ),
    .C1(_1454_),
    .X(_1455_));
 sky130_fd_sc_hd__o22a_2 _4507_ (.A1(net89),
    .A2(_1377_),
    .B1(_1452_),
    .B2(_1455_),
    .X(_1456_));
 sky130_fd_sc_hd__buf_4 _4508_ (.A(_1456_),
    .X(_1457_));
 sky130_fd_sc_hd__inv_2 _4509_ (.A(_1457_),
    .Y(_1458_));
 sky130_fd_sc_hd__clkbuf_4 _4510_ (.A(_1400_),
    .X(_1459_));
 sky130_fd_sc_hd__and3_1 _4511_ (.A(\core_1.execute.rf.reg_outputs[1][9] ),
    .B(_0694_),
    .C(_1459_),
    .X(_1460_));
 sky130_fd_sc_hd__a22o_1 _4512_ (.A1(\core_1.execute.rf.reg_outputs[5][9] ),
    .A2(_1379_),
    .B1(_1380_),
    .B2(\core_1.execute.rf.reg_outputs[2][9] ),
    .X(_1461_));
 sky130_fd_sc_hd__or2b_1 _4513_ (.A(\core_1.execute.rf.reg_outputs[4][9] ),
    .B_N(_0717_),
    .X(_1462_));
 sky130_fd_sc_hd__a22o_1 _4514_ (.A1(\core_1.execute.rf.reg_outputs[6][9] ),
    .A2(_1340_),
    .B1(_1462_),
    .B2(_0700_),
    .X(_1463_));
 sky130_fd_sc_hd__a221o_1 _4515_ (.A1(\core_1.execute.rf.reg_outputs[7][9] ),
    .A2(_1382_),
    .B1(_1383_),
    .B2(\core_1.execute.rf.reg_outputs[3][9] ),
    .C1(_1463_),
    .X(_1464_));
 sky130_fd_sc_hd__o32a_4 _4516_ (.A1(_1460_),
    .A2(_1461_),
    .A3(_1464_),
    .B1(_1376_),
    .B2(net103),
    .X(_1465_));
 sky130_fd_sc_hd__inv_2 _4517_ (.A(_1465_),
    .Y(_1466_));
 sky130_fd_sc_hd__mux2_1 _4518_ (.A0(_1458_),
    .A1(_1466_),
    .S(_1324_),
    .X(_1467_));
 sky130_fd_sc_hd__o21ai_4 _4519_ (.A1(_1079_),
    .A2(_0623_),
    .B1(_1361_),
    .Y(_1468_));
 sky130_fd_sc_hd__or3b_1 _4520_ (.A(_1468_),
    .B(_1359_),
    .C_N(_1374_),
    .X(_1469_));
 sky130_fd_sc_hd__or2_2 _4521_ (.A(_1319_),
    .B(_1469_),
    .X(_1470_));
 sky130_fd_sc_hd__a22o_1 _4522_ (.A1(\core_1.execute.rf.reg_outputs[7][12] ),
    .A2(_1382_),
    .B1(_1384_),
    .B2(\core_1.execute.rf.reg_outputs[6][12] ),
    .X(_1471_));
 sky130_fd_sc_hd__and2b_4 _4523_ (.A_N(\core_1.dec_l_reg_sel[2] ),
    .B(\core_1.dec_l_reg_sel[1] ),
    .X(_1472_));
 sky130_fd_sc_hd__and3_1 _4524_ (.A(\core_1.execute.rf.reg_outputs[3][12] ),
    .B(_0701_),
    .C(_1472_),
    .X(_1473_));
 sky130_fd_sc_hd__or2_1 _4525_ (.A(\core_1.execute.rf.reg_outputs[4][12] ),
    .B(_0693_),
    .X(_1474_));
 sky130_fd_sc_hd__a22o_1 _4526_ (.A1(\core_1.execute.rf.reg_outputs[1][12] ),
    .A2(_1378_),
    .B1(_1474_),
    .B2(_0700_),
    .X(_1475_));
 sky130_fd_sc_hd__a221o_1 _4527_ (.A1(\core_1.execute.rf.reg_outputs[5][12] ),
    .A2(_1379_),
    .B1(_1380_),
    .B2(\core_1.execute.rf.reg_outputs[2][12] ),
    .C1(_1475_),
    .X(_1476_));
 sky130_fd_sc_hd__o32a_4 _4528_ (.A1(_1471_),
    .A2(_1473_),
    .A3(_1476_),
    .B1(_1377_),
    .B2(net91),
    .X(_1477_));
 sky130_fd_sc_hd__inv_2 _4529_ (.A(_1477_),
    .Y(_1478_));
 sky130_fd_sc_hd__and3_1 _4530_ (.A(\core_1.execute.rf.reg_outputs[1][11] ),
    .B(_0694_),
    .C(_1400_),
    .X(_1479_));
 sky130_fd_sc_hd__a221o_2 _4531_ (.A1(\core_1.execute.rf.reg_outputs[5][11] ),
    .A2(_1379_),
    .B1(_1380_),
    .B2(\core_1.execute.rf.reg_outputs[2][11] ),
    .C1(_1479_),
    .X(_1480_));
 sky130_fd_sc_hd__or2b_1 _4532_ (.A(\core_1.execute.rf.reg_outputs[4][11] ),
    .B_N(_0717_),
    .X(_1481_));
 sky130_fd_sc_hd__a22o_1 _4533_ (.A1(\core_1.execute.rf.reg_outputs[6][11] ),
    .A2(_1384_),
    .B1(_1481_),
    .B2(_0700_),
    .X(_1482_));
 sky130_fd_sc_hd__a221o_2 _4534_ (.A1(\core_1.execute.rf.reg_outputs[7][11] ),
    .A2(_1382_),
    .B1(_1383_),
    .B2(\core_1.execute.rf.reg_outputs[3][11] ),
    .C1(_1482_),
    .X(_1483_));
 sky130_fd_sc_hd__o22ai_4 _4535_ (.A1(net90),
    .A2(_1376_),
    .B1(_1480_),
    .B2(_1483_),
    .Y(_1484_));
 sky130_fd_sc_hd__mux2_1 _4536_ (.A0(_1478_),
    .A1(_1484_),
    .S(_1406_),
    .X(_1485_));
 sky130_fd_sc_hd__or2_2 _4537_ (.A(_1427_),
    .B(_1469_),
    .X(_1486_));
 sky130_fd_sc_hd__o22a_1 _4538_ (.A1(_1467_),
    .A2(_1470_),
    .B1(_1485_),
    .B2(_1486_),
    .X(_1487_));
 sky130_fd_sc_hd__clkbuf_4 _4539_ (.A(_1328_),
    .X(_1488_));
 sky130_fd_sc_hd__a22o_1 _4540_ (.A1(\core_1.execute.rf.reg_outputs[3][13] ),
    .A2(_1383_),
    .B1(_1380_),
    .B2(\core_1.execute.rf.reg_outputs[2][13] ),
    .X(_1489_));
 sky130_fd_sc_hd__o21a_1 _4541_ (.A1(\core_1.execute.rf.reg_outputs[4][13] ),
    .A2(_0693_),
    .B1(_0700_),
    .X(_1490_));
 sky130_fd_sc_hd__a221o_1 _4542_ (.A1(\core_1.execute.rf.reg_outputs[5][13] ),
    .A2(_1379_),
    .B1(_1378_),
    .B2(\core_1.execute.rf.reg_outputs[1][13] ),
    .C1(_1490_),
    .X(_1491_));
 sky130_fd_sc_hd__a221o_1 _4543_ (.A1(\core_1.execute.rf.reg_outputs[7][13] ),
    .A2(_1382_),
    .B1(_1384_),
    .B2(\core_1.execute.rf.reg_outputs[6][13] ),
    .C1(_1491_),
    .X(_1492_));
 sky130_fd_sc_hd__o22a_4 _4544_ (.A1(net92),
    .A2(_1377_),
    .B1(_1489_),
    .B2(_1492_),
    .X(_1493_));
 sky130_fd_sc_hd__inv_2 _4545_ (.A(_1493_),
    .Y(_1494_));
 sky130_fd_sc_hd__a22o_1 _4546_ (.A1(\core_1.execute.rf.reg_outputs[5][14] ),
    .A2(_1379_),
    .B1(_1380_),
    .B2(\core_1.execute.rf.reg_outputs[2][14] ),
    .X(_1495_));
 sky130_fd_sc_hd__or2_1 _4547_ (.A(\core_1.execute.rf.reg_outputs[4][14] ),
    .B(_0693_),
    .X(_1496_));
 sky130_fd_sc_hd__a22o_1 _4548_ (.A1(\core_1.execute.rf.reg_outputs[6][14] ),
    .A2(_1384_),
    .B1(_1496_),
    .B2(_0700_),
    .X(_1497_));
 sky130_fd_sc_hd__a221o_1 _4549_ (.A1(\core_1.execute.rf.reg_outputs[7][14] ),
    .A2(_1382_),
    .B1(_1383_),
    .B2(\core_1.execute.rf.reg_outputs[3][14] ),
    .C1(_1497_),
    .X(_1498_));
 sky130_fd_sc_hd__a211o_2 _4550_ (.A1(\core_1.execute.rf.reg_outputs[1][14] ),
    .A2(_1378_),
    .B1(_1495_),
    .C1(_1498_),
    .X(_1499_));
 sky130_fd_sc_hd__o21ai_4 _4551_ (.A1(net93),
    .A2(_1377_),
    .B1(_1499_),
    .Y(_1500_));
 sky130_fd_sc_hd__mux2_1 _4552_ (.A0(_1494_),
    .A1(_1500_),
    .S(_1328_),
    .X(_1501_));
 sky130_fd_sc_hd__o32a_1 _4553_ (.A1(_1488_),
    .A2(_1389_),
    .A3(_1486_),
    .B1(_1501_),
    .B2(_1470_),
    .X(_1502_));
 sky130_fd_sc_hd__mux2_1 _4554_ (.A0(_1487_),
    .A1(_1502_),
    .S(_1413_),
    .X(_1503_));
 sky130_fd_sc_hd__buf_6 _4555_ (.A(_1366_),
    .X(_1504_));
 sky130_fd_sc_hd__buf_4 _4556_ (.A(_1413_),
    .X(_1505_));
 sky130_fd_sc_hd__buf_2 _4557_ (.A(_1469_),
    .X(_1506_));
 sky130_fd_sc_hd__or2_1 _4558_ (.A(_1505_),
    .B(_1506_),
    .X(_1507_));
 sky130_fd_sc_hd__a22o_1 _4559_ (.A1(\core_1.execute.rf.reg_outputs[1][6] ),
    .A2(_1400_),
    .B1(_1340_),
    .B2(\core_1.execute.rf.reg_outputs[6][6] ),
    .X(_1508_));
 sky130_fd_sc_hd__a22o_1 _4560_ (.A1(\core_1.execute.rf.reg_outputs[2][6] ),
    .A2(_1336_),
    .B1(_1337_),
    .B2(\core_1.execute.rf.reg_outputs[4][6] ),
    .X(_1509_));
 sky130_fd_sc_hd__o21a_2 _4561_ (.A1(_1508_),
    .A2(_1509_),
    .B1(_1344_),
    .X(_1510_));
 sky130_fd_sc_hd__and2b_2 _4562_ (.A_N(\core_1.dec_l_reg_sel[1] ),
    .B(\core_1.dec_l_reg_sel[2] ),
    .X(_1511_));
 sky130_fd_sc_hd__and3_1 _4563_ (.A(\core_1.execute.rf.reg_outputs[7][6] ),
    .B(_0716_),
    .C(_0698_),
    .X(_1512_));
 sky130_fd_sc_hd__a221o_1 _4564_ (.A1(\core_1.execute.rf.reg_outputs[5][6] ),
    .A2(_1511_),
    .B1(_1472_),
    .B2(\core_1.execute.rf.reg_outputs[3][6] ),
    .C1(_1512_),
    .X(_1513_));
 sky130_fd_sc_hd__and2_1 _4565_ (.A(_0694_),
    .B(_1513_),
    .X(_1514_));
 sky130_fd_sc_hd__a211oi_4 _4566_ (.A1(net100),
    .A2(_1341_),
    .B1(_1510_),
    .C1(_1514_),
    .Y(_1515_));
 sky130_fd_sc_hd__and3_1 _4567_ (.A(\core_1.execute.rf.reg_outputs[7][5] ),
    .B(\core_1.dec_l_reg_sel[2] ),
    .C(\core_1.dec_l_reg_sel[1] ),
    .X(_1516_));
 sky130_fd_sc_hd__a221o_1 _4568_ (.A1(\core_1.execute.rf.reg_outputs[5][5] ),
    .A2(_1511_),
    .B1(_1472_),
    .B2(\core_1.execute.rf.reg_outputs[3][5] ),
    .C1(_1516_),
    .X(_1517_));
 sky130_fd_sc_hd__and2_1 _4569_ (.A(_0694_),
    .B(_1517_),
    .X(_1518_));
 sky130_fd_sc_hd__a221o_1 _4570_ (.A1(\core_1.execute.rf.reg_outputs[1][5] ),
    .A2(_1400_),
    .B1(_1337_),
    .B2(\core_1.execute.rf.reg_outputs[4][5] ),
    .C1(_1341_),
    .X(_1519_));
 sky130_fd_sc_hd__a22o_1 _4571_ (.A1(\core_1.execute.rf.reg_outputs[6][5] ),
    .A2(_1340_),
    .B1(_1336_),
    .B2(\core_1.execute.rf.reg_outputs[2][5] ),
    .X(_1520_));
 sky130_fd_sc_hd__o32a_1 _4572_ (.A1(_1518_),
    .A2(_1519_),
    .A3(_1520_),
    .B1(_1376_),
    .B2(net99),
    .X(_1521_));
 sky130_fd_sc_hd__buf_6 _4573_ (.A(_1521_),
    .X(_1522_));
 sky130_fd_sc_hd__inv_2 _4574_ (.A(_1522_),
    .Y(_1523_));
 sky130_fd_sc_hd__mux2_1 _4575_ (.A0(_1515_),
    .A1(_1523_),
    .S(_1406_),
    .X(_1524_));
 sky130_fd_sc_hd__a22o_1 _4576_ (.A1(\core_1.execute.rf.reg_outputs[1][7] ),
    .A2(_1400_),
    .B1(_1384_),
    .B2(\core_1.execute.rf.reg_outputs[6][7] ),
    .X(_1525_));
 sky130_fd_sc_hd__a221o_1 _4577_ (.A1(\core_1.execute.rf.reg_outputs[2][7] ),
    .A2(_1380_),
    .B1(_1337_),
    .B2(\core_1.execute.rf.reg_outputs[4][7] ),
    .C1(_1525_),
    .X(_1526_));
 sky130_fd_sc_hd__and3_1 _4578_ (.A(\core_1.execute.rf.reg_outputs[7][7] ),
    .B(_0716_),
    .C(_0695_),
    .X(_1527_));
 sky130_fd_sc_hd__a221o_1 _4579_ (.A1(\core_1.execute.rf.reg_outputs[5][7] ),
    .A2(_1511_),
    .B1(_1472_),
    .B2(\core_1.execute.rf.reg_outputs[3][7] ),
    .C1(_1527_),
    .X(_1528_));
 sky130_fd_sc_hd__a22o_1 _4580_ (.A1(net101),
    .A2(_1341_),
    .B1(_1528_),
    .B2(_0701_),
    .X(_1529_));
 sky130_fd_sc_hd__a21o_2 _4581_ (.A1(_1376_),
    .A2(_1526_),
    .B1(_1529_),
    .X(_1530_));
 sky130_fd_sc_hd__buf_4 _4582_ (.A(_1530_),
    .X(_1531_));
 sky130_fd_sc_hd__and3_1 _4583_ (.A(\core_1.execute.rf.reg_outputs[1][8] ),
    .B(_0694_),
    .C(_1400_),
    .X(_1532_));
 sky130_fd_sc_hd__a221o_4 _4584_ (.A1(\core_1.execute.rf.reg_outputs[5][8] ),
    .A2(_1379_),
    .B1(_1380_),
    .B2(\core_1.execute.rf.reg_outputs[2][8] ),
    .C1(_1532_),
    .X(_1533_));
 sky130_fd_sc_hd__or2b_1 _4585_ (.A(\core_1.execute.rf.reg_outputs[4][8] ),
    .B_N(_0717_),
    .X(_1534_));
 sky130_fd_sc_hd__a22o_1 _4586_ (.A1(\core_1.execute.rf.reg_outputs[6][8] ),
    .A2(_1340_),
    .B1(_1534_),
    .B2(_0700_),
    .X(_1535_));
 sky130_fd_sc_hd__a221o_4 _4587_ (.A1(\core_1.execute.rf.reg_outputs[7][8] ),
    .A2(_1382_),
    .B1(_1383_),
    .B2(\core_1.execute.rf.reg_outputs[3][8] ),
    .C1(_1535_),
    .X(_1536_));
 sky130_fd_sc_hd__o22ai_4 _4588_ (.A1(net102),
    .A2(_1377_),
    .B1(_1533_),
    .B2(_1536_),
    .Y(_1537_));
 sky130_fd_sc_hd__nand2_1 _4589_ (.A(_1328_),
    .B(_1537_),
    .Y(_1538_));
 sky130_fd_sc_hd__o21ai_2 _4590_ (.A1(_1328_),
    .A2(_1531_),
    .B1(_1538_),
    .Y(_1539_));
 sky130_fd_sc_hd__o22a_1 _4591_ (.A1(_1470_),
    .A2(_1524_),
    .B1(_1539_),
    .B2(_1486_),
    .X(_1540_));
 sky130_fd_sc_hd__a22o_1 _4592_ (.A1(\core_1.execute.rf.reg_outputs[1][4] ),
    .A2(_1400_),
    .B1(_1384_),
    .B2(\core_1.execute.rf.reg_outputs[6][4] ),
    .X(_1541_));
 sky130_fd_sc_hd__a22o_1 _4593_ (.A1(\core_1.execute.rf.reg_outputs[2][4] ),
    .A2(_1336_),
    .B1(_1337_),
    .B2(\core_1.execute.rf.reg_outputs[4][4] ),
    .X(_1542_));
 sky130_fd_sc_hd__o21a_2 _4594_ (.A1(_1541_),
    .A2(_1542_),
    .B1(_1376_),
    .X(_1543_));
 sky130_fd_sc_hd__and3_1 _4595_ (.A(\core_1.execute.rf.reg_outputs[7][4] ),
    .B(_0716_),
    .C(_0698_),
    .X(_1544_));
 sky130_fd_sc_hd__a221o_1 _4596_ (.A1(\core_1.execute.rf.reg_outputs[5][4] ),
    .A2(_1511_),
    .B1(_1472_),
    .B2(\core_1.execute.rf.reg_outputs[3][4] ),
    .C1(_1544_),
    .X(_1545_));
 sky130_fd_sc_hd__and2_1 _4597_ (.A(_0694_),
    .B(_1545_),
    .X(_1546_));
 sky130_fd_sc_hd__a211oi_4 _4598_ (.A1(net98),
    .A2(_1341_),
    .B1(_1543_),
    .C1(_1546_),
    .Y(_1547_));
 sky130_fd_sc_hd__and3_1 _4599_ (.A(\core_1.execute.rf.reg_outputs[7][3] ),
    .B(_0717_),
    .C(_0695_),
    .X(_1548_));
 sky130_fd_sc_hd__a221o_2 _4600_ (.A1(\core_1.execute.rf.reg_outputs[5][3] ),
    .A2(_1511_),
    .B1(_1472_),
    .B2(\core_1.execute.rf.reg_outputs[3][3] ),
    .C1(_1548_),
    .X(_1549_));
 sky130_fd_sc_hd__a221o_1 _4601_ (.A1(\core_1.execute.rf.reg_outputs[1][3] ),
    .A2(_1400_),
    .B1(_1380_),
    .B2(\core_1.execute.rf.reg_outputs[2][3] ),
    .C1(_1341_),
    .X(_1550_));
 sky130_fd_sc_hd__a22o_1 _4602_ (.A1(\core_1.execute.rf.reg_outputs[6][3] ),
    .A2(_1384_),
    .B1(_1337_),
    .B2(\core_1.execute.rf.reg_outputs[4][3] ),
    .X(_1551_));
 sky130_fd_sc_hd__a211o_1 _4603_ (.A1(_0701_),
    .A2(_1549_),
    .B1(_1550_),
    .C1(_1551_),
    .X(_1552_));
 sky130_fd_sc_hd__o21ai_4 _4604_ (.A1(net97),
    .A2(_1376_),
    .B1(_1552_),
    .Y(_1553_));
 sky130_fd_sc_hd__mux2_1 _4605_ (.A0(_1547_),
    .A1(_1553_),
    .S(_1406_),
    .X(_1554_));
 sky130_fd_sc_hd__buf_4 _4606_ (.A(_1427_),
    .X(_1555_));
 sky130_fd_sc_hd__and3_1 _4607_ (.A(\core_1.execute.rf.reg_outputs[7][2] ),
    .B(_0717_),
    .C(_0695_),
    .X(_1556_));
 sky130_fd_sc_hd__a21o_1 _4608_ (.A1(\core_1.execute.rf.reg_outputs[5][2] ),
    .A2(_1511_),
    .B1(_1556_),
    .X(_1557_));
 sky130_fd_sc_hd__and2_1 _4609_ (.A(\core_1.execute.rf.reg_outputs[3][2] ),
    .B(_1472_),
    .X(_1558_));
 sky130_fd_sc_hd__o21a_1 _4610_ (.A1(_1557_),
    .A2(_1558_),
    .B1(_0701_),
    .X(_1559_));
 sky130_fd_sc_hd__a221o_1 _4611_ (.A1(\core_1.execute.rf.reg_outputs[1][2] ),
    .A2(_1400_),
    .B1(_1336_),
    .B2(\core_1.execute.rf.reg_outputs[2][2] ),
    .C1(_1341_),
    .X(_1560_));
 sky130_fd_sc_hd__a221o_2 _4612_ (.A1(\core_1.execute.rf.reg_outputs[6][2] ),
    .A2(_1384_),
    .B1(_1337_),
    .B2(\core_1.execute.rf.reg_outputs[4][2] ),
    .C1(_1560_),
    .X(_1561_));
 sky130_fd_sc_hd__o22ai_4 _4613_ (.A1(net96),
    .A2(_1376_),
    .B1(_1559_),
    .B2(_1561_),
    .Y(_1562_));
 sky130_fd_sc_hd__and3_1 _4614_ (.A(_1555_),
    .B(_1488_),
    .C(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__a221o_1 _4615_ (.A1(_1364_),
    .A2(_1403_),
    .B1(_1554_),
    .B2(_1319_),
    .C1(_1563_),
    .X(_1564_));
 sky130_fd_sc_hd__a21o_2 _4616_ (.A1(_1350_),
    .A2(_0629_),
    .B1(_1368_),
    .X(_1565_));
 sky130_fd_sc_hd__o21ai_4 _4617_ (.A1(_0822_),
    .A2(\core_1.decode.oc_alu_mode[1] ),
    .B1(_1565_),
    .Y(_1566_));
 sky130_fd_sc_hd__a21o_1 _4618_ (.A1(_1414_),
    .A2(_1564_),
    .B1(_1566_),
    .X(_1567_));
 sky130_fd_sc_hd__a31o_1 _4619_ (.A1(_1504_),
    .A2(_1507_),
    .A3(_1540_),
    .B1(_1567_),
    .X(_1568_));
 sky130_fd_sc_hd__a21o_1 _4620_ (.A1(_1451_),
    .A2(_1503_),
    .B1(_1568_),
    .X(_1569_));
 sky130_fd_sc_hd__o211ai_4 _4621_ (.A1(_1409_),
    .A2(_1425_),
    .B1(_1450_),
    .C1(_1569_),
    .Y(_1570_));
 sky130_fd_sc_hd__a21o_1 _4622_ (.A1(_0859_),
    .A2(\core_1.execute.alu_mul_div.mul_res[1] ),
    .B1(\core_1.execute.alu_mul_div.i_div ),
    .X(_1571_));
 sky130_fd_sc_hd__a21o_1 _4623_ (.A1(_1316_),
    .A2(_1570_),
    .B1(_1571_),
    .X(_1572_));
 sky130_fd_sc_hd__a22o_4 _4624_ (.A1(\core_1.execute.alu_mul_div.div_cur[1] ),
    .A2(_0835_),
    .B1(_1315_),
    .B2(_1572_),
    .X(_1573_));
 sky130_fd_sc_hd__nand2_1 _4625_ (.A(_1311_),
    .B(_1573_),
    .Y(_1574_));
 sky130_fd_sc_hd__o211a_1 _4626_ (.A1(_0650_),
    .A2(_1309_),
    .B1(_1310_),
    .C1(_1574_),
    .X(_1575_));
 sky130_fd_sc_hd__or2_1 _4627_ (.A(\core_1.dec_pc_inc ),
    .B(_1041_),
    .X(_1576_));
 sky130_fd_sc_hd__and3_1 _4628_ (.A(net72),
    .B(_0734_),
    .C(_1576_),
    .X(_1577_));
 sky130_fd_sc_hd__and2_1 _4629_ (.A(net79),
    .B(_1577_),
    .X(_1578_));
 sky130_fd_sc_hd__nor2_1 _4630_ (.A(net79),
    .B(_1577_),
    .Y(_1579_));
 sky130_fd_sc_hd__inv_2 _4631_ (.A(_1306_),
    .Y(_1580_));
 sky130_fd_sc_hd__or3_1 _4632_ (.A(_1578_),
    .B(_1579_),
    .C(_1580_),
    .X(_1581_));
 sky130_fd_sc_hd__o211a_1 _4633_ (.A1(_1307_),
    .A2(_1575_),
    .B1(_1581_),
    .C1(_0668_),
    .X(_1582_));
 sky130_fd_sc_hd__nor2_1 _4634_ (.A(_1056_),
    .B(_1582_),
    .Y(_0171_));
 sky130_fd_sc_hd__nor2_1 _4635_ (.A(\core_1.execute.alu_mul_div.div_cur[15] ),
    .B(_1358_),
    .Y(_1583_));
 sky130_fd_sc_hd__and2b_1 _4636_ (.A_N(\core_1.execute.alu_mul_div.div_cur[14] ),
    .B(_1351_),
    .X(_1584_));
 sky130_fd_sc_hd__inv_2 _4637_ (.A(_1371_),
    .Y(_1585_));
 sky130_fd_sc_hd__and2_1 _4638_ (.A(\core_1.execute.alu_mul_div.div_cur[13] ),
    .B(_1585_),
    .X(_1586_));
 sky130_fd_sc_hd__clkinv_2 _4639_ (.A(_1373_),
    .Y(_1587_));
 sky130_fd_sc_hd__inv_2 _4640_ (.A(net180),
    .Y(_1588_));
 sky130_fd_sc_hd__mux2_8 _4641_ (.A0(_1588_),
    .A1(_0582_),
    .S(_1350_),
    .X(_1589_));
 sky130_fd_sc_hd__or2_1 _4642_ (.A(\core_1.execute.alu_mul_div.div_cur[11] ),
    .B(_1589_),
    .X(_1590_));
 sky130_fd_sc_hd__inv_2 _4643_ (.A(_1352_),
    .Y(_1591_));
 sky130_fd_sc_hd__and2_1 _4644_ (.A(\core_1.execute.alu_mul_div.div_cur[10] ),
    .B(_1591_),
    .X(_1592_));
 sky130_fd_sc_hd__nor2_1 _4645_ (.A(\core_1.execute.alu_mul_div.div_cur[10] ),
    .B(_1591_),
    .Y(_1593_));
 sky130_fd_sc_hd__nor2_1 _4646_ (.A(_1592_),
    .B(_1593_),
    .Y(_1594_));
 sky130_fd_sc_hd__or2b_1 _4647_ (.A(\core_1.execute.alu_mul_div.div_cur[9] ),
    .B_N(_1354_),
    .X(_1595_));
 sky130_fd_sc_hd__inv_2 _4648_ (.A(_1347_),
    .Y(_1596_));
 sky130_fd_sc_hd__or2_1 _4649_ (.A(\core_1.execute.alu_mul_div.div_cur[7] ),
    .B(_1596_),
    .X(_1597_));
 sky130_fd_sc_hd__and2_1 _4650_ (.A(\core_1.execute.alu_mul_div.div_cur[7] ),
    .B(_1596_),
    .X(_1598_));
 sky130_fd_sc_hd__buf_4 _4651_ (.A(_1348_),
    .X(_1599_));
 sky130_fd_sc_hd__and2b_1 _4652_ (.A_N(_1599_),
    .B(\core_1.execute.alu_mul_div.div_cur[6] ),
    .X(_1600_));
 sky130_fd_sc_hd__and2b_1 _4653_ (.A_N(\core_1.execute.alu_mul_div.div_cur[6] ),
    .B(_1599_),
    .X(_1601_));
 sky130_fd_sc_hd__nor2_1 _4654_ (.A(_1600_),
    .B(_1601_),
    .Y(_1602_));
 sky130_fd_sc_hd__or2_1 _4655_ (.A(\core_1.execute.alu_mul_div.div_cur[5] ),
    .B(_1363_),
    .X(_1603_));
 sky130_fd_sc_hd__and2_1 _4656_ (.A(\core_1.execute.alu_mul_div.div_cur[4] ),
    .B(_1565_),
    .X(_1604_));
 sky130_fd_sc_hd__nor2_1 _4657_ (.A(\core_1.execute.alu_mul_div.div_cur[4] ),
    .B(_1565_),
    .Y(_1605_));
 sky130_fd_sc_hd__nor2_1 _4658_ (.A(_1604_),
    .B(_1605_),
    .Y(_1606_));
 sky130_fd_sc_hd__or2_1 _4659_ (.A(\core_1.execute.alu_mul_div.div_cur[3] ),
    .B(_1366_),
    .X(_1607_));
 sky130_fd_sc_hd__xnor2_1 _4660_ (.A(\core_1.execute.alu_mul_div.div_cur[2] ),
    .B(_1412_),
    .Y(_1608_));
 sky130_fd_sc_hd__a21o_1 _4661_ (.A1(_1317_),
    .A2(_1318_),
    .B1(\core_1.execute.alu_mul_div.div_cur[1] ),
    .X(_1609_));
 sky130_fd_sc_hd__a21o_1 _4662_ (.A1(_1326_),
    .A2(_1327_),
    .B1(\core_1.execute.alu_mul_div.div_cur[0] ),
    .X(_1610_));
 sky130_fd_sc_hd__and3_1 _4663_ (.A(\core_1.execute.alu_mul_div.div_cur[1] ),
    .B(_1317_),
    .C(_1318_),
    .X(_1611_));
 sky130_fd_sc_hd__a21o_1 _4664_ (.A1(_1609_),
    .A2(_1610_),
    .B1(_1611_),
    .X(_1612_));
 sky130_fd_sc_hd__and2_1 _4665_ (.A(\core_1.execute.alu_mul_div.div_cur[3] ),
    .B(_1366_),
    .X(_1613_));
 sky130_fd_sc_hd__and2_1 _4666_ (.A(\core_1.execute.alu_mul_div.div_cur[2] ),
    .B(_1367_),
    .X(_1614_));
 sky130_fd_sc_hd__a211o_1 _4667_ (.A1(_1608_),
    .A2(_1612_),
    .B1(_1613_),
    .C1(_1614_),
    .X(_1615_));
 sky130_fd_sc_hd__and2_1 _4668_ (.A(\core_1.execute.alu_mul_div.div_cur[5] ),
    .B(_1363_),
    .X(_1616_));
 sky130_fd_sc_hd__a311o_1 _4669_ (.A1(_1606_),
    .A2(_1607_),
    .A3(_1615_),
    .B1(_1604_),
    .C1(_1616_),
    .X(_1617_));
 sky130_fd_sc_hd__a31o_1 _4670_ (.A1(_1602_),
    .A2(_1603_),
    .A3(_1617_),
    .B1(_1600_),
    .X(_1618_));
 sky130_fd_sc_hd__or2_1 _4671_ (.A(_1598_),
    .B(_1618_),
    .X(_1619_));
 sky130_fd_sc_hd__and2b_1 _4672_ (.A_N(_1355_),
    .B(\core_1.execute.alu_mul_div.div_cur[8] ),
    .X(_1620_));
 sky130_fd_sc_hd__and2b_1 _4673_ (.A_N(\core_1.execute.alu_mul_div.div_cur[8] ),
    .B(_1355_),
    .X(_1621_));
 sky130_fd_sc_hd__nor2_1 _4674_ (.A(_1620_),
    .B(_1621_),
    .Y(_1622_));
 sky130_fd_sc_hd__a31o_1 _4675_ (.A1(_1597_),
    .A2(_1619_),
    .A3(_1622_),
    .B1(_1620_),
    .X(_1623_));
 sky130_fd_sc_hd__and2b_1 _4676_ (.A_N(_1354_),
    .B(\core_1.execute.alu_mul_div.div_cur[9] ),
    .X(_1624_));
 sky130_fd_sc_hd__a21o_1 _4677_ (.A1(_1595_),
    .A2(_1623_),
    .B1(_1624_),
    .X(_1625_));
 sky130_fd_sc_hd__a21o_1 _4678_ (.A1(_1594_),
    .A2(_1625_),
    .B1(_1592_),
    .X(_1626_));
 sky130_fd_sc_hd__and2_1 _4679_ (.A(\core_1.execute.alu_mul_div.div_cur[11] ),
    .B(_1589_),
    .X(_1627_));
 sky130_fd_sc_hd__a21oi_1 _4680_ (.A1(_1590_),
    .A2(_1626_),
    .B1(_1627_),
    .Y(_1628_));
 sky130_fd_sc_hd__xnor2_1 _4681_ (.A(\core_1.execute.alu_mul_div.div_cur[12] ),
    .B(_1373_),
    .Y(_1629_));
 sky130_fd_sc_hd__and2b_1 _4682_ (.A_N(_1628_),
    .B(_1629_),
    .X(_1630_));
 sky130_fd_sc_hd__a21o_1 _4683_ (.A1(\core_1.execute.alu_mul_div.div_cur[12] ),
    .A2(_1587_),
    .B1(_1630_),
    .X(_1631_));
 sky130_fd_sc_hd__or2_1 _4684_ (.A(\core_1.execute.alu_mul_div.div_cur[13] ),
    .B(_1585_),
    .X(_1632_));
 sky130_fd_sc_hd__o21ai_2 _4685_ (.A1(_1586_),
    .A2(_1631_),
    .B1(_1632_),
    .Y(_1633_));
 sky130_fd_sc_hd__or2b_1 _4686_ (.A(_1351_),
    .B_N(\core_1.execute.alu_mul_div.div_cur[14] ),
    .X(_1634_));
 sky130_fd_sc_hd__o21a_1 _4687_ (.A1(_1584_),
    .A2(_1633_),
    .B1(_1634_),
    .X(_1635_));
 sky130_fd_sc_hd__nand2_1 _4688_ (.A(\core_1.execute.alu_mul_div.div_cur[15] ),
    .B(_1358_),
    .Y(_1636_));
 sky130_fd_sc_hd__o21ai_4 _4689_ (.A1(_1583_),
    .A2(_1635_),
    .B1(_1636_),
    .Y(_1637_));
 sky130_fd_sc_hd__and2_1 _4690_ (.A(\core_1.execute.alu_mul_div.comp ),
    .B(_1314_),
    .X(_1638_));
 sky130_fd_sc_hd__o21a_2 _4691_ (.A1(_1196_),
    .A2(_1637_),
    .B1(_1638_),
    .X(_1639_));
 sky130_fd_sc_hd__clkbuf_4 _4692_ (.A(_1639_),
    .X(_1640_));
 sky130_fd_sc_hd__o21a_4 _4693_ (.A1(_1583_),
    .A2(_1635_),
    .B1(_1636_),
    .X(_1641_));
 sky130_fd_sc_hd__o21ai_4 _4694_ (.A1(_1197_),
    .A2(_1637_),
    .B1(_1638_),
    .Y(_1642_));
 sky130_fd_sc_hd__clkbuf_4 _4695_ (.A(_1642_),
    .X(_1643_));
 sky130_fd_sc_hd__and2b_1 _4696_ (.A_N(_1611_),
    .B(_1609_),
    .X(_1644_));
 sky130_fd_sc_hd__nor2_1 _4697_ (.A(\core_1.execute.alu_mul_div.div_cur[0] ),
    .B(_1407_),
    .Y(_1645_));
 sky130_fd_sc_hd__xnor2_2 _4698_ (.A(_1644_),
    .B(_1645_),
    .Y(_1646_));
 sky130_fd_sc_hd__and3_1 _4699_ (.A(\core_1.execute.alu_mul_div.div_cur[0] ),
    .B(_1326_),
    .C(_1327_),
    .X(_1647_));
 sky130_fd_sc_hd__nor2_1 _4700_ (.A(_1645_),
    .B(_1647_),
    .Y(_1648_));
 sky130_fd_sc_hd__nand2_1 _4701_ (.A(_1197_),
    .B(_1648_),
    .Y(_1649_));
 sky130_fd_sc_hd__clkbuf_4 _4702_ (.A(_1637_),
    .X(_1650_));
 sky130_fd_sc_hd__o211a_1 _4703_ (.A1(_1197_),
    .A2(_1646_),
    .B1(_1649_),
    .C1(_1650_),
    .X(_1651_));
 sky130_fd_sc_hd__a211o_1 _4704_ (.A1(\core_1.execute.alu_mul_div.div_cur[0] ),
    .A2(_1641_),
    .B1(_1643_),
    .C1(_1651_),
    .X(_1652_));
 sky130_fd_sc_hd__buf_2 _4705_ (.A(_0728_),
    .X(_1653_));
 sky130_fd_sc_hd__clkbuf_4 _4706_ (.A(_1653_),
    .X(_1654_));
 sky130_fd_sc_hd__o211a_1 _4707_ (.A1(\core_1.execute.alu_mul_div.div_cur[1] ),
    .A2(_1640_),
    .B1(_1652_),
    .C1(_1654_),
    .X(_0172_));
 sky130_fd_sc_hd__and2_1 _4708_ (.A(_1188_),
    .B(_1195_),
    .X(_1655_));
 sky130_fd_sc_hd__buf_2 _4709_ (.A(_1655_),
    .X(_1656_));
 sky130_fd_sc_hd__and2_1 _4710_ (.A(_1608_),
    .B(_1612_),
    .X(_1657_));
 sky130_fd_sc_hd__nor2_1 _4711_ (.A(_1608_),
    .B(_1612_),
    .Y(_1658_));
 sky130_fd_sc_hd__nor2_1 _4712_ (.A(_1657_),
    .B(_1658_),
    .Y(_1659_));
 sky130_fd_sc_hd__or2_1 _4713_ (.A(_1196_),
    .B(_1659_),
    .X(_1660_));
 sky130_fd_sc_hd__o211a_1 _4714_ (.A1(_1656_),
    .A2(_1646_),
    .B1(_1660_),
    .C1(_1650_),
    .X(_1661_));
 sky130_fd_sc_hd__a211o_1 _4715_ (.A1(\core_1.execute.alu_mul_div.div_cur[1] ),
    .A2(_1641_),
    .B1(_1643_),
    .C1(_1661_),
    .X(_1662_));
 sky130_fd_sc_hd__o211a_1 _4716_ (.A1(\core_1.execute.alu_mul_div.div_cur[2] ),
    .A2(_1640_),
    .B1(_1662_),
    .C1(_1654_),
    .X(_0173_));
 sky130_fd_sc_hd__or2_1 _4717_ (.A(_1614_),
    .B(_1657_),
    .X(_1663_));
 sky130_fd_sc_hd__nor2_1 _4718_ (.A(\core_1.execute.alu_mul_div.div_cur[3] ),
    .B(_1504_),
    .Y(_1664_));
 sky130_fd_sc_hd__nor2_1 _4719_ (.A(_1664_),
    .B(_1613_),
    .Y(_1665_));
 sky130_fd_sc_hd__xor2_2 _4720_ (.A(_1663_),
    .B(_1665_),
    .X(_1666_));
 sky130_fd_sc_hd__or2_1 _4721_ (.A(_1656_),
    .B(_1659_),
    .X(_1667_));
 sky130_fd_sc_hd__o211a_1 _4722_ (.A1(_1197_),
    .A2(_1666_),
    .B1(_1667_),
    .C1(_1650_),
    .X(_1668_));
 sky130_fd_sc_hd__a211o_1 _4723_ (.A1(\core_1.execute.alu_mul_div.div_cur[2] ),
    .A2(_1641_),
    .B1(_1643_),
    .C1(_1668_),
    .X(_1669_));
 sky130_fd_sc_hd__o211a_1 _4724_ (.A1(\core_1.execute.alu_mul_div.div_cur[3] ),
    .A2(_1640_),
    .B1(_1669_),
    .C1(_1654_),
    .X(_0174_));
 sky130_fd_sc_hd__and3_1 _4725_ (.A(_1606_),
    .B(_1607_),
    .C(_1615_),
    .X(_1670_));
 sky130_fd_sc_hd__a21oi_1 _4726_ (.A1(_1607_),
    .A2(_1615_),
    .B1(_1606_),
    .Y(_1671_));
 sky130_fd_sc_hd__nor2_1 _4727_ (.A(_1670_),
    .B(_1671_),
    .Y(_1672_));
 sky130_fd_sc_hd__or2_1 _4728_ (.A(_1196_),
    .B(_1672_),
    .X(_1673_));
 sky130_fd_sc_hd__o211a_1 _4729_ (.A1(_1656_),
    .A2(_1666_),
    .B1(_1673_),
    .C1(_1650_),
    .X(_1674_));
 sky130_fd_sc_hd__a211o_1 _4730_ (.A1(\core_1.execute.alu_mul_div.div_cur[3] ),
    .A2(_1641_),
    .B1(_1643_),
    .C1(_1674_),
    .X(_1675_));
 sky130_fd_sc_hd__o211a_1 _4731_ (.A1(\core_1.execute.alu_mul_div.div_cur[4] ),
    .A2(_1640_),
    .B1(_1675_),
    .C1(_1654_),
    .X(_0175_));
 sky130_fd_sc_hd__or2_1 _4732_ (.A(_1604_),
    .B(_1670_),
    .X(_1676_));
 sky130_fd_sc_hd__or2b_1 _4733_ (.A(_1616_),
    .B_N(_1603_),
    .X(_1677_));
 sky130_fd_sc_hd__xnor2_1 _4734_ (.A(_1676_),
    .B(_1677_),
    .Y(_1678_));
 sky130_fd_sc_hd__or2_1 _4735_ (.A(_1656_),
    .B(_1672_),
    .X(_1679_));
 sky130_fd_sc_hd__o211a_1 _4736_ (.A1(_1197_),
    .A2(_1678_),
    .B1(_1679_),
    .C1(_1650_),
    .X(_1680_));
 sky130_fd_sc_hd__a211o_1 _4737_ (.A1(\core_1.execute.alu_mul_div.div_cur[4] ),
    .A2(_1641_),
    .B1(_1643_),
    .C1(_1680_),
    .X(_1681_));
 sky130_fd_sc_hd__o211a_1 _4738_ (.A1(\core_1.execute.alu_mul_div.div_cur[5] ),
    .A2(_1640_),
    .B1(_1681_),
    .C1(_1654_),
    .X(_0176_));
 sky130_fd_sc_hd__nand2_1 _4739_ (.A(_1603_),
    .B(_1617_),
    .Y(_1682_));
 sky130_fd_sc_hd__xnor2_1 _4740_ (.A(_1602_),
    .B(_1682_),
    .Y(_1683_));
 sky130_fd_sc_hd__mux2_1 _4741_ (.A0(_1678_),
    .A1(_1683_),
    .S(_1656_),
    .X(_1684_));
 sky130_fd_sc_hd__mux2_1 _4742_ (.A0(\core_1.execute.alu_mul_div.div_cur[5] ),
    .A1(_1684_),
    .S(_1650_),
    .X(_1685_));
 sky130_fd_sc_hd__or2_1 _4743_ (.A(_1643_),
    .B(_1685_),
    .X(_1686_));
 sky130_fd_sc_hd__clkbuf_4 _4744_ (.A(_1653_),
    .X(_1687_));
 sky130_fd_sc_hd__o211a_1 _4745_ (.A1(\core_1.execute.alu_mul_div.div_cur[6] ),
    .A2(_1640_),
    .B1(_1686_),
    .C1(_1687_),
    .X(_0177_));
 sky130_fd_sc_hd__inv_2 _4746_ (.A(_1597_),
    .Y(_1688_));
 sky130_fd_sc_hd__nor2_1 _4747_ (.A(_1688_),
    .B(_1598_),
    .Y(_1689_));
 sky130_fd_sc_hd__xor2_1 _4748_ (.A(_1618_),
    .B(_1689_),
    .X(_1690_));
 sky130_fd_sc_hd__mux2_1 _4749_ (.A0(_1683_),
    .A1(_1690_),
    .S(_1656_),
    .X(_1691_));
 sky130_fd_sc_hd__mux2_1 _4750_ (.A0(\core_1.execute.alu_mul_div.div_cur[6] ),
    .A1(_1691_),
    .S(_1650_),
    .X(_1692_));
 sky130_fd_sc_hd__or2_1 _4751_ (.A(_1642_),
    .B(_1692_),
    .X(_1693_));
 sky130_fd_sc_hd__o211a_1 _4752_ (.A1(\core_1.execute.alu_mul_div.div_cur[7] ),
    .A2(_1640_),
    .B1(_1693_),
    .C1(_1687_),
    .X(_0178_));
 sky130_fd_sc_hd__nand2_1 _4753_ (.A(_1597_),
    .B(_1619_),
    .Y(_1694_));
 sky130_fd_sc_hd__xnor2_1 _4754_ (.A(_1694_),
    .B(_1622_),
    .Y(_1695_));
 sky130_fd_sc_hd__or2_1 _4755_ (.A(_1196_),
    .B(_1695_),
    .X(_1696_));
 sky130_fd_sc_hd__o211a_1 _4756_ (.A1(_1656_),
    .A2(_1690_),
    .B1(_1696_),
    .C1(_1650_),
    .X(_1697_));
 sky130_fd_sc_hd__a211o_1 _4757_ (.A1(\core_1.execute.alu_mul_div.div_cur[7] ),
    .A2(_1641_),
    .B1(_1643_),
    .C1(_1697_),
    .X(_1698_));
 sky130_fd_sc_hd__o211a_1 _4758_ (.A1(\core_1.execute.alu_mul_div.div_cur[8] ),
    .A2(_1640_),
    .B1(_1698_),
    .C1(_1687_),
    .X(_0179_));
 sky130_fd_sc_hd__and2b_1 _4759_ (.A_N(_1624_),
    .B(_1595_),
    .X(_1699_));
 sky130_fd_sc_hd__xor2_1 _4760_ (.A(_1623_),
    .B(_1699_),
    .X(_1700_));
 sky130_fd_sc_hd__mux2_1 _4761_ (.A0(_1695_),
    .A1(_1700_),
    .S(_1656_),
    .X(_1701_));
 sky130_fd_sc_hd__mux2_1 _4762_ (.A0(\core_1.execute.alu_mul_div.div_cur[8] ),
    .A1(_1701_),
    .S(_1637_),
    .X(_1702_));
 sky130_fd_sc_hd__or2_1 _4763_ (.A(_1642_),
    .B(_1702_),
    .X(_1703_));
 sky130_fd_sc_hd__o211a_1 _4764_ (.A1(\core_1.execute.alu_mul_div.div_cur[9] ),
    .A2(_1640_),
    .B1(_1703_),
    .C1(_1687_),
    .X(_0180_));
 sky130_fd_sc_hd__xor2_1 _4765_ (.A(_1594_),
    .B(_1625_),
    .X(_1704_));
 sky130_fd_sc_hd__or2_1 _4766_ (.A(_1196_),
    .B(_1704_),
    .X(_1705_));
 sky130_fd_sc_hd__o211a_1 _4767_ (.A1(_1656_),
    .A2(_1700_),
    .B1(_1705_),
    .C1(_1650_),
    .X(_1706_));
 sky130_fd_sc_hd__a211o_1 _4768_ (.A1(\core_1.execute.alu_mul_div.div_cur[9] ),
    .A2(_1641_),
    .B1(_1643_),
    .C1(_1706_),
    .X(_1707_));
 sky130_fd_sc_hd__o211a_1 _4769_ (.A1(\core_1.execute.alu_mul_div.div_cur[10] ),
    .A2(_1640_),
    .B1(_1707_),
    .C1(_1687_),
    .X(_0181_));
 sky130_fd_sc_hd__or2b_1 _4770_ (.A(_1627_),
    .B_N(_1590_),
    .X(_1708_));
 sky130_fd_sc_hd__xnor2_1 _4771_ (.A(_1626_),
    .B(_1708_),
    .Y(_1709_));
 sky130_fd_sc_hd__mux2_1 _4772_ (.A0(_1704_),
    .A1(_1709_),
    .S(_1655_),
    .X(_1710_));
 sky130_fd_sc_hd__mux2_1 _4773_ (.A0(\core_1.execute.alu_mul_div.div_cur[10] ),
    .A1(_1710_),
    .S(_1637_),
    .X(_1711_));
 sky130_fd_sc_hd__or2_1 _4774_ (.A(_1642_),
    .B(_1711_),
    .X(_1712_));
 sky130_fd_sc_hd__o211a_1 _4775_ (.A1(\core_1.execute.alu_mul_div.div_cur[11] ),
    .A2(_1639_),
    .B1(_1712_),
    .C1(_1687_),
    .X(_0182_));
 sky130_fd_sc_hd__xnor2_1 _4776_ (.A(_1629_),
    .B(_1628_),
    .Y(_1713_));
 sky130_fd_sc_hd__mux2_1 _4777_ (.A0(_1709_),
    .A1(_1713_),
    .S(_1655_),
    .X(_1714_));
 sky130_fd_sc_hd__mux2_1 _4778_ (.A0(\core_1.execute.alu_mul_div.div_cur[11] ),
    .A1(_1714_),
    .S(_1637_),
    .X(_1715_));
 sky130_fd_sc_hd__or2_1 _4779_ (.A(_1642_),
    .B(_1715_),
    .X(_1716_));
 sky130_fd_sc_hd__o211a_1 _4780_ (.A1(\core_1.execute.alu_mul_div.div_cur[12] ),
    .A2(_1639_),
    .B1(_1716_),
    .C1(_1687_),
    .X(_0183_));
 sky130_fd_sc_hd__nor2_1 _4781_ (.A(\core_1.execute.alu_mul_div.div_cur[13] ),
    .B(_1585_),
    .Y(_1717_));
 sky130_fd_sc_hd__or2_1 _4782_ (.A(_1717_),
    .B(_1586_),
    .X(_1718_));
 sky130_fd_sc_hd__xnor2_1 _4783_ (.A(_1631_),
    .B(_1718_),
    .Y(_1719_));
 sky130_fd_sc_hd__or2_1 _4784_ (.A(_1656_),
    .B(_1713_),
    .X(_1720_));
 sky130_fd_sc_hd__o211a_1 _4785_ (.A1(_1197_),
    .A2(_1719_),
    .B1(_1720_),
    .C1(_1650_),
    .X(_1721_));
 sky130_fd_sc_hd__a211o_1 _4786_ (.A1(\core_1.execute.alu_mul_div.div_cur[12] ),
    .A2(_1641_),
    .B1(_1643_),
    .C1(_1721_),
    .X(_1722_));
 sky130_fd_sc_hd__o211a_1 _4787_ (.A1(\core_1.execute.alu_mul_div.div_cur[13] ),
    .A2(_1639_),
    .B1(_1722_),
    .C1(_1687_),
    .X(_0184_));
 sky130_fd_sc_hd__and2b_1 _4788_ (.A_N(_1351_),
    .B(\core_1.execute.alu_mul_div.div_cur[14] ),
    .X(_1723_));
 sky130_fd_sc_hd__nor2_1 _4789_ (.A(_1723_),
    .B(_1584_),
    .Y(_1724_));
 sky130_fd_sc_hd__xnor2_1 _4790_ (.A(_1724_),
    .B(_1633_),
    .Y(_1725_));
 sky130_fd_sc_hd__mux2_1 _4791_ (.A0(_1719_),
    .A1(_1725_),
    .S(_1655_),
    .X(_1726_));
 sky130_fd_sc_hd__mux2_1 _4792_ (.A0(\core_1.execute.alu_mul_div.div_cur[13] ),
    .A1(_1726_),
    .S(_1637_),
    .X(_1727_));
 sky130_fd_sc_hd__or2_1 _4793_ (.A(_1642_),
    .B(_1727_),
    .X(_1728_));
 sky130_fd_sc_hd__o211a_1 _4794_ (.A1(\core_1.execute.alu_mul_div.div_cur[14] ),
    .A2(_1639_),
    .B1(_1728_),
    .C1(_1687_),
    .X(_0185_));
 sky130_fd_sc_hd__nand2_1 _4795_ (.A(_1197_),
    .B(_1725_),
    .Y(_1729_));
 sky130_fd_sc_hd__or3_1 _4796_ (.A(_1196_),
    .B(_1636_),
    .C(_1635_),
    .X(_1730_));
 sky130_fd_sc_hd__a21oi_1 _4797_ (.A1(_1729_),
    .A2(_1730_),
    .B1(_1641_),
    .Y(_1731_));
 sky130_fd_sc_hd__a211o_1 _4798_ (.A1(\core_1.execute.alu_mul_div.div_cur[14] ),
    .A2(_1641_),
    .B1(_1643_),
    .C1(_1731_),
    .X(_1732_));
 sky130_fd_sc_hd__o211a_1 _4799_ (.A1(\core_1.execute.alu_mul_div.div_cur[15] ),
    .A2(_1639_),
    .B1(_1732_),
    .C1(_1687_),
    .X(_0186_));
 sky130_fd_sc_hd__o21a_4 _4800_ (.A1(net94),
    .A2(_1377_),
    .B1(_1388_),
    .X(_1733_));
 sky130_fd_sc_hd__o22a_4 _4801_ (.A1(net90),
    .A2(_1377_),
    .B1(_1480_),
    .B2(_1483_),
    .X(_1734_));
 sky130_fd_sc_hd__mux2_1 _4802_ (.A0(_1477_),
    .A1(_1734_),
    .S(_1192_),
    .X(_1735_));
 sky130_fd_sc_hd__clkinv_2 _4803_ (.A(\core_1.execute.alu_mul_div.cbit[0] ),
    .Y(_1736_));
 sky130_fd_sc_hd__buf_4 _4804_ (.A(_1736_),
    .X(_1737_));
 sky130_fd_sc_hd__nor2_4 _4805_ (.A(_1737_),
    .B(_1193_),
    .Y(_1738_));
 sky130_fd_sc_hd__a22o_1 _4806_ (.A1(_1193_),
    .A2(_1735_),
    .B1(_1738_),
    .B2(_1493_),
    .X(_1739_));
 sky130_fd_sc_hd__and2_1 _4807_ (.A(_1191_),
    .B(_1739_),
    .X(_1740_));
 sky130_fd_sc_hd__clkbuf_4 _4808_ (.A(\core_1.execute.alu_mul_div.cbit[2] ),
    .X(_1741_));
 sky130_fd_sc_hd__or2_1 _4809_ (.A(\core_1.execute.alu_mul_div.cbit[0] ),
    .B(\core_1.execute.alu_mul_div.cbit[1] ),
    .X(_1742_));
 sky130_fd_sc_hd__clkbuf_4 _4810_ (.A(_1742_),
    .X(_1743_));
 sky130_fd_sc_hd__nor2_2 _4811_ (.A(_1741_),
    .B(_1743_),
    .Y(_1744_));
 sky130_fd_sc_hd__o21a_4 _4812_ (.A1(net93),
    .A2(_1377_),
    .B1(_1499_),
    .X(_1745_));
 sky130_fd_sc_hd__o22a_4 _4813_ (.A1(net102),
    .A2(_1376_),
    .B1(_1533_),
    .B2(_1536_),
    .X(_1746_));
 sky130_fd_sc_hd__mux4_1 _4814_ (.A0(_1457_),
    .A1(_1465_),
    .A2(_1746_),
    .A3(_1531_),
    .S0(_1192_),
    .S1(_1193_),
    .X(_1747_));
 sky130_fd_sc_hd__a221o_1 _4815_ (.A1(_1744_),
    .A2(_1745_),
    .B1(_1747_),
    .B2(_1741_),
    .C1(_1188_),
    .X(_1748_));
 sky130_fd_sc_hd__mux4_2 _4816_ (.A0(_1515_),
    .A1(_1523_),
    .A2(_1547_),
    .A3(_1553_),
    .S0(_1192_),
    .S1(_1193_),
    .X(_1749_));
 sky130_fd_sc_hd__mux2_1 _4817_ (.A0(_1403_),
    .A1(_1562_),
    .S(_1737_),
    .X(_1750_));
 sky130_fd_sc_hd__inv_2 _4818_ (.A(\core_1.execute.alu_mul_div.cbit[1] ),
    .Y(_1751_));
 sky130_fd_sc_hd__nor2_2 _4819_ (.A(\core_1.execute.alu_mul_div.cbit[0] ),
    .B(_1751_),
    .Y(_1752_));
 sky130_fd_sc_hd__a2bb2o_1 _4820_ (.A1_N(\core_1.execute.alu_mul_div.cbit[1] ),
    .A2_N(_1750_),
    .B1(_1752_),
    .B2(_1346_),
    .X(_1753_));
 sky130_fd_sc_hd__inv_2 _4821_ (.A(_1753_),
    .Y(_1754_));
 sky130_fd_sc_hd__mux2_1 _4822_ (.A0(_1749_),
    .A1(_1754_),
    .S(\core_1.execute.alu_mul_div.cbit[2] ),
    .X(_1755_));
 sky130_fd_sc_hd__a2bb2o_2 _4823_ (.A1_N(_1740_),
    .A2_N(_1748_),
    .B1(_1755_),
    .B2(_1188_),
    .X(_1756_));
 sky130_fd_sc_hd__o21ai_1 _4824_ (.A1(_1197_),
    .A2(_1648_),
    .B1(_1756_),
    .Y(_1757_));
 sky130_fd_sc_hd__mux2_1 _4825_ (.A0(\core_1.execute.alu_mul_div.div_cur[0] ),
    .A1(_1757_),
    .S(_1639_),
    .X(_1758_));
 sky130_fd_sc_hd__mux2_1 _4826_ (.A0(_1733_),
    .A1(_1758_),
    .S(_1653_),
    .X(_1759_));
 sky130_fd_sc_hd__clkbuf_1 _4827_ (.A(_1759_),
    .X(_0187_));
 sky130_fd_sc_hd__or4b_4 _4828_ (.A(\core_1.decode.i_flush ),
    .B(_0659_),
    .C(_0688_),
    .D_N(_0731_),
    .X(_1760_));
 sky130_fd_sc_hd__nor2_1 _4829_ (.A(_0730_),
    .B(_1760_),
    .Y(_1761_));
 sky130_fd_sc_hd__and2_1 _4830_ (.A(_1193_),
    .B(_1760_),
    .X(_1762_));
 sky130_fd_sc_hd__a31o_1 _4831_ (.A1(_1194_),
    .A2(_1743_),
    .A3(_1761_),
    .B1(_1762_),
    .X(_0188_));
 sky130_fd_sc_hd__buf_2 _4832_ (.A(_1741_),
    .X(_1763_));
 sky130_fd_sc_hd__clkbuf_4 _4833_ (.A(_1751_),
    .X(_1764_));
 sky130_fd_sc_hd__nor2_2 _4834_ (.A(_1737_),
    .B(_1764_),
    .Y(_1765_));
 sky130_fd_sc_hd__nor2_1 _4835_ (.A(_1763_),
    .B(_1765_),
    .Y(_1766_));
 sky130_fd_sc_hd__or4_1 _4836_ (.A(_0730_),
    .B(_1198_),
    .C(_1195_),
    .D(_1766_),
    .X(_1767_));
 sky130_fd_sc_hd__a21bo_1 _4837_ (.A1(_1763_),
    .A2(_1760_),
    .B1_N(_1767_),
    .X(_0189_));
 sky130_fd_sc_hd__inv_2 _4838_ (.A(\core_1.execute.alu_mul_div.cbit[3] ),
    .Y(_1768_));
 sky130_fd_sc_hd__buf_4 _4839_ (.A(_1768_),
    .X(_1769_));
 sky130_fd_sc_hd__xnor2_1 _4840_ (.A(_1769_),
    .B(_1195_),
    .Y(_1770_));
 sky130_fd_sc_hd__a22o_1 _4841_ (.A1(_1188_),
    .A2(_1760_),
    .B1(_1761_),
    .B2(_1770_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _4842_ (.A0(\core_1.dec_mem_long ),
    .A1(_0806_),
    .S(_0811_),
    .X(_1771_));
 sky130_fd_sc_hd__clkbuf_1 _4843_ (.A(_1771_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _4844_ (.A0(\core_1.execute.sreg_data_page ),
    .A1(net104),
    .S(_0726_),
    .X(_1772_));
 sky130_fd_sc_hd__and2_1 _4845_ (.A(_1178_),
    .B(_1772_),
    .X(_1773_));
 sky130_fd_sc_hd__clkbuf_1 _4846_ (.A(_1773_),
    .X(_0192_));
 sky130_fd_sc_hd__clkinv_2 _4847_ (.A(_1043_),
    .Y(_1774_));
 sky130_fd_sc_hd__or2_1 _4848_ (.A(net72),
    .B(_1043_),
    .X(_1775_));
 sky130_fd_sc_hd__clkbuf_4 _4849_ (.A(_1155_),
    .X(_1776_));
 sky130_fd_sc_hd__o211a_1 _4850_ (.A1(\core_1.execute.mem_stage_pc[0] ),
    .A2(_1774_),
    .B1(_1775_),
    .C1(_1776_),
    .X(_0193_));
 sky130_fd_sc_hd__buf_6 _4851_ (.A(_0733_),
    .X(_1777_));
 sky130_fd_sc_hd__buf_4 _4852_ (.A(_1777_),
    .X(_1778_));
 sky130_fd_sc_hd__or2_1 _4853_ (.A(\core_1.execute.mem_stage_pc[1] ),
    .B(_1007_),
    .X(_1779_));
 sky130_fd_sc_hd__o211a_1 _4854_ (.A1(net79),
    .A2(_1778_),
    .B1(_1779_),
    .C1(_1776_),
    .X(_0194_));
 sky130_fd_sc_hd__or2_1 _4855_ (.A(\core_1.execute.mem_stage_pc[2] ),
    .B(_1007_),
    .X(_1780_));
 sky130_fd_sc_hd__o211a_1 _4856_ (.A1(net80),
    .A2(_1778_),
    .B1(_1780_),
    .C1(_1776_),
    .X(_0195_));
 sky130_fd_sc_hd__or2_1 _4857_ (.A(\core_1.execute.mem_stage_pc[3] ),
    .B(_1007_),
    .X(_1781_));
 sky130_fd_sc_hd__o211a_1 _4858_ (.A1(net81),
    .A2(_1778_),
    .B1(_1781_),
    .C1(_1776_),
    .X(_0196_));
 sky130_fd_sc_hd__or2_1 _4859_ (.A(\core_1.execute.mem_stage_pc[4] ),
    .B(_1007_),
    .X(_1782_));
 sky130_fd_sc_hd__o211a_1 _4860_ (.A1(net82),
    .A2(_1778_),
    .B1(_1782_),
    .C1(_1776_),
    .X(_0197_));
 sky130_fd_sc_hd__or2_1 _4861_ (.A(\core_1.execute.mem_stage_pc[5] ),
    .B(_1007_),
    .X(_1783_));
 sky130_fd_sc_hd__o211a_1 _4862_ (.A1(net83),
    .A2(_1778_),
    .B1(_1783_),
    .C1(_1776_),
    .X(_0198_));
 sky130_fd_sc_hd__or2_1 _4863_ (.A(\core_1.execute.mem_stage_pc[6] ),
    .B(_1007_),
    .X(_1784_));
 sky130_fd_sc_hd__o211a_1 _4864_ (.A1(net84),
    .A2(_1778_),
    .B1(_1784_),
    .C1(_1776_),
    .X(_0199_));
 sky130_fd_sc_hd__or2_1 _4865_ (.A(\core_1.execute.mem_stage_pc[7] ),
    .B(_1007_),
    .X(_1785_));
 sky130_fd_sc_hd__o211a_1 _4866_ (.A1(net85),
    .A2(_1778_),
    .B1(_1785_),
    .C1(_1776_),
    .X(_0200_));
 sky130_fd_sc_hd__or2_1 _4867_ (.A(\core_1.execute.mem_stage_pc[8] ),
    .B(_1007_),
    .X(_1786_));
 sky130_fd_sc_hd__o211a_1 _4868_ (.A1(net86),
    .A2(_1778_),
    .B1(_1786_),
    .C1(_1776_),
    .X(_0201_));
 sky130_fd_sc_hd__or2_1 _4869_ (.A(\core_1.execute.mem_stage_pc[9] ),
    .B(_1007_),
    .X(_1787_));
 sky130_fd_sc_hd__clkbuf_4 _4870_ (.A(_1155_),
    .X(_1788_));
 sky130_fd_sc_hd__clkbuf_8 _4871_ (.A(_1788_),
    .X(_1789_));
 sky130_fd_sc_hd__o211a_1 _4872_ (.A1(net87),
    .A2(_1778_),
    .B1(_1787_),
    .C1(_1789_),
    .X(_0202_));
 sky130_fd_sc_hd__or2_1 _4873_ (.A(\core_1.execute.mem_stage_pc[10] ),
    .B(_1006_),
    .X(_1790_));
 sky130_fd_sc_hd__o211a_1 _4874_ (.A1(net73),
    .A2(_1778_),
    .B1(_1790_),
    .C1(_1789_),
    .X(_0203_));
 sky130_fd_sc_hd__or2_1 _4875_ (.A(\core_1.execute.mem_stage_pc[11] ),
    .B(_1006_),
    .X(_1791_));
 sky130_fd_sc_hd__o211a_1 _4876_ (.A1(net74),
    .A2(_1777_),
    .B1(_1791_),
    .C1(_1789_),
    .X(_0204_));
 sky130_fd_sc_hd__or2_1 _4877_ (.A(\core_1.execute.mem_stage_pc[12] ),
    .B(_1006_),
    .X(_1792_));
 sky130_fd_sc_hd__o211a_1 _4878_ (.A1(net75),
    .A2(_1777_),
    .B1(_1792_),
    .C1(_1789_),
    .X(_0205_));
 sky130_fd_sc_hd__or2_1 _4879_ (.A(\core_1.execute.mem_stage_pc[13] ),
    .B(_1006_),
    .X(_1793_));
 sky130_fd_sc_hd__o211a_1 _4880_ (.A1(net76),
    .A2(_1777_),
    .B1(_1793_),
    .C1(_1789_),
    .X(_0206_));
 sky130_fd_sc_hd__or2_1 _4881_ (.A(\core_1.execute.mem_stage_pc[14] ),
    .B(_1006_),
    .X(_1794_));
 sky130_fd_sc_hd__o211a_1 _4882_ (.A1(net77),
    .A2(_1777_),
    .B1(_1794_),
    .C1(_1789_),
    .X(_0207_));
 sky130_fd_sc_hd__or2_1 _4883_ (.A(\core_1.execute.mem_stage_pc[15] ),
    .B(_1006_),
    .X(_1795_));
 sky130_fd_sc_hd__o211a_1 _4884_ (.A1(net78),
    .A2(_1777_),
    .B1(_1795_),
    .C1(_1789_),
    .X(_0208_));
 sky130_fd_sc_hd__nor2_1 _4885_ (.A(_1056_),
    .B(_0684_),
    .Y(_0209_));
 sky130_fd_sc_hd__nor2_1 _4886_ (.A(_1056_),
    .B(_0674_),
    .Y(_0210_));
 sky130_fd_sc_hd__nor2_1 _4887_ (.A(_1056_),
    .B(_0672_),
    .Y(_0211_));
 sky130_fd_sc_hd__nor2_1 _4888_ (.A(_1056_),
    .B(_0669_),
    .Y(_0212_));
 sky130_fd_sc_hd__nor2_1 _4889_ (.A(_1056_),
    .B(_0680_),
    .Y(_0213_));
 sky130_fd_sc_hd__nor2_1 _4890_ (.A(_1056_),
    .B(_0677_),
    .Y(_0214_));
 sky130_fd_sc_hd__nor2_1 _4891_ (.A(_1056_),
    .B(_0671_),
    .Y(_0215_));
 sky130_fd_sc_hd__nor2_1 _4892_ (.A(_1165_),
    .B(_0675_),
    .Y(_0216_));
 sky130_fd_sc_hd__or2_2 _4893_ (.A(_0659_),
    .B(_1777_),
    .X(_1796_));
 sky130_fd_sc_hd__inv_2 _4894_ (.A(_1796_),
    .Y(_0228_));
 sky130_fd_sc_hd__and2_1 _4895_ (.A(\core_1.execute.trap_flag ),
    .B(_0228_),
    .X(_1797_));
 sky130_fd_sc_hd__clkbuf_1 _4896_ (.A(_1797_),
    .X(_0217_));
 sky130_fd_sc_hd__and2_1 _4897_ (.A(\core_1.dec_sys ),
    .B(_0228_),
    .X(_1798_));
 sky130_fd_sc_hd__clkbuf_1 _4898_ (.A(_1798_),
    .X(_0218_));
 sky130_fd_sc_hd__and2_1 _4899_ (.A(_1154_),
    .B(_1006_),
    .X(_1799_));
 sky130_fd_sc_hd__buf_2 _4900_ (.A(_1799_),
    .X(_1800_));
 sky130_fd_sc_hd__buf_6 _4901_ (.A(_1800_),
    .X(_1801_));
 sky130_fd_sc_hd__mux2_1 _4902_ (.A0(net159),
    .A1(\core_1.dec_mem_we ),
    .S(_1801_),
    .X(_1802_));
 sky130_fd_sc_hd__clkbuf_1 _4903_ (.A(_1802_),
    .X(_0219_));
 sky130_fd_sc_hd__a2111o_4 _4904_ (.A1(\core_1.execute.rf.reg_outputs[1][0] ),
    .A2(_1459_),
    .B1(_1332_),
    .C1(_1333_),
    .D1(_1334_),
    .X(_1803_));
 sky130_fd_sc_hd__mux2_4 _4905_ (.A0(net184),
    .A1(net200),
    .S(_1350_),
    .X(_1804_));
 sky130_fd_sc_hd__a21oi_1 _4906_ (.A1(_1364_),
    .A2(_1414_),
    .B1(_1369_),
    .Y(_1805_));
 sky130_fd_sc_hd__o21ai_1 _4907_ (.A1(_1363_),
    .A2(_1805_),
    .B1(\core_1.decode.oc_alu_mode[13] ),
    .Y(_1806_));
 sky130_fd_sc_hd__a21oi_1 _4908_ (.A1(_1363_),
    .A2(_1805_),
    .B1(_1806_),
    .Y(_1807_));
 sky130_fd_sc_hd__o21ai_1 _4909_ (.A1(_0822_),
    .A2(_1531_),
    .B1(_1393_),
    .Y(_1808_));
 sky130_fd_sc_hd__o21ai_1 _4910_ (.A1(_1331_),
    .A2(_1746_),
    .B1(_1392_),
    .Y(_1809_));
 sky130_fd_sc_hd__mux2_1 _4911_ (.A0(_1808_),
    .A1(_1809_),
    .S(_1407_),
    .X(_1810_));
 sky130_fd_sc_hd__a211o_4 _4912_ (.A1(net100),
    .A2(_1341_),
    .B1(_1510_),
    .C1(_1514_),
    .X(_1811_));
 sky130_fd_sc_hd__o21ai_1 _4913_ (.A1(_0822_),
    .A2(_1811_),
    .B1(_1393_),
    .Y(_1812_));
 sky130_fd_sc_hd__o21ai_1 _4914_ (.A1(_0822_),
    .A2(_1522_),
    .B1(_1393_),
    .Y(_1813_));
 sky130_fd_sc_hd__mux2_1 _4915_ (.A0(_1812_),
    .A1(_1813_),
    .S(_1488_),
    .X(_1814_));
 sky130_fd_sc_hd__a211o_4 _4916_ (.A1(net98),
    .A2(_1341_),
    .B1(_1543_),
    .C1(_1546_),
    .X(_1815_));
 sky130_fd_sc_hd__o21ai_1 _4917_ (.A1(_1331_),
    .A2(_1815_),
    .B1(_1393_),
    .Y(_1816_));
 sky130_fd_sc_hd__inv_2 _4918_ (.A(_1553_),
    .Y(_1817_));
 sky130_fd_sc_hd__o21ai_1 _4919_ (.A1(_1331_),
    .A2(_1817_),
    .B1(_1393_),
    .Y(_1818_));
 sky130_fd_sc_hd__mux2_1 _4920_ (.A0(_1816_),
    .A1(_1818_),
    .S(_1488_),
    .X(_1819_));
 sky130_fd_sc_hd__clkinv_2 _4921_ (.A(_1562_),
    .Y(_1820_));
 sky130_fd_sc_hd__o21ai_1 _4922_ (.A1(_1331_),
    .A2(_1820_),
    .B1(_1393_),
    .Y(_1821_));
 sky130_fd_sc_hd__mux2_1 _4923_ (.A0(_1405_),
    .A1(_1821_),
    .S(_1407_),
    .X(_1822_));
 sky130_fd_sc_hd__xnor2_4 _4924_ (.A(_1418_),
    .B(_1423_),
    .Y(_1823_));
 sky130_fd_sc_hd__mux4_1 _4925_ (.A0(_1810_),
    .A1(_1814_),
    .A2(_1819_),
    .A3(_1822_),
    .S0(_1330_),
    .S1(_1823_),
    .X(_1824_));
 sky130_fd_sc_hd__nand2_1 _4926_ (.A(_1421_),
    .B(_1824_),
    .Y(_1825_));
 sky130_fd_sc_hd__clkbuf_4 _4927_ (.A(_1424_),
    .X(_1826_));
 sky130_fd_sc_hd__buf_4 _4928_ (.A(_1488_),
    .X(_1827_));
 sky130_fd_sc_hd__inv_2 _4929_ (.A(_1330_),
    .Y(_1828_));
 sky130_fd_sc_hd__clkbuf_4 _4930_ (.A(_1828_),
    .X(_1829_));
 sky130_fd_sc_hd__and3b_1 _4931_ (.A_N(_1359_),
    .B(_1375_),
    .C(_1733_),
    .X(_1830_));
 sky130_fd_sc_hd__o21ai_1 _4932_ (.A1(_0822_),
    .A2(_1745_),
    .B1(_1393_),
    .Y(_1831_));
 sky130_fd_sc_hd__o21ai_1 _4933_ (.A1(_1331_),
    .A2(_1493_),
    .B1(_1392_),
    .Y(_1832_));
 sky130_fd_sc_hd__mux2_1 _4934_ (.A0(_1831_),
    .A1(_1832_),
    .S(_1827_),
    .X(_1833_));
 sky130_fd_sc_hd__nor2_1 _4935_ (.A(_1829_),
    .B(_1833_),
    .Y(_1834_));
 sky130_fd_sc_hd__a31o_1 _4936_ (.A1(_1827_),
    .A2(_1829_),
    .A3(_1830_),
    .B1(_1834_),
    .X(_1835_));
 sky130_fd_sc_hd__o21ai_1 _4937_ (.A1(_1331_),
    .A2(_1465_),
    .B1(_1392_),
    .Y(_1836_));
 sky130_fd_sc_hd__o21ai_1 _4938_ (.A1(_1331_),
    .A2(_1457_),
    .B1(_1393_),
    .Y(_1837_));
 sky130_fd_sc_hd__mux2_1 _4939_ (.A0(_1836_),
    .A1(_1837_),
    .S(_1407_),
    .X(_1838_));
 sky130_fd_sc_hd__o21ai_1 _4940_ (.A1(_1331_),
    .A2(_1734_),
    .B1(_1392_),
    .Y(_1839_));
 sky130_fd_sc_hd__o21ai_1 _4941_ (.A1(_1331_),
    .A2(_1477_),
    .B1(_1392_),
    .Y(_1840_));
 sky130_fd_sc_hd__mux2_1 _4942_ (.A0(_1839_),
    .A1(_1840_),
    .S(_1407_),
    .X(_1841_));
 sky130_fd_sc_hd__mux2_1 _4943_ (.A0(_1838_),
    .A1(_1841_),
    .S(_1829_),
    .X(_1842_));
 sky130_fd_sc_hd__nor2_1 _4944_ (.A(_1826_),
    .B(_1842_),
    .Y(_1843_));
 sky130_fd_sc_hd__a211o_1 _4945_ (.A1(_1826_),
    .A2(_1835_),
    .B1(_1843_),
    .C1(_1421_),
    .X(_1844_));
 sky130_fd_sc_hd__xnor2_4 _4946_ (.A(_1504_),
    .B(_1420_),
    .Y(_1845_));
 sky130_fd_sc_hd__nor2_1 _4947_ (.A(_1419_),
    .B(_1394_),
    .Y(_1846_));
 sky130_fd_sc_hd__and3b_1 _4948_ (.A_N(_1416_),
    .B(_1845_),
    .C(_1846_),
    .X(_1847_));
 sky130_fd_sc_hd__a31o_1 _4949_ (.A1(_1416_),
    .A2(_1825_),
    .A3(_1844_),
    .B1(_1847_),
    .X(_1848_));
 sky130_fd_sc_hd__nor2_1 _4950_ (.A(_1804_),
    .B(_1733_),
    .Y(_1849_));
 sky130_fd_sc_hd__nor2_1 _4951_ (.A(_1358_),
    .B(_1389_),
    .Y(_1850_));
 sky130_fd_sc_hd__or2_1 _4952_ (.A(_1849_),
    .B(_1850_),
    .X(_1851_));
 sky130_fd_sc_hd__a21oi_1 _4953_ (.A1(_1351_),
    .A2(_1500_),
    .B1(_1851_),
    .Y(_1852_));
 sky130_fd_sc_hd__and2_1 _4954_ (.A(_1351_),
    .B(_1745_),
    .X(_1853_));
 sky130_fd_sc_hd__or2_1 _4955_ (.A(_1351_),
    .B(_1745_),
    .X(_1854_));
 sky130_fd_sc_hd__nor2b_2 _4956_ (.A(_1853_),
    .B_N(_1854_),
    .Y(_1855_));
 sky130_fd_sc_hd__o21a_1 _4957_ (.A1(_1585_),
    .A2(_1493_),
    .B1(_1855_),
    .X(_1856_));
 sky130_fd_sc_hd__inv_2 _4958_ (.A(_1856_),
    .Y(_1857_));
 sky130_fd_sc_hd__or2_1 _4959_ (.A(_1371_),
    .B(_1493_),
    .X(_1858_));
 sky130_fd_sc_hd__nand2_1 _4960_ (.A(_1371_),
    .B(_1493_),
    .Y(_1859_));
 sky130_fd_sc_hd__nand2_1 _4961_ (.A(_1858_),
    .B(_1859_),
    .Y(_1860_));
 sky130_fd_sc_hd__a21o_1 _4962_ (.A1(_1373_),
    .A2(_1478_),
    .B1(_1860_),
    .X(_1861_));
 sky130_fd_sc_hd__nor2_1 _4963_ (.A(_1587_),
    .B(_1478_),
    .Y(_1862_));
 sky130_fd_sc_hd__nor2_1 _4964_ (.A(_1373_),
    .B(_1477_),
    .Y(_1863_));
 sky130_fd_sc_hd__or2_1 _4965_ (.A(_1862_),
    .B(_1863_),
    .X(_1864_));
 sky130_fd_sc_hd__a21o_1 _4966_ (.A1(_1353_),
    .A2(_1484_),
    .B1(_1864_),
    .X(_1865_));
 sky130_fd_sc_hd__xnor2_4 _4967_ (.A(_1362_),
    .B(_1522_),
    .Y(_1866_));
 sky130_fd_sc_hd__nand2_1 _4968_ (.A(_1410_),
    .B(_1547_),
    .Y(_1867_));
 sky130_fd_sc_hd__xnor2_1 _4969_ (.A(_1410_),
    .B(_1547_),
    .Y(_1868_));
 sky130_fd_sc_hd__o221a_1 _4970_ (.A1(_1366_),
    .A2(_1817_),
    .B1(_1866_),
    .B2(_1867_),
    .C1(_1868_),
    .X(_1869_));
 sky130_fd_sc_hd__a21o_1 _4971_ (.A1(_1866_),
    .A2(_1867_),
    .B1(_1869_),
    .X(_1870_));
 sky130_fd_sc_hd__xnor2_1 _4972_ (.A(_1347_),
    .B(_1530_),
    .Y(_1871_));
 sky130_fd_sc_hd__and3_1 _4973_ (.A(_1599_),
    .B(_1515_),
    .C(_1871_),
    .X(_1872_));
 sky130_fd_sc_hd__a21o_1 _4974_ (.A1(_1599_),
    .A2(_1515_),
    .B1(_1871_),
    .X(_1873_));
 sky130_fd_sc_hd__and2b_1 _4975_ (.A_N(_1872_),
    .B(_1873_),
    .X(_1874_));
 sky130_fd_sc_hd__xnor2_2 _4976_ (.A(_1348_),
    .B(_1515_),
    .Y(_1875_));
 sky130_fd_sc_hd__o21ai_1 _4977_ (.A1(_1363_),
    .A2(_1522_),
    .B1(_1875_),
    .Y(_1876_));
 sky130_fd_sc_hd__or3_1 _4978_ (.A(_1363_),
    .B(_1522_),
    .C(_1875_),
    .X(_1877_));
 sky130_fd_sc_hd__and2_1 _4979_ (.A(_1876_),
    .B(_1877_),
    .X(_1878_));
 sky130_fd_sc_hd__o21ai_1 _4980_ (.A1(_1872_),
    .A2(_1876_),
    .B1(_1873_),
    .Y(_1879_));
 sky130_fd_sc_hd__a31o_1 _4981_ (.A1(_1870_),
    .A2(_1874_),
    .A3(_1878_),
    .B1(_1879_),
    .X(_1880_));
 sky130_fd_sc_hd__nand2_1 _4982_ (.A(_1412_),
    .B(_1562_),
    .Y(_1881_));
 sky130_fd_sc_hd__o21bai_2 _4983_ (.A1(_1403_),
    .A2(_1432_),
    .B1_N(_1431_),
    .Y(_1882_));
 sky130_fd_sc_hd__nor2_1 _4984_ (.A(_1413_),
    .B(_1562_),
    .Y(_1883_));
 sky130_fd_sc_hd__nor2_1 _4985_ (.A(_1366_),
    .B(_1553_),
    .Y(_1884_));
 sky130_fd_sc_hd__nand2_1 _4986_ (.A(_1366_),
    .B(_1553_),
    .Y(_1885_));
 sky130_fd_sc_hd__and2b_1 _4987_ (.A_N(_1884_),
    .B(_1885_),
    .X(_1886_));
 sky130_fd_sc_hd__a211o_2 _4988_ (.A1(_1881_),
    .A2(_1882_),
    .B1(_1883_),
    .C1(_1886_),
    .X(_1887_));
 sky130_fd_sc_hd__xor2_1 _4989_ (.A(_1866_),
    .B(_1867_),
    .X(_1888_));
 sky130_fd_sc_hd__and2_1 _4990_ (.A(_1411_),
    .B(_1553_),
    .X(_1889_));
 sky130_fd_sc_hd__xnor2_1 _4991_ (.A(_1868_),
    .B(_1889_),
    .Y(_1890_));
 sky130_fd_sc_hd__and2_1 _4992_ (.A(_1888_),
    .B(_1890_),
    .X(_1891_));
 sky130_fd_sc_hd__and4_1 _4993_ (.A(_1887_),
    .B(_1891_),
    .C(_1874_),
    .D(_1878_),
    .X(_1892_));
 sky130_fd_sc_hd__nor2_2 _4994_ (.A(_1354_),
    .B(_1465_),
    .Y(_1893_));
 sky130_fd_sc_hd__and2_1 _4995_ (.A(_1354_),
    .B(_1465_),
    .X(_1894_));
 sky130_fd_sc_hd__or2_1 _4996_ (.A(_1893_),
    .B(_1894_),
    .X(_1895_));
 sky130_fd_sc_hd__a21o_1 _4997_ (.A1(_1355_),
    .A2(_1537_),
    .B1(_1895_),
    .X(_1896_));
 sky130_fd_sc_hd__and3_1 _4998_ (.A(_1355_),
    .B(_1537_),
    .C(_1895_),
    .X(_1897_));
 sky130_fd_sc_hd__inv_2 _4999_ (.A(_1897_),
    .Y(_1898_));
 sky130_fd_sc_hd__and2_1 _5000_ (.A(_1355_),
    .B(_1746_),
    .X(_1899_));
 sky130_fd_sc_hd__or2_1 _5001_ (.A(_1355_),
    .B(_1746_),
    .X(_1900_));
 sky130_fd_sc_hd__nor2b_2 _5002_ (.A(_1899_),
    .B_N(_1900_),
    .Y(_1901_));
 sky130_fd_sc_hd__o21ai_1 _5003_ (.A1(_1596_),
    .A2(_1531_),
    .B1(_1901_),
    .Y(_1902_));
 sky130_fd_sc_hd__or3_1 _5004_ (.A(_1596_),
    .B(_1530_),
    .C(_1901_),
    .X(_1903_));
 sky130_fd_sc_hd__and2_1 _5005_ (.A(_1902_),
    .B(_1903_),
    .X(_1904_));
 sky130_fd_sc_hd__o2111ai_4 _5006_ (.A1(_1880_),
    .A2(_1892_),
    .B1(_1896_),
    .C1(_1898_),
    .D1(_1904_),
    .Y(_1905_));
 sky130_fd_sc_hd__a21o_1 _5007_ (.A1(_1896_),
    .A2(_1902_),
    .B1(_1897_),
    .X(_1906_));
 sky130_fd_sc_hd__and2_1 _5008_ (.A(_1352_),
    .B(_1456_),
    .X(_1907_));
 sky130_fd_sc_hd__nor2_1 _5009_ (.A(_1352_),
    .B(_1457_),
    .Y(_1908_));
 sky130_fd_sc_hd__or2_2 _5010_ (.A(_1907_),
    .B(_1908_),
    .X(_1909_));
 sky130_fd_sc_hd__and2_1 _5011_ (.A(_1466_),
    .B(_1909_),
    .X(_1910_));
 sky130_fd_sc_hd__a21oi_1 _5012_ (.A1(_1354_),
    .A2(_1466_),
    .B1(_1909_),
    .Y(_1911_));
 sky130_fd_sc_hd__a21o_1 _5013_ (.A1(_1354_),
    .A2(_1910_),
    .B1(_1911_),
    .X(_1912_));
 sky130_fd_sc_hd__nor2_1 _5014_ (.A(_1353_),
    .B(_1734_),
    .Y(_1913_));
 sky130_fd_sc_hd__nor2_1 _5015_ (.A(_1589_),
    .B(_1484_),
    .Y(_1914_));
 sky130_fd_sc_hd__nor2_2 _5016_ (.A(_1913_),
    .B(_1914_),
    .Y(_1915_));
 sky130_fd_sc_hd__o21a_1 _5017_ (.A1(_1591_),
    .A2(_1457_),
    .B1(_1915_),
    .X(_1916_));
 sky130_fd_sc_hd__or3_1 _5018_ (.A(_1591_),
    .B(_1457_),
    .C(_1915_),
    .X(_1917_));
 sky130_fd_sc_hd__and2b_1 _5019_ (.A_N(_1916_),
    .B(_1917_),
    .X(_1918_));
 sky130_fd_sc_hd__inv_2 _5020_ (.A(_1918_),
    .Y(_1919_));
 sky130_fd_sc_hd__a211o_1 _5021_ (.A1(_1905_),
    .A2(_1906_),
    .B1(_1912_),
    .C1(_1919_),
    .X(_1920_));
 sky130_fd_sc_hd__a21o_1 _5022_ (.A1(_1917_),
    .A2(_1911_),
    .B1(_1916_),
    .X(_1921_));
 sky130_fd_sc_hd__inv_2 _5023_ (.A(_1921_),
    .Y(_1922_));
 sky130_fd_sc_hd__nand2_1 _5024_ (.A(_1484_),
    .B(_1864_),
    .Y(_1923_));
 sky130_fd_sc_hd__o21a_1 _5025_ (.A1(_1589_),
    .A2(_1923_),
    .B1(_1865_),
    .X(_1924_));
 sky130_fd_sc_hd__a21bo_2 _5026_ (.A1(_1920_),
    .A2(_1922_),
    .B1_N(_1924_),
    .X(_1925_));
 sky130_fd_sc_hd__and3_1 _5027_ (.A(_1373_),
    .B(_1478_),
    .C(_1860_),
    .X(_1926_));
 sky130_fd_sc_hd__nor2_1 _5028_ (.A(_1493_),
    .B(_1855_),
    .Y(_1927_));
 sky130_fd_sc_hd__a21o_1 _5029_ (.A1(_1371_),
    .A2(_1927_),
    .B1(_1856_),
    .X(_1928_));
 sky130_fd_sc_hd__a311o_1 _5030_ (.A1(_1861_),
    .A2(_1865_),
    .A3(_1925_),
    .B1(_1926_),
    .C1(_1928_),
    .X(_1929_));
 sky130_fd_sc_hd__and3b_1 _5031_ (.A_N(_1852_),
    .B(_1857_),
    .C(_1929_),
    .X(_1930_));
 sky130_fd_sc_hd__nor2_1 _5032_ (.A(_1358_),
    .B(_1733_),
    .Y(_1931_));
 sky130_fd_sc_hd__and3_1 _5033_ (.A(_1351_),
    .B(_1500_),
    .C(_1851_),
    .X(_1932_));
 sky130_fd_sc_hd__o31a_1 _5034_ (.A1(_1930_),
    .A2(_1931_),
    .A3(_1932_),
    .B1(_0862_),
    .X(_1933_));
 sky130_fd_sc_hd__nor2_1 _5035_ (.A(_1585_),
    .B(_1494_),
    .Y(_1934_));
 sky130_fd_sc_hd__nor2_1 _5036_ (.A(_1894_),
    .B(_1899_),
    .Y(_1935_));
 sky130_fd_sc_hd__and2_2 _5037_ (.A(_1347_),
    .B(_1530_),
    .X(_1936_));
 sky130_fd_sc_hd__inv_2 _5038_ (.A(_1866_),
    .Y(_1937_));
 sky130_fd_sc_hd__nor2_1 _5039_ (.A(_1565_),
    .B(_1547_),
    .Y(_1938_));
 sky130_fd_sc_hd__nor2_1 _5040_ (.A(_1410_),
    .B(_1815_),
    .Y(_1939_));
 sky130_fd_sc_hd__or2_2 _5041_ (.A(_1938_),
    .B(_1939_),
    .X(_1940_));
 sky130_fd_sc_hd__nand2_2 _5042_ (.A(_1418_),
    .B(_1562_),
    .Y(_1941_));
 sky130_fd_sc_hd__nor2_1 _5043_ (.A(_1367_),
    .B(_1562_),
    .Y(_1942_));
 sky130_fd_sc_hd__a211o_1 _5044_ (.A1(_1436_),
    .A2(_1441_),
    .B1(_1942_),
    .C1(_1435_),
    .X(_1943_));
 sky130_fd_sc_hd__a31oi_4 _5045_ (.A1(_1885_),
    .A2(_1941_),
    .A3(_1943_),
    .B1(_1884_),
    .Y(_1944_));
 sky130_fd_sc_hd__or2_1 _5046_ (.A(_1347_),
    .B(_1530_),
    .X(_1945_));
 sky130_fd_sc_hd__and2b_1 _5047_ (.A_N(_1936_),
    .B(_1945_),
    .X(_1946_));
 sky130_fd_sc_hd__nand2_1 _5048_ (.A(_1946_),
    .B(_1875_),
    .Y(_1947_));
 sky130_fd_sc_hd__nor4_2 _5049_ (.A(_1937_),
    .B(_1940_),
    .C(_1944_),
    .D(_1947_),
    .Y(_1948_));
 sky130_fd_sc_hd__and2_1 _5050_ (.A(_1599_),
    .B(_1811_),
    .X(_1949_));
 sky130_fd_sc_hd__nand2_1 _5051_ (.A(_1468_),
    .B(_1522_),
    .Y(_1950_));
 sky130_fd_sc_hd__inv_2 _5052_ (.A(_1938_),
    .Y(_1951_));
 sky130_fd_sc_hd__nor2_1 _5053_ (.A(_1468_),
    .B(_1522_),
    .Y(_1952_));
 sky130_fd_sc_hd__a21oi_2 _5054_ (.A1(_1950_),
    .A2(_1951_),
    .B1(_1952_),
    .Y(_1953_));
 sky130_fd_sc_hd__nor2_1 _5055_ (.A(_1599_),
    .B(_1811_),
    .Y(_1954_));
 sky130_fd_sc_hd__inv_2 _5056_ (.A(_1954_),
    .Y(_1955_));
 sky130_fd_sc_hd__o211a_1 _5057_ (.A1(_1949_),
    .A2(_1953_),
    .B1(_1955_),
    .C1(_1945_),
    .X(_1956_));
 sky130_fd_sc_hd__o31ai_4 _5058_ (.A1(_1936_),
    .A2(_1948_),
    .A3(_1956_),
    .B1(_1901_),
    .Y(_1957_));
 sky130_fd_sc_hd__a211oi_4 _5059_ (.A1(_1935_),
    .A2(_1957_),
    .B1(_1893_),
    .C1(_1909_),
    .Y(_1958_));
 sky130_fd_sc_hd__nand2_1 _5060_ (.A(_1589_),
    .B(_1484_),
    .Y(_1959_));
 sky130_fd_sc_hd__inv_2 _5061_ (.A(_1864_),
    .Y(_1960_));
 sky130_fd_sc_hd__o311a_1 _5062_ (.A1(_1914_),
    .A2(_1907_),
    .A3(_1958_),
    .B1(_1959_),
    .C1(_1960_),
    .X(_1961_));
 sky130_fd_sc_hd__o31a_1 _5063_ (.A1(_1934_),
    .A2(_1862_),
    .A3(_1961_),
    .B1(_1858_),
    .X(_1962_));
 sky130_fd_sc_hd__and2_1 _5064_ (.A(_1855_),
    .B(_1962_),
    .X(_1963_));
 sky130_fd_sc_hd__nand2_1 _5065_ (.A(_1358_),
    .B(_1389_),
    .Y(_1964_));
 sky130_fd_sc_hd__o311a_1 _5066_ (.A1(_1850_),
    .A2(_1853_),
    .A3(_1963_),
    .B1(_1964_),
    .C1(_0780_),
    .X(_1965_));
 sky130_fd_sc_hd__a211o_4 _5067_ (.A1(_1807_),
    .A2(_1848_),
    .B1(_1933_),
    .C1(_1965_),
    .X(_1966_));
 sky130_fd_sc_hd__nor2_1 _5068_ (.A(_1804_),
    .B(_1966_),
    .Y(_1967_));
 sky130_fd_sc_hd__xnor2_1 _5069_ (.A(_1803_),
    .B(_1967_),
    .Y(_1968_));
 sky130_fd_sc_hd__mux2_1 _5070_ (.A0(\core_1.ew_addr_high[0] ),
    .A1(_1968_),
    .S(_1801_),
    .X(_1969_));
 sky130_fd_sc_hd__clkbuf_1 _5071_ (.A(_1969_),
    .X(_0220_));
 sky130_fd_sc_hd__and2_1 _5072_ (.A(\core_1.execute.rf.reg_outputs[1][1] ),
    .B(_1459_),
    .X(_1970_));
 sky130_fd_sc_hd__or3_1 _5073_ (.A(_1396_),
    .B(_1397_),
    .C(_1398_),
    .X(_1971_));
 sky130_fd_sc_hd__or3_1 _5074_ (.A(_1970_),
    .B(_1971_),
    .C(_1803_),
    .X(_1972_));
 sky130_fd_sc_hd__inv_2 _5075_ (.A(_1972_),
    .Y(_1973_));
 sky130_fd_sc_hd__o21a_1 _5076_ (.A1(_1970_),
    .A2(_1971_),
    .B1(_1803_),
    .X(_1974_));
 sky130_fd_sc_hd__or2_2 _5077_ (.A(_1973_),
    .B(_1974_),
    .X(_1975_));
 sky130_fd_sc_hd__o21ba_1 _5078_ (.A1(_1804_),
    .A2(_1803_),
    .B1_N(_1966_),
    .X(_1976_));
 sky130_fd_sc_hd__xnor2_4 _5079_ (.A(_1975_),
    .B(_1976_),
    .Y(_1977_));
 sky130_fd_sc_hd__mux2_1 _5080_ (.A0(net132),
    .A1(_1977_),
    .S(_1801_),
    .X(_1978_));
 sky130_fd_sc_hd__clkbuf_1 _5081_ (.A(_1978_),
    .X(_0221_));
 sky130_fd_sc_hd__nor2_2 _5082_ (.A(_1358_),
    .B(_1966_),
    .Y(_1979_));
 sky130_fd_sc_hd__o22a_1 _5083_ (.A1(_1966_),
    .A2(_1973_),
    .B1(_1974_),
    .B2(_1979_),
    .X(_1980_));
 sky130_fd_sc_hd__a221o_2 _5084_ (.A1(\core_1.execute.rf.reg_outputs[1][2] ),
    .A2(_1459_),
    .B1(_1472_),
    .B2(\core_1.execute.rf.reg_outputs[3][2] ),
    .C1(_1557_),
    .X(_1981_));
 sky130_fd_sc_hd__xor2_4 _5085_ (.A(_1980_),
    .B(_1981_),
    .X(_1982_));
 sky130_fd_sc_hd__mux2_1 _5086_ (.A0(net133),
    .A1(_1982_),
    .S(_1801_),
    .X(_1983_));
 sky130_fd_sc_hd__clkbuf_1 _5087_ (.A(_1983_),
    .X(_0222_));
 sky130_fd_sc_hd__nor2_1 _5088_ (.A(_1972_),
    .B(_1981_),
    .Y(_1984_));
 sky130_fd_sc_hd__and2_1 _5089_ (.A(_1979_),
    .B(_1984_),
    .X(_1985_));
 sky130_fd_sc_hd__and3_1 _5090_ (.A(_1966_),
    .B(_1974_),
    .C(_1981_),
    .X(_1986_));
 sky130_fd_sc_hd__or2_2 _5091_ (.A(_1985_),
    .B(_1986_),
    .X(_1987_));
 sky130_fd_sc_hd__a21oi_4 _5092_ (.A1(\core_1.execute.rf.reg_outputs[1][3] ),
    .A2(_1459_),
    .B1(_1549_),
    .Y(_1988_));
 sky130_fd_sc_hd__xnor2_4 _5093_ (.A(_1987_),
    .B(_1988_),
    .Y(_1989_));
 sky130_fd_sc_hd__mux2_1 _5094_ (.A0(net134),
    .A1(_1989_),
    .S(_1801_),
    .X(_1990_));
 sky130_fd_sc_hd__clkbuf_1 _5095_ (.A(_1990_),
    .X(_0223_));
 sky130_fd_sc_hd__a21o_1 _5096_ (.A1(\core_1.execute.rf.reg_outputs[1][4] ),
    .A2(_1459_),
    .B1(_1545_),
    .X(_1991_));
 sky130_fd_sc_hd__a21o_1 _5097_ (.A1(\core_1.execute.rf.reg_outputs[1][3] ),
    .A2(_1459_),
    .B1(_1549_),
    .X(_1992_));
 sky130_fd_sc_hd__nand2_1 _5098_ (.A(_1986_),
    .B(_1992_),
    .Y(_1993_));
 sky130_fd_sc_hd__a21bo_1 _5099_ (.A1(_1985_),
    .A2(_1988_),
    .B1_N(_1993_),
    .X(_1994_));
 sky130_fd_sc_hd__a21oi_1 _5100_ (.A1(_1991_),
    .A2(_1994_),
    .B1(_1796_),
    .Y(_1995_));
 sky130_fd_sc_hd__o21a_1 _5101_ (.A1(_1991_),
    .A2(_1994_),
    .B1(_1995_),
    .X(_1996_));
 sky130_fd_sc_hd__a21o_1 _5102_ (.A1(net135),
    .A2(_1796_),
    .B1(_1996_),
    .X(_0224_));
 sky130_fd_sc_hd__a21o_1 _5103_ (.A1(\core_1.execute.rf.reg_outputs[1][5] ),
    .A2(_1459_),
    .B1(_1517_),
    .X(_1997_));
 sky130_fd_sc_hd__a31oi_1 _5104_ (.A1(_1979_),
    .A2(_1984_),
    .A3(_1988_),
    .B1(_1991_),
    .Y(_1998_));
 sky130_fd_sc_hd__a21oi_1 _5105_ (.A1(_1993_),
    .A2(_1991_),
    .B1(_1998_),
    .Y(_1999_));
 sky130_fd_sc_hd__xor2_1 _5106_ (.A(_1997_),
    .B(_1999_),
    .X(_2000_));
 sky130_fd_sc_hd__mux2_1 _5107_ (.A0(net136),
    .A1(_2000_),
    .S(_1801_),
    .X(_2001_));
 sky130_fd_sc_hd__clkbuf_1 _5108_ (.A(_2001_),
    .X(_0225_));
 sky130_fd_sc_hd__a21o_1 _5109_ (.A1(\core_1.execute.rf.reg_outputs[1][6] ),
    .A2(_1459_),
    .B1(_1513_),
    .X(_2002_));
 sky130_fd_sc_hd__xor2_1 _5110_ (.A(_1979_),
    .B(_1997_),
    .X(_2003_));
 sky130_fd_sc_hd__nand2_1 _5111_ (.A(_1999_),
    .B(_2003_),
    .Y(_2004_));
 sky130_fd_sc_hd__xnor2_1 _5112_ (.A(_2002_),
    .B(_2004_),
    .Y(_2005_));
 sky130_fd_sc_hd__mux2_1 _5113_ (.A0(net137),
    .A1(_2005_),
    .S(_1801_),
    .X(_2006_));
 sky130_fd_sc_hd__clkbuf_1 _5114_ (.A(_2006_),
    .X(_0226_));
 sky130_fd_sc_hd__a21oi_1 _5115_ (.A1(\core_1.execute.rf.reg_outputs[1][7] ),
    .A2(_1459_),
    .B1(_1528_),
    .Y(_2007_));
 sky130_fd_sc_hd__xnor2_1 _5116_ (.A(_1979_),
    .B(_2002_),
    .Y(_2008_));
 sky130_fd_sc_hd__nor2_1 _5117_ (.A(_2004_),
    .B(_2008_),
    .Y(_2009_));
 sky130_fd_sc_hd__xnor2_1 _5118_ (.A(_2007_),
    .B(_2009_),
    .Y(_2010_));
 sky130_fd_sc_hd__mux2_1 _5119_ (.A0(net138),
    .A1(_2010_),
    .S(_1801_),
    .X(_2011_));
 sky130_fd_sc_hd__clkbuf_1 _5120_ (.A(_2011_),
    .X(_0227_));
 sky130_fd_sc_hd__and3b_1 _5121_ (.A_N(net187),
    .B(net186),
    .C(_1011_),
    .X(_2012_));
 sky130_fd_sc_hd__and3_2 _5122_ (.A(_1009_),
    .B(_1016_),
    .C(_2012_),
    .X(_2013_));
 sky130_fd_sc_hd__nand2_1 _5123_ (.A(net187),
    .B(_1011_),
    .Y(_2014_));
 sky130_fd_sc_hd__and4bb_2 _5124_ (.A_N(_1009_),
    .B_N(_2014_),
    .C(_1010_),
    .D(_1016_),
    .X(_2015_));
 sky130_fd_sc_hd__and4b_2 _5125_ (.A_N(net192),
    .B(_1013_),
    .C(_1014_),
    .D(net185),
    .X(_2016_));
 sky130_fd_sc_hd__and3_1 _5126_ (.A(net211),
    .B(_1012_),
    .C(_2016_),
    .X(_2017_));
 sky130_fd_sc_hd__buf_2 _5127_ (.A(_2017_),
    .X(_2018_));
 sky130_fd_sc_hd__a22o_1 _5128_ (.A1(net72),
    .A2(_1017_),
    .B1(_2018_),
    .B2(\core_1.execute.sreg_irq_pc.o_d[0] ),
    .X(_2019_));
 sky130_fd_sc_hd__a221o_1 _5129_ (.A1(\core_1.execute.alu_flag_reg.o_d[0] ),
    .A2(_2013_),
    .B1(_2015_),
    .B2(net1),
    .C1(_2019_),
    .X(_2020_));
 sky130_fd_sc_hd__and3_2 _5130_ (.A(_1009_),
    .B(_2016_),
    .C(_2012_),
    .X(_2021_));
 sky130_fd_sc_hd__and3_1 _5131_ (.A(net187),
    .B(net186),
    .C(_1011_),
    .X(_2022_));
 sky130_fd_sc_hd__and3_1 _5132_ (.A(_1008_),
    .B(_1015_),
    .C(_2022_),
    .X(_2023_));
 sky130_fd_sc_hd__clkbuf_4 _5133_ (.A(_2023_),
    .X(_2024_));
 sky130_fd_sc_hd__a22o_1 _5134_ (.A1(\core_1.execute.sreg_scratch.o_d[0] ),
    .A2(_2021_),
    .B1(_2024_),
    .B2(\core_1.execute.pc_high_out[0] ),
    .X(_2025_));
 sky130_fd_sc_hd__and3_1 _5135_ (.A(net211),
    .B(_1015_),
    .C(_2012_),
    .X(_2026_));
 sky130_fd_sc_hd__and3_2 _5136_ (.A(_1009_),
    .B(_1012_),
    .C(_2016_),
    .X(_2027_));
 sky130_fd_sc_hd__a22o_1 _5137_ (.A1(\core_1.execute.sreg_irq_flags.o_d[0] ),
    .A2(_2026_),
    .B1(_2027_),
    .B2(net106),
    .X(_2028_));
 sky130_fd_sc_hd__nor2_1 _5138_ (.A(net186),
    .B(_2014_),
    .Y(_2029_));
 sky130_fd_sc_hd__and3_2 _5139_ (.A(net211),
    .B(_2016_),
    .C(_2012_),
    .X(_2030_));
 sky130_fd_sc_hd__a311o_1 _5140_ (.A1(_1009_),
    .A2(_1016_),
    .A3(_2029_),
    .B1(_2030_),
    .C1(\core_1.dec_sreg_jal_over ),
    .X(_2031_));
 sky130_fd_sc_hd__and3_2 _5141_ (.A(net211),
    .B(_1016_),
    .C(_2022_),
    .X(_2032_));
 sky130_fd_sc_hd__a22o_1 _5142_ (.A1(\core_1.execute.sreg_priv_control.o_d[0] ),
    .A2(_1144_),
    .B1(_2032_),
    .B2(\core_1.execute.pc_high_buff_out[0] ),
    .X(_2033_));
 sky130_fd_sc_hd__or4_1 _5143_ (.A(_2025_),
    .B(_2028_),
    .C(_2031_),
    .D(_2033_),
    .X(_2034_));
 sky130_fd_sc_hd__o22a_1 _5144_ (.A1(net72),
    .A2(_1137_),
    .B1(_2020_),
    .B2(_2034_),
    .X(_2035_));
 sky130_fd_sc_hd__or2_1 _5145_ (.A(\core_1.execute.sreg_irq_pc.o_d[0] ),
    .B(_1140_),
    .X(_2036_));
 sky130_fd_sc_hd__o21ai_1 _5146_ (.A1(_1146_),
    .A2(_2035_),
    .B1(_2036_),
    .Y(_2037_));
 sky130_fd_sc_hd__xnor2_1 _5147_ (.A(\core_1.dec_sreg_jal_over ),
    .B(_2037_),
    .Y(_2038_));
 sky130_fd_sc_hd__o211a_2 _5148_ (.A1(_0822_),
    .A2(\core_1.decode.oc_alu_mode[13] ),
    .B1(_1363_),
    .C1(_1416_),
    .X(_2039_));
 sky130_fd_sc_hd__and2b_1 _5149_ (.A_N(_1440_),
    .B(_1439_),
    .X(_2040_));
 sky130_fd_sc_hd__nand2_2 _5150_ (.A(_1343_),
    .B(_1345_),
    .Y(_2041_));
 sky130_fd_sc_hd__nor2_2 _5151_ (.A(\core_1.decode.oc_alu_mode[3] ),
    .B(_1445_),
    .Y(_2042_));
 sky130_fd_sc_hd__nor2_1 _5152_ (.A(_2041_),
    .B(_2042_),
    .Y(_2043_));
 sky130_fd_sc_hd__a221o_1 _5153_ (.A1(_0846_),
    .A2(_1827_),
    .B1(_1439_),
    .B2(\core_1.decode.oc_alu_mode[9] ),
    .C1(_2043_),
    .X(_2044_));
 sky130_fd_sc_hd__and2_1 _5154_ (.A(_1438_),
    .B(_2040_),
    .X(_2045_));
 sky130_fd_sc_hd__inv_2 _5155_ (.A(\core_1.decode.oc_alu_mode[4] ),
    .Y(_2046_));
 sky130_fd_sc_hd__clkinv_2 _5156_ (.A(\core_1.decode.oc_alu_mode[11] ),
    .Y(_2047_));
 sky130_fd_sc_hd__a2bb2o_1 _5157_ (.A1_N(_1438_),
    .A2_N(_2040_),
    .B1(_2046_),
    .B2(_2047_),
    .X(_2048_));
 sky130_fd_sc_hd__a2bb2o_1 _5158_ (.A1_N(_2045_),
    .A2_N(_2048_),
    .B1(\core_1.decode.oc_alu_mode[2] ),
    .B2(_1440_),
    .X(_2049_));
 sky130_fd_sc_hd__a211o_1 _5159_ (.A1(_0832_),
    .A2(_2040_),
    .B1(_2044_),
    .C1(_2049_),
    .X(_2050_));
 sky130_fd_sc_hd__a31o_1 _5160_ (.A1(_2039_),
    .A2(_1845_),
    .A3(_1846_),
    .B1(_2050_),
    .X(_2051_));
 sky130_fd_sc_hd__mux2_1 _5161_ (.A0(_1466_),
    .A1(_1537_),
    .S(_1406_),
    .X(_2052_));
 sky130_fd_sc_hd__mux2_1 _5162_ (.A0(_1458_),
    .A1(_1484_),
    .S(_1328_),
    .X(_2053_));
 sky130_fd_sc_hd__o22a_1 _5163_ (.A1(_1470_),
    .A2(_2052_),
    .B1(_2053_),
    .B2(_1486_),
    .X(_2054_));
 sky130_fd_sc_hd__mux2_1 _5164_ (.A0(_1478_),
    .A1(_1494_),
    .S(_1488_),
    .X(_2055_));
 sky130_fd_sc_hd__mux2_1 _5165_ (.A0(_1389_),
    .A1(_1500_),
    .S(_1406_),
    .X(_2056_));
 sky130_fd_sc_hd__o22a_1 _5166_ (.A1(_1470_),
    .A2(_2055_),
    .B1(_2056_),
    .B2(_1486_),
    .X(_2057_));
 sky130_fd_sc_hd__mux2_1 _5167_ (.A0(_2054_),
    .A1(_2057_),
    .S(_1505_),
    .X(_2058_));
 sky130_fd_sc_hd__mux2_1 _5168_ (.A0(_1523_),
    .A1(_1547_),
    .S(_1406_),
    .X(_2059_));
 sky130_fd_sc_hd__mux2_1 _5169_ (.A0(_1811_),
    .A1(_1531_),
    .S(_1328_),
    .X(_2060_));
 sky130_fd_sc_hd__inv_2 _5170_ (.A(_2060_),
    .Y(_2061_));
 sky130_fd_sc_hd__o22a_1 _5171_ (.A1(_1470_),
    .A2(_2059_),
    .B1(_2061_),
    .B2(_1486_),
    .X(_2062_));
 sky130_fd_sc_hd__mux2_2 _5172_ (.A0(_1817_),
    .A1(_1820_),
    .S(_1407_),
    .X(_2063_));
 sky130_fd_sc_hd__nand2_1 _5173_ (.A(_1555_),
    .B(_1407_),
    .Y(_2064_));
 sky130_fd_sc_hd__nor2_1 _5174_ (.A(_1827_),
    .B(_2041_),
    .Y(_2065_));
 sky130_fd_sc_hd__a21o_1 _5175_ (.A1(_2064_),
    .A2(_1436_),
    .B1(_2065_),
    .X(_2066_));
 sky130_fd_sc_hd__o21ai_1 _5176_ (.A1(_1555_),
    .A2(_2063_),
    .B1(_2066_),
    .Y(_2067_));
 sky130_fd_sc_hd__a21o_1 _5177_ (.A1(_1414_),
    .A2(_2067_),
    .B1(_1566_),
    .X(_2068_));
 sky130_fd_sc_hd__a31o_1 _5178_ (.A1(_1504_),
    .A2(_1507_),
    .A3(_2062_),
    .B1(_2068_),
    .X(_2069_));
 sky130_fd_sc_hd__a21oi_1 _5179_ (.A1(_1451_),
    .A2(_2058_),
    .B1(_2069_),
    .Y(_2070_));
 sky130_fd_sc_hd__or2_2 _5180_ (.A(_2051_),
    .B(_2070_),
    .X(_2071_));
 sky130_fd_sc_hd__or2_1 _5181_ (.A(\core_1.execute.alu_mul_div.i_mul ),
    .B(_2071_),
    .X(_2072_));
 sky130_fd_sc_hd__inv_2 _5182_ (.A(\core_1.execute.alu_mul_div.mul_res[0] ),
    .Y(_2073_));
 sky130_fd_sc_hd__a21oi_1 _5183_ (.A1(_0859_),
    .A2(_2073_),
    .B1(\core_1.execute.alu_mul_div.i_div ),
    .Y(_2074_));
 sky130_fd_sc_hd__a221o_1 _5184_ (.A1(\core_1.execute.alu_mul_div.div_res[0] ),
    .A2(\core_1.execute.alu_mul_div.i_div ),
    .B1(_2072_),
    .B2(_2074_),
    .C1(\core_1.execute.alu_mul_div.i_mod ),
    .X(_2075_));
 sky130_fd_sc_hd__o21a_4 _5185_ (.A1(_1313_),
    .A2(\core_1.execute.alu_mul_div.div_cur[0] ),
    .B1(_2075_),
    .X(_2076_));
 sky130_fd_sc_hd__nor2_4 _5186_ (.A(\core_1.dec_sreg_load ),
    .B(\core_1.dec_sreg_jal_over ),
    .Y(_2077_));
 sky130_fd_sc_hd__buf_6 _5187_ (.A(_2077_),
    .X(_2078_));
 sky130_fd_sc_hd__mux2_1 _5188_ (.A0(_2038_),
    .A1(_2076_),
    .S(_2078_),
    .X(_2079_));
 sky130_fd_sc_hd__clkinv_2 _5189_ (.A(\core_1.dec_mem_access ),
    .Y(_2080_));
 sky130_fd_sc_hd__buf_4 _5190_ (.A(_2080_),
    .X(_2081_));
 sky130_fd_sc_hd__mux2_1 _5191_ (.A0(net194),
    .A1(_2079_),
    .S(_2081_),
    .X(_2082_));
 sky130_fd_sc_hd__mux2_1 _5192_ (.A0(\core_1.ew_data[0] ),
    .A1(_2082_),
    .S(_1801_),
    .X(_2083_));
 sky130_fd_sc_hd__clkbuf_1 _5193_ (.A(_2083_),
    .X(_0229_));
 sky130_fd_sc_hd__buf_4 _5194_ (.A(_2077_),
    .X(_2084_));
 sky130_fd_sc_hd__nor2_1 _5195_ (.A(net79),
    .B(_1137_),
    .Y(_2085_));
 sky130_fd_sc_hd__a22o_1 _5196_ (.A1(net79),
    .A2(_1017_),
    .B1(_2027_),
    .B2(\core_1.execute.trap_flag ),
    .X(_2086_));
 sky130_fd_sc_hd__and4_1 _5197_ (.A(\core_1.execute.pc_high_buff_out[1] ),
    .B(net211),
    .C(_1016_),
    .D(_2022_),
    .X(_2087_));
 sky130_fd_sc_hd__and4_1 _5198_ (.A(\core_1.execute.sreg_irq_flags.o_d[1] ),
    .B(net211),
    .C(_1016_),
    .D(_2012_),
    .X(_2088_));
 sky130_fd_sc_hd__and4_1 _5199_ (.A(\core_1.execute.sreg_scratch.o_d[1] ),
    .B(_1009_),
    .C(_2016_),
    .D(_2012_),
    .X(_2089_));
 sky130_fd_sc_hd__a2111o_1 _5200_ (.A1(net8),
    .A2(_2015_),
    .B1(_2087_),
    .C1(_2088_),
    .D1(_2089_),
    .X(_2090_));
 sky130_fd_sc_hd__and4_1 _5201_ (.A(\core_1.execute.alu_flag_reg.o_d[1] ),
    .B(_1009_),
    .C(_1016_),
    .D(_2012_),
    .X(_2091_));
 sky130_fd_sc_hd__and4_1 _5202_ (.A(\core_1.execute.pc_high_out[1] ),
    .B(_1009_),
    .C(_1016_),
    .D(_2022_),
    .X(_2092_));
 sky130_fd_sc_hd__a2111o_1 _5203_ (.A1(\core_1.execute.sreg_data_page ),
    .A2(_1144_),
    .B1(_2091_),
    .C1(_2092_),
    .D1(\core_1.dec_sreg_jal_over ),
    .X(_2093_));
 sky130_fd_sc_hd__a2111oi_2 _5204_ (.A1(\core_1.execute.sreg_irq_pc.o_d[1] ),
    .A2(_2018_),
    .B1(_2086_),
    .C1(_2090_),
    .D1(_2093_),
    .Y(_2094_));
 sky130_fd_sc_hd__o31ai_1 _5205_ (.A1(\core_1.dec_sreg_irt ),
    .A2(_2085_),
    .A3(_2094_),
    .B1(_1310_),
    .Y(_2095_));
 sky130_fd_sc_hd__o2111a_1 _5206_ (.A1(_1018_),
    .A2(_2035_),
    .B1(_2036_),
    .C1(_2095_),
    .D1(\core_1.dec_sreg_jal_over ),
    .X(_2096_));
 sky130_fd_sc_hd__o21ba_1 _5207_ (.A1(_1138_),
    .A2(_2037_),
    .B1_N(_2095_),
    .X(_2097_));
 sky130_fd_sc_hd__nand2_1 _5208_ (.A(_1573_),
    .B(_2084_),
    .Y(_2098_));
 sky130_fd_sc_hd__o31ai_1 _5209_ (.A1(_2084_),
    .A2(_2096_),
    .A3(_2097_),
    .B1(_2098_),
    .Y(_2099_));
 sky130_fd_sc_hd__mux2_1 _5210_ (.A0(net201),
    .A1(_2099_),
    .S(_2081_),
    .X(_2100_));
 sky130_fd_sc_hd__clkbuf_8 _5211_ (.A(_1800_),
    .X(_2101_));
 sky130_fd_sc_hd__mux2_1 _5212_ (.A0(\core_1.ew_data[1] ),
    .A1(_2100_),
    .S(_2101_),
    .X(_2102_));
 sky130_fd_sc_hd__clkbuf_1 _5213_ (.A(_2102_),
    .X(_0230_));
 sky130_fd_sc_hd__a21bo_1 _5214_ (.A1(\core_1.execute.alu_mul_div.div_res[2] ),
    .A2(_1313_),
    .B1_N(_1314_),
    .X(_2103_));
 sky130_fd_sc_hd__buf_2 _5215_ (.A(\core_1.execute.alu_mul_div.i_mul ),
    .X(_2104_));
 sky130_fd_sc_hd__mux2_1 _5216_ (.A0(_1405_),
    .A1(_1821_),
    .S(_1407_),
    .X(_2105_));
 sky130_fd_sc_hd__o32a_1 _5217_ (.A1(_1555_),
    .A2(_1827_),
    .A3(_1394_),
    .B1(_2105_),
    .B2(_1330_),
    .X(_2106_));
 sky130_fd_sc_hd__or3_1 _5218_ (.A(_1319_),
    .B(_1506_),
    .C(_2056_),
    .X(_2107_));
 sky130_fd_sc_hd__or3_1 _5219_ (.A(_1319_),
    .B(_1506_),
    .C(_2053_),
    .X(_2108_));
 sky130_fd_sc_hd__o311a_1 _5220_ (.A1(_1555_),
    .A2(_1506_),
    .A3(_2055_),
    .B1(_2108_),
    .C1(_1418_),
    .X(_2109_));
 sky130_fd_sc_hd__a21oi_2 _5221_ (.A1(_1505_),
    .A2(_2107_),
    .B1(_2109_),
    .Y(_2110_));
 sky130_fd_sc_hd__mux2_1 _5222_ (.A0(_2052_),
    .A1(_2061_),
    .S(_1555_),
    .X(_2111_));
 sky130_fd_sc_hd__nor2_1 _5223_ (.A(_1506_),
    .B(_2111_),
    .Y(_2112_));
 sky130_fd_sc_hd__a21oi_1 _5224_ (.A1(_1319_),
    .A2(_2059_),
    .B1(_1506_),
    .Y(_2113_));
 sky130_fd_sc_hd__o211a_1 _5225_ (.A1(_1319_),
    .A2(_2063_),
    .B1(_2113_),
    .C1(_1418_),
    .X(_2114_));
 sky130_fd_sc_hd__a211o_1 _5226_ (.A1(_1505_),
    .A2(_2112_),
    .B1(_2114_),
    .C1(_1451_),
    .X(_2115_));
 sky130_fd_sc_hd__inv_2 _5227_ (.A(_1566_),
    .Y(_2116_));
 sky130_fd_sc_hd__o211ai_4 _5228_ (.A1(_1504_),
    .A2(_2110_),
    .B1(_2115_),
    .C1(_2116_),
    .Y(_2117_));
 sky130_fd_sc_hd__inv_2 _5229_ (.A(_1882_),
    .Y(_2118_));
 sky130_fd_sc_hd__a21o_1 _5230_ (.A1(_1436_),
    .A2(_1441_),
    .B1(_1435_),
    .X(_2119_));
 sky130_fd_sc_hd__or2_1 _5231_ (.A(_1413_),
    .B(_1562_),
    .X(_2120_));
 sky130_fd_sc_hd__nand2_1 _5232_ (.A(_1881_),
    .B(_2120_),
    .Y(_2121_));
 sky130_fd_sc_hd__a221o_1 _5233_ (.A1(_0862_),
    .A2(_2118_),
    .B1(_2119_),
    .B2(\core_1.decode.oc_alu_mode[4] ),
    .C1(_2121_),
    .X(_2122_));
 sky130_fd_sc_hd__a2bb2o_1 _5234_ (.A1_N(_2046_),
    .A2_N(_2119_),
    .B1(_1882_),
    .B2(_0862_),
    .X(_2123_));
 sky130_fd_sc_hd__or3b_1 _5235_ (.A(\core_1.decode.oc_alu_mode[6] ),
    .B(_2123_),
    .C_N(_2121_),
    .X(_2124_));
 sky130_fd_sc_hd__a22o_1 _5236_ (.A1(\core_1.decode.oc_alu_mode[7] ),
    .A2(_1413_),
    .B1(_1446_),
    .B2(_1820_),
    .X(_2125_));
 sky130_fd_sc_hd__a221o_1 _5237_ (.A1(_0814_),
    .A2(_1941_),
    .B1(_1942_),
    .B2(\core_1.decode.oc_alu_mode[2] ),
    .C1(_2125_),
    .X(_2126_));
 sky130_fd_sc_hd__a21oi_1 _5238_ (.A1(_2122_),
    .A2(_2124_),
    .B1(_2126_),
    .Y(_2127_));
 sky130_fd_sc_hd__o211a_1 _5239_ (.A1(_1425_),
    .A2(_2106_),
    .B1(_2117_),
    .C1(_2127_),
    .X(_2128_));
 sky130_fd_sc_hd__nor2_1 _5240_ (.A(_2104_),
    .B(_2128_),
    .Y(_2129_));
 sky130_fd_sc_hd__a211o_1 _5241_ (.A1(_0860_),
    .A2(\core_1.execute.alu_mul_div.mul_res[2] ),
    .B1(_2129_),
    .C1(_0831_),
    .X(_2130_));
 sky130_fd_sc_hd__a22o_2 _5242_ (.A1(\core_1.execute.alu_mul_div.div_cur[2] ),
    .A2(_0835_),
    .B1(_2103_),
    .B2(_2130_),
    .X(_2131_));
 sky130_fd_sc_hd__or2_1 _5243_ (.A(\core_1.dec_sreg_jal_over ),
    .B(_1017_),
    .X(_2132_));
 sky130_fd_sc_hd__a22o_1 _5244_ (.A1(\core_1.execute.alu_flag_reg.o_d[2] ),
    .A2(_2013_),
    .B1(_2027_),
    .B2(net105),
    .X(_2133_));
 sky130_fd_sc_hd__a22o_1 _5245_ (.A1(\core_1.execute.irq_en ),
    .A2(_1144_),
    .B1(_2015_),
    .B2(net9),
    .X(_2134_));
 sky130_fd_sc_hd__a22o_1 _5246_ (.A1(\core_1.execute.sreg_irq_flags.o_d[2] ),
    .A2(_2026_),
    .B1(_2032_),
    .B2(\core_1.execute.pc_high_buff_out[2] ),
    .X(_2135_));
 sky130_fd_sc_hd__a2111o_1 _5247_ (.A1(\core_1.execute.pc_high_out[2] ),
    .A2(_2024_),
    .B1(_2133_),
    .C1(_2134_),
    .D1(_2135_),
    .X(_2136_));
 sky130_fd_sc_hd__a221o_1 _5248_ (.A1(\core_1.execute.sreg_irq_pc.o_d[2] ),
    .A2(_2018_),
    .B1(_2021_),
    .B2(\core_1.execute.sreg_scratch.o_d[2] ),
    .C1(_2136_),
    .X(_2137_));
 sky130_fd_sc_hd__a22o_1 _5249_ (.A1(net80),
    .A2(_2132_),
    .B1(_2137_),
    .B2(_1137_),
    .X(_2138_));
 sky130_fd_sc_hd__or2_1 _5250_ (.A(\core_1.execute.sreg_irq_pc.o_d[2] ),
    .B(_1140_),
    .X(_2139_));
 sky130_fd_sc_hd__o21a_1 _5251_ (.A1(_1146_),
    .A2(_2138_),
    .B1(_2139_),
    .X(_2140_));
 sky130_fd_sc_hd__or2_1 _5252_ (.A(_2096_),
    .B(_2140_),
    .X(_2141_));
 sky130_fd_sc_hd__o211a_1 _5253_ (.A1(_1018_),
    .A2(_2138_),
    .B1(_2139_),
    .C1(_2096_),
    .X(_2142_));
 sky130_fd_sc_hd__nor2_1 _5254_ (.A(_2077_),
    .B(_2142_),
    .Y(_2143_));
 sky130_fd_sc_hd__a22o_1 _5255_ (.A1(_2084_),
    .A2(_2131_),
    .B1(_2141_),
    .B2(_2143_),
    .X(_2144_));
 sky130_fd_sc_hd__mux2_1 _5256_ (.A0(net202),
    .A1(_2144_),
    .S(_2081_),
    .X(_2145_));
 sky130_fd_sc_hd__mux2_1 _5257_ (.A0(\core_1.ew_data[2] ),
    .A1(_2145_),
    .S(_2101_),
    .X(_2146_));
 sky130_fd_sc_hd__clkbuf_1 _5258_ (.A(_2146_),
    .X(_0231_));
 sky130_fd_sc_hd__a22o_1 _5259_ (.A1(\core_1.execute.sreg_long_ptr_en ),
    .A2(_1144_),
    .B1(_2013_),
    .B2(\core_1.execute.alu_flag_reg.o_d[3] ),
    .X(_2147_));
 sky130_fd_sc_hd__a221o_1 _5260_ (.A1(\core_1.execute.sreg_irq_pc.o_d[3] ),
    .A2(_2018_),
    .B1(_2026_),
    .B2(\core_1.execute.sreg_irq_flags.o_d[3] ),
    .C1(_2147_),
    .X(_2148_));
 sky130_fd_sc_hd__a22o_1 _5261_ (.A1(net10),
    .A2(_2015_),
    .B1(_2032_),
    .B2(\core_1.execute.pc_high_buff_out[3] ),
    .X(_2149_));
 sky130_fd_sc_hd__a221o_1 _5262_ (.A1(\core_1.execute.sreg_scratch.o_d[3] ),
    .A2(_2021_),
    .B1(_2024_),
    .B2(\core_1.execute.pc_high_out[3] ),
    .C1(_2149_),
    .X(_2150_));
 sky130_fd_sc_hd__nor2_1 _5263_ (.A(_2148_),
    .B(_2150_),
    .Y(_2151_));
 sky130_fd_sc_hd__o2bb2a_1 _5264_ (.A1_N(net81),
    .A2_N(_2132_),
    .B1(_2151_),
    .B2(\core_1.dec_sreg_jal_over ),
    .X(_2152_));
 sky130_fd_sc_hd__nand2_1 _5265_ (.A(\core_1.execute.sreg_irq_pc.o_d[3] ),
    .B(_1018_),
    .Y(_2153_));
 sky130_fd_sc_hd__o21a_1 _5266_ (.A1(_1018_),
    .A2(_2152_),
    .B1(_2153_),
    .X(_2154_));
 sky130_fd_sc_hd__xnor2_1 _5267_ (.A(_2142_),
    .B(_2154_),
    .Y(_2155_));
 sky130_fd_sc_hd__a21bo_1 _5268_ (.A1(\core_1.execute.alu_mul_div.div_res[3] ),
    .A2(_1313_),
    .B1_N(_1314_),
    .X(_2156_));
 sky130_fd_sc_hd__mux2_1 _5269_ (.A0(_1818_),
    .A1(_1821_),
    .S(_1488_),
    .X(_2157_));
 sky130_fd_sc_hd__mux2_1 _5270_ (.A0(_1408_),
    .A1(_2157_),
    .S(_1829_),
    .X(_2158_));
 sky130_fd_sc_hd__or2_1 _5271_ (.A(_1425_),
    .B(_2158_),
    .X(_2159_));
 sky130_fd_sc_hd__or2_1 _5272_ (.A(_1389_),
    .B(_1506_),
    .X(_2160_));
 sky130_fd_sc_hd__or3_1 _5273_ (.A(_2064_),
    .B(_1418_),
    .C(_2160_),
    .X(_2161_));
 sky130_fd_sc_hd__mux2_1 _5274_ (.A0(_1485_),
    .A1(_1501_),
    .S(_1319_),
    .X(_2162_));
 sky130_fd_sc_hd__or3_1 _5275_ (.A(_1413_),
    .B(_1506_),
    .C(_2162_),
    .X(_2163_));
 sky130_fd_sc_hd__mux2_1 _5276_ (.A0(_1524_),
    .A1(_1554_),
    .S(_1555_),
    .X(_2164_));
 sky130_fd_sc_hd__mux2_1 _5277_ (.A0(_1467_),
    .A1(_1539_),
    .S(_1555_),
    .X(_2165_));
 sky130_fd_sc_hd__nor2_1 _5278_ (.A(_1506_),
    .B(_2165_),
    .Y(_2166_));
 sky130_fd_sc_hd__nand2_1 _5279_ (.A(_1413_),
    .B(_2166_),
    .Y(_2167_));
 sky130_fd_sc_hd__o311a_1 _5280_ (.A1(_1413_),
    .A2(_1506_),
    .A3(_2164_),
    .B1(_2167_),
    .C1(_1504_),
    .X(_2168_));
 sky130_fd_sc_hd__a31o_1 _5281_ (.A1(_1451_),
    .A2(_2161_),
    .A3(_2163_),
    .B1(_2168_),
    .X(_2169_));
 sky130_fd_sc_hd__a21o_1 _5282_ (.A1(_1881_),
    .A2(_1882_),
    .B1(_1883_),
    .X(_2170_));
 sky130_fd_sc_hd__nand2_1 _5283_ (.A(_1941_),
    .B(_1943_),
    .Y(_2171_));
 sky130_fd_sc_hd__o22a_1 _5284_ (.A1(_2047_),
    .A2(_2170_),
    .B1(_2171_),
    .B2(_2046_),
    .X(_2172_));
 sky130_fd_sc_hd__a221o_1 _5285_ (.A1(_0862_),
    .A2(_2170_),
    .B1(_2171_),
    .B2(\core_1.decode.oc_alu_mode[4] ),
    .C1(\core_1.decode.oc_alu_mode[6] ),
    .X(_2173_));
 sky130_fd_sc_hd__a221o_1 _5286_ (.A1(\core_1.decode.oc_alu_mode[7] ),
    .A2(_1451_),
    .B1(_1884_),
    .B2(\core_1.decode.oc_alu_mode[2] ),
    .C1(\core_1.decode.oc_alu_mode[9] ),
    .X(_2174_));
 sky130_fd_sc_hd__a22oi_1 _5287_ (.A1(_1886_),
    .A2(_2173_),
    .B1(_2174_),
    .B2(_1885_),
    .Y(_2175_));
 sky130_fd_sc_hd__o221a_1 _5288_ (.A1(_1566_),
    .A2(_2169_),
    .B1(_2172_),
    .B2(_1886_),
    .C1(_2175_),
    .X(_2176_));
 sky130_fd_sc_hd__o211a_1 _5289_ (.A1(_2042_),
    .A2(_1553_),
    .B1(_2159_),
    .C1(_2176_),
    .X(_2177_));
 sky130_fd_sc_hd__nor2_1 _5290_ (.A(_2104_),
    .B(_2177_),
    .Y(_2178_));
 sky130_fd_sc_hd__a211o_1 _5291_ (.A1(_2104_),
    .A2(\core_1.execute.alu_mul_div.mul_res[3] ),
    .B1(_2178_),
    .C1(_0831_),
    .X(_2179_));
 sky130_fd_sc_hd__a22o_2 _5292_ (.A1(\core_1.execute.alu_mul_div.div_cur[3] ),
    .A2(_0835_),
    .B1(_2156_),
    .B2(_2179_),
    .X(_2180_));
 sky130_fd_sc_hd__mux2_1 _5293_ (.A0(_2155_),
    .A1(_2180_),
    .S(_2078_),
    .X(_2181_));
 sky130_fd_sc_hd__mux2_1 _5294_ (.A0(net203),
    .A1(_2181_),
    .S(_2081_),
    .X(_2182_));
 sky130_fd_sc_hd__mux2_1 _5295_ (.A0(\core_1.ew_data[3] ),
    .A1(_2182_),
    .S(_2101_),
    .X(_2183_));
 sky130_fd_sc_hd__clkbuf_1 _5296_ (.A(_2183_),
    .X(_0232_));
 sky130_fd_sc_hd__a221o_1 _5297_ (.A1(\core_1.execute.sreg_irq_pc.o_d[4] ),
    .A2(_2018_),
    .B1(_2032_),
    .B2(\core_1.execute.pc_high_buff_out[4] ),
    .C1(_2030_),
    .X(_2184_));
 sky130_fd_sc_hd__a22o_1 _5298_ (.A1(net11),
    .A2(_2015_),
    .B1(_2021_),
    .B2(\core_1.execute.sreg_scratch.o_d[4] ),
    .X(_2185_));
 sky130_fd_sc_hd__a22o_1 _5299_ (.A1(\core_1.execute.sreg_priv_control.o_d[4] ),
    .A2(_1144_),
    .B1(_2026_),
    .B2(\core_1.execute.sreg_irq_flags.o_d[4] ),
    .X(_2186_));
 sky130_fd_sc_hd__a21o_1 _5300_ (.A1(\core_1.execute.pc_high_out[4] ),
    .A2(_2024_),
    .B1(_2186_),
    .X(_2187_));
 sky130_fd_sc_hd__a2111o_1 _5301_ (.A1(\core_1.execute.alu_flag_reg.o_d[4] ),
    .A2(_2013_),
    .B1(_2184_),
    .C1(_2185_),
    .D1(_2187_),
    .X(_2188_));
 sky130_fd_sc_hd__a22o_1 _5302_ (.A1(net82),
    .A2(_2132_),
    .B1(_2188_),
    .B2(_1137_),
    .X(_2189_));
 sky130_fd_sc_hd__nand2_1 _5303_ (.A(\core_1.execute.sreg_irq_pc.o_d[4] ),
    .B(_1018_),
    .Y(_2190_));
 sky130_fd_sc_hd__a21boi_1 _5304_ (.A1(_1140_),
    .A2(_2189_),
    .B1_N(_2190_),
    .Y(_2191_));
 sky130_fd_sc_hd__nor3b_1 _5305_ (.A(_2154_),
    .B(_2191_),
    .C_N(_2142_),
    .Y(_2192_));
 sky130_fd_sc_hd__or2b_1 _5306_ (.A(_2154_),
    .B_N(_2142_),
    .X(_2193_));
 sky130_fd_sc_hd__a21o_1 _5307_ (.A1(_2193_),
    .A2(_2191_),
    .B1(_2077_),
    .X(_2194_));
 sky130_fd_sc_hd__a21bo_1 _5308_ (.A1(\core_1.execute.alu_mul_div.div_res[4] ),
    .A2(_1313_),
    .B1_N(_1314_),
    .X(_2195_));
 sky130_fd_sc_hd__mux2_1 _5309_ (.A0(_1816_),
    .A1(_1818_),
    .S(_1488_),
    .X(_2196_));
 sky130_fd_sc_hd__mux2_1 _5310_ (.A0(_2105_),
    .A1(_2196_),
    .S(_1829_),
    .X(_2197_));
 sky130_fd_sc_hd__or3_1 _5311_ (.A(_2064_),
    .B(_1418_),
    .C(_1394_),
    .X(_2198_));
 sky130_fd_sc_hd__o21ai_2 _5312_ (.A1(_1823_),
    .A2(_2197_),
    .B1(_2198_),
    .Y(_2199_));
 sky130_fd_sc_hd__nor2_1 _5313_ (.A(_1940_),
    .B(_1944_),
    .Y(_2200_));
 sky130_fd_sc_hd__a21o_1 _5314_ (.A1(_1940_),
    .A2(_1944_),
    .B1(_2046_),
    .X(_2201_));
 sky130_fd_sc_hd__nor2_1 _5315_ (.A(_2200_),
    .B(_2201_),
    .Y(_2202_));
 sky130_fd_sc_hd__a221o_1 _5316_ (.A1(\core_1.decode.oc_alu_mode[7] ),
    .A2(_1410_),
    .B1(_1446_),
    .B2(_1815_),
    .C1(\core_1.decode.oc_alu_mode[9] ),
    .X(_2203_));
 sky130_fd_sc_hd__and2b_1 _5317_ (.A_N(_1939_),
    .B(_2203_),
    .X(_2204_));
 sky130_fd_sc_hd__a221o_1 _5318_ (.A1(_0839_),
    .A2(_1938_),
    .B1(_1868_),
    .B2(_0832_),
    .C1(_2204_),
    .X(_2205_));
 sky130_fd_sc_hd__nor2_1 _5319_ (.A(_1505_),
    .B(_2057_),
    .Y(_2206_));
 sky130_fd_sc_hd__nor2_1 _5320_ (.A(_1451_),
    .B(_1418_),
    .Y(_2207_));
 sky130_fd_sc_hd__a221o_1 _5321_ (.A1(_1414_),
    .A2(_2062_),
    .B1(_2207_),
    .B2(_2054_),
    .C1(_1566_),
    .X(_2208_));
 sky130_fd_sc_hd__o21ba_1 _5322_ (.A1(_1504_),
    .A2(_2206_),
    .B1_N(_2208_),
    .X(_2209_));
 sky130_fd_sc_hd__or3_1 _5323_ (.A(_2202_),
    .B(_2205_),
    .C(_2209_),
    .X(_2210_));
 sky130_fd_sc_hd__nand2_1 _5324_ (.A(_1887_),
    .B(_1890_),
    .Y(_2211_));
 sky130_fd_sc_hd__o211a_1 _5325_ (.A1(_1940_),
    .A2(_1887_),
    .B1(_2211_),
    .C1(_0863_),
    .X(_2212_));
 sky130_fd_sc_hd__a211oi_4 _5326_ (.A1(_1422_),
    .A2(_2199_),
    .B1(_2210_),
    .C1(_2212_),
    .Y(_2213_));
 sky130_fd_sc_hd__nor2_1 _5327_ (.A(_2104_),
    .B(_2213_),
    .Y(_2214_));
 sky130_fd_sc_hd__a211o_1 _5328_ (.A1(_0860_),
    .A2(\core_1.execute.alu_mul_div.mul_res[4] ),
    .B1(_2214_),
    .C1(_0831_),
    .X(_2215_));
 sky130_fd_sc_hd__a22o_2 _5329_ (.A1(\core_1.execute.alu_mul_div.div_cur[4] ),
    .A2(_0835_),
    .B1(_2195_),
    .B2(_2215_),
    .X(_2216_));
 sky130_fd_sc_hd__a2bb2o_1 _5330_ (.A1_N(_2192_),
    .A2_N(_2194_),
    .B1(_2084_),
    .B2(_2216_),
    .X(_2217_));
 sky130_fd_sc_hd__mux2_1 _5331_ (.A0(net204),
    .A1(_2217_),
    .S(_2081_),
    .X(_2218_));
 sky130_fd_sc_hd__mux2_1 _5332_ (.A0(\core_1.ew_data[4] ),
    .A1(_2218_),
    .S(_2101_),
    .X(_2219_));
 sky130_fd_sc_hd__clkbuf_1 _5333_ (.A(_2219_),
    .X(_0233_));
 sky130_fd_sc_hd__a22o_1 _5334_ (.A1(\core_1.execute.sreg_irq_pc.o_d[5] ),
    .A2(_2018_),
    .B1(_2024_),
    .B2(\core_1.execute.pc_high_out[5] ),
    .X(_2220_));
 sky130_fd_sc_hd__a221o_1 _5335_ (.A1(net12),
    .A2(_2015_),
    .B1(_2021_),
    .B2(\core_1.execute.sreg_scratch.o_d[5] ),
    .C1(_2220_),
    .X(_2221_));
 sky130_fd_sc_hd__a221o_1 _5336_ (.A1(\core_1.execute.sreg_priv_control.o_d[5] ),
    .A2(_1144_),
    .B1(_2032_),
    .B2(\core_1.execute.pc_high_buff_out[5] ),
    .C1(_2221_),
    .X(_2222_));
 sky130_fd_sc_hd__a22o_1 _5337_ (.A1(net83),
    .A2(_2132_),
    .B1(_2222_),
    .B2(_1137_),
    .X(_2223_));
 sky130_fd_sc_hd__nand2_1 _5338_ (.A(\core_1.execute.sreg_irq_pc.o_d[5] ),
    .B(_1018_),
    .Y(_2224_));
 sky130_fd_sc_hd__a21bo_1 _5339_ (.A1(_1140_),
    .A2(_2223_),
    .B1_N(_2224_),
    .X(_2225_));
 sky130_fd_sc_hd__nor2_1 _5340_ (.A(_2192_),
    .B(_2225_),
    .Y(_2226_));
 sky130_fd_sc_hd__nand2_2 _5341_ (.A(_2192_),
    .B(_2225_),
    .Y(_2227_));
 sky130_fd_sc_hd__and2b_1 _5342_ (.A_N(_2226_),
    .B(_2227_),
    .X(_2228_));
 sky130_fd_sc_hd__a21bo_1 _5343_ (.A1(\core_1.execute.alu_mul_div.div_res[5] ),
    .A2(_1313_),
    .B1_N(_0727_),
    .X(_2229_));
 sky130_fd_sc_hd__nand2_1 _5344_ (.A(_2039_),
    .B(_1845_),
    .Y(_2230_));
 sky130_fd_sc_hd__mux2_1 _5345_ (.A0(_1813_),
    .A1(_1816_),
    .S(_1488_),
    .X(_2231_));
 sky130_fd_sc_hd__mux2_1 _5346_ (.A0(_2157_),
    .A1(_2231_),
    .S(_1828_),
    .X(_2232_));
 sky130_fd_sc_hd__mux2_1 _5347_ (.A0(_1409_),
    .A1(_2232_),
    .S(_1424_),
    .X(_2233_));
 sky130_fd_sc_hd__o21a_1 _5348_ (.A1(_1938_),
    .A2(_2200_),
    .B1(_1866_),
    .X(_2234_));
 sky130_fd_sc_hd__o211a_1 _5349_ (.A1(_1940_),
    .A2(_1944_),
    .B1(_1937_),
    .C1(_1951_),
    .X(_2235_));
 sky130_fd_sc_hd__nor2_1 _5350_ (.A(_1886_),
    .B(_2170_),
    .Y(_2236_));
 sky130_fd_sc_hd__o21a_1 _5351_ (.A1(_1889_),
    .A2(_2236_),
    .B1(_1940_),
    .X(_2237_));
 sky130_fd_sc_hd__xnor2_1 _5352_ (.A(_1888_),
    .B(_2237_),
    .Y(_2238_));
 sky130_fd_sc_hd__nand2_1 _5353_ (.A(_0863_),
    .B(_2238_),
    .Y(_2239_));
 sky130_fd_sc_hd__a21oi_1 _5354_ (.A1(_0832_),
    .A2(_1950_),
    .B1(_0814_),
    .Y(_2240_));
 sky130_fd_sc_hd__a21oi_1 _5355_ (.A1(_0839_),
    .A2(_1522_),
    .B1(_0846_),
    .Y(_2241_));
 sky130_fd_sc_hd__o22a_1 _5356_ (.A1(_2042_),
    .A2(_1523_),
    .B1(_2241_),
    .B2(_1363_),
    .X(_2242_));
 sky130_fd_sc_hd__nor2_1 _5357_ (.A(_1505_),
    .B(_1502_),
    .Y(_2243_));
 sky130_fd_sc_hd__a21oi_1 _5358_ (.A1(_1505_),
    .A2(_1487_),
    .B1(_1451_),
    .Y(_2244_));
 sky130_fd_sc_hd__a21oi_1 _5359_ (.A1(_1414_),
    .A2(_1540_),
    .B1(_1566_),
    .Y(_2245_));
 sky130_fd_sc_hd__o21ai_1 _5360_ (.A1(_2243_),
    .A2(_2244_),
    .B1(_2245_),
    .Y(_2246_));
 sky130_fd_sc_hd__o211a_1 _5361_ (.A1(_1952_),
    .A2(_2240_),
    .B1(_2242_),
    .C1(_2246_),
    .X(_2247_));
 sky130_fd_sc_hd__o311a_1 _5362_ (.A1(_2046_),
    .A2(_2234_),
    .A3(_2235_),
    .B1(_2239_),
    .C1(_2247_),
    .X(_2248_));
 sky130_fd_sc_hd__o21ai_4 _5363_ (.A1(_2230_),
    .A2(_2233_),
    .B1(_2248_),
    .Y(_2249_));
 sky130_fd_sc_hd__a21o_1 _5364_ (.A1(_0859_),
    .A2(\core_1.execute.alu_mul_div.mul_res[5] ),
    .B1(\core_1.execute.alu_mul_div.i_div ),
    .X(_2250_));
 sky130_fd_sc_hd__a21o_1 _5365_ (.A1(_1316_),
    .A2(_2249_),
    .B1(_2250_),
    .X(_2251_));
 sky130_fd_sc_hd__a22o_2 _5366_ (.A1(\core_1.execute.alu_mul_div.div_cur[5] ),
    .A2(_0835_),
    .B1(_2229_),
    .B2(_2251_),
    .X(_2252_));
 sky130_fd_sc_hd__mux2_1 _5367_ (.A0(_2228_),
    .A1(_2252_),
    .S(_2078_),
    .X(_2253_));
 sky130_fd_sc_hd__mux2_1 _5368_ (.A0(net205),
    .A1(_2253_),
    .S(_2081_),
    .X(_2254_));
 sky130_fd_sc_hd__mux2_1 _5369_ (.A0(\core_1.ew_data[5] ),
    .A1(_2254_),
    .S(_2101_),
    .X(_2255_));
 sky130_fd_sc_hd__clkbuf_1 _5370_ (.A(_2255_),
    .X(_0234_));
 sky130_fd_sc_hd__clkbuf_4 _5371_ (.A(_2132_),
    .X(_2256_));
 sky130_fd_sc_hd__buf_4 _5372_ (.A(_2015_),
    .X(_2257_));
 sky130_fd_sc_hd__a22o_1 _5373_ (.A1(\core_1.execute.sreg_irq_pc.o_d[6] ),
    .A2(_2018_),
    .B1(_2024_),
    .B2(\core_1.execute.pc_high_out[6] ),
    .X(_2258_));
 sky130_fd_sc_hd__a221o_1 _5374_ (.A1(\core_1.execute.sreg_priv_control.o_d[6] ),
    .A2(_1144_),
    .B1(_2021_),
    .B2(\core_1.execute.sreg_scratch.o_d[6] ),
    .C1(_2258_),
    .X(_2259_));
 sky130_fd_sc_hd__a221o_1 _5375_ (.A1(net13),
    .A2(_2257_),
    .B1(_2032_),
    .B2(\core_1.execute.pc_high_buff_out[6] ),
    .C1(_2259_),
    .X(_2260_));
 sky130_fd_sc_hd__a22o_1 _5376_ (.A1(net84),
    .A2(_2256_),
    .B1(_2260_),
    .B2(_1137_),
    .X(_2261_));
 sky130_fd_sc_hd__nand2_1 _5377_ (.A(\core_1.execute.sreg_irq_pc.o_d[6] ),
    .B(_1018_),
    .Y(_2262_));
 sky130_fd_sc_hd__a21bo_2 _5378_ (.A1(_1140_),
    .A2(_2261_),
    .B1_N(_2262_),
    .X(_2263_));
 sky130_fd_sc_hd__xnor2_1 _5379_ (.A(_2227_),
    .B(_2263_),
    .Y(_2264_));
 sky130_fd_sc_hd__a21bo_1 _5380_ (.A1(\core_1.execute.alu_mul_div.div_res[6] ),
    .A2(_1312_),
    .B1_N(_0727_),
    .X(_2265_));
 sky130_fd_sc_hd__o32a_1 _5381_ (.A1(_1555_),
    .A2(_1827_),
    .A3(_1394_),
    .B1(_1822_),
    .B2(_1330_),
    .X(_2266_));
 sky130_fd_sc_hd__mux2_1 _5382_ (.A0(_1814_),
    .A1(_1819_),
    .S(_1330_),
    .X(_2267_));
 sky130_fd_sc_hd__mux2_1 _5383_ (.A0(_2266_),
    .A1(_2267_),
    .S(_1826_),
    .X(_2268_));
 sky130_fd_sc_hd__nand2_1 _5384_ (.A(_1504_),
    .B(_1418_),
    .Y(_2269_));
 sky130_fd_sc_hd__o22a_1 _5385_ (.A1(_1470_),
    .A2(_2053_),
    .B1(_2055_),
    .B2(_1486_),
    .X(_2270_));
 sky130_fd_sc_hd__a2bb2o_1 _5386_ (.A1_N(_2269_),
    .A2_N(_2112_),
    .B1(_2207_),
    .B2(_2270_),
    .X(_2271_));
 sky130_fd_sc_hd__o21a_1 _5387_ (.A1(_1505_),
    .A2(_2107_),
    .B1(_1451_),
    .X(_2272_));
 sky130_fd_sc_hd__inv_2 _5388_ (.A(\core_1.decode.oc_alu_mode[6] ),
    .Y(_2273_));
 sky130_fd_sc_hd__a21oi_1 _5389_ (.A1(_0839_),
    .A2(_1599_),
    .B1(_1446_),
    .Y(_2274_));
 sky130_fd_sc_hd__a21oi_1 _5390_ (.A1(_0846_),
    .A2(_1599_),
    .B1(_0814_),
    .Y(_2275_));
 sky130_fd_sc_hd__o221a_1 _5391_ (.A1(_2273_),
    .A2(_1949_),
    .B1(_2274_),
    .B2(_1515_),
    .C1(_2275_),
    .X(_2276_));
 sky130_fd_sc_hd__o32a_1 _5392_ (.A1(_1566_),
    .A2(_2271_),
    .A3(_2272_),
    .B1(_1954_),
    .B2(_2276_),
    .X(_2277_));
 sky130_fd_sc_hd__and2_1 _5393_ (.A(_1866_),
    .B(_2200_),
    .X(_2278_));
 sky130_fd_sc_hd__o21ai_1 _5394_ (.A1(_2278_),
    .A2(_1953_),
    .B1(_1875_),
    .Y(_2279_));
 sky130_fd_sc_hd__or3_1 _5395_ (.A(_1875_),
    .B(_2278_),
    .C(_1953_),
    .X(_2280_));
 sky130_fd_sc_hd__a21o_1 _5396_ (.A1(_1887_),
    .A2(_1891_),
    .B1(_1870_),
    .X(_2281_));
 sky130_fd_sc_hd__xor2_1 _5397_ (.A(_2281_),
    .B(_1878_),
    .X(_2282_));
 sky130_fd_sc_hd__a32o_1 _5398_ (.A1(_0780_),
    .A2(_2279_),
    .A3(_2280_),
    .B1(_0862_),
    .B2(_2282_),
    .X(_2283_));
 sky130_fd_sc_hd__inv_2 _5399_ (.A(_2283_),
    .Y(_2284_));
 sky130_fd_sc_hd__o211a_2 _5400_ (.A1(_2230_),
    .A2(_2268_),
    .B1(_2277_),
    .C1(_2284_),
    .X(_2285_));
 sky130_fd_sc_hd__nor2_1 _5401_ (.A(_0859_),
    .B(_2285_),
    .Y(_2286_));
 sky130_fd_sc_hd__a211o_1 _5402_ (.A1(_2104_),
    .A2(\core_1.execute.alu_mul_div.mul_res[6] ),
    .B1(_2286_),
    .C1(_0831_),
    .X(_2287_));
 sky130_fd_sc_hd__a22o_2 _5403_ (.A1(\core_1.execute.alu_mul_div.div_cur[6] ),
    .A2(\core_1.execute.alu_mul_div.i_mod ),
    .B1(_2265_),
    .B2(_2287_),
    .X(_2288_));
 sky130_fd_sc_hd__mux2_1 _5404_ (.A0(_2264_),
    .A1(_2288_),
    .S(_2078_),
    .X(_2289_));
 sky130_fd_sc_hd__mux2_1 _5405_ (.A0(net206),
    .A1(_2289_),
    .S(_2081_),
    .X(_2290_));
 sky130_fd_sc_hd__mux2_1 _5406_ (.A0(\core_1.ew_data[6] ),
    .A1(_2290_),
    .S(_2101_),
    .X(_2291_));
 sky130_fd_sc_hd__clkbuf_1 _5407_ (.A(_2291_),
    .X(_0235_));
 sky130_fd_sc_hd__or2b_1 _5408_ (.A(_2227_),
    .B_N(_2263_),
    .X(_2292_));
 sky130_fd_sc_hd__buf_4 _5409_ (.A(_2021_),
    .X(_2293_));
 sky130_fd_sc_hd__buf_4 _5410_ (.A(_2018_),
    .X(_2294_));
 sky130_fd_sc_hd__a22o_1 _5411_ (.A1(\core_1.execute.sreg_irq_pc.o_d[7] ),
    .A2(_2294_),
    .B1(_2024_),
    .B2(\core_1.execute.pc_high_out[7] ),
    .X(_2295_));
 sky130_fd_sc_hd__a221o_1 _5412_ (.A1(\core_1.execute.sreg_priv_control.o_d[7] ),
    .A2(_1145_),
    .B1(_2293_),
    .B2(\core_1.execute.sreg_scratch.o_d[7] ),
    .C1(_2295_),
    .X(_2296_));
 sky130_fd_sc_hd__a221o_1 _5413_ (.A1(net14),
    .A2(_2257_),
    .B1(_2032_),
    .B2(\core_1.execute.pc_high_buff_out[7] ),
    .C1(_2296_),
    .X(_2297_));
 sky130_fd_sc_hd__a22o_1 _5414_ (.A1(net85),
    .A2(_2256_),
    .B1(_2297_),
    .B2(_1138_),
    .X(_2298_));
 sky130_fd_sc_hd__nand2_1 _5415_ (.A(\core_1.execute.sreg_irq_pc.o_d[7] ),
    .B(_1018_),
    .Y(_2299_));
 sky130_fd_sc_hd__a21bo_2 _5416_ (.A1(_1140_),
    .A2(_2298_),
    .B1_N(_2299_),
    .X(_2300_));
 sky130_fd_sc_hd__xnor2_1 _5417_ (.A(_2292_),
    .B(_2300_),
    .Y(_2301_));
 sky130_fd_sc_hd__a21bo_1 _5418_ (.A1(\core_1.execute.alu_mul_div.div_res[7] ),
    .A2(_1312_),
    .B1_N(_0727_),
    .X(_2302_));
 sky130_fd_sc_hd__or3b_1 _5419_ (.A(_1946_),
    .B(_1949_),
    .C_N(_2279_),
    .X(_2303_));
 sky130_fd_sc_hd__nand2_1 _5420_ (.A(_1599_),
    .B(_1811_),
    .Y(_2304_));
 sky130_fd_sc_hd__a21o_1 _5421_ (.A1(_2304_),
    .A2(_2279_),
    .B1(_1871_),
    .X(_2305_));
 sky130_fd_sc_hd__a21bo_1 _5422_ (.A1(_2281_),
    .A2(_1878_),
    .B1_N(_1876_),
    .X(_2306_));
 sky130_fd_sc_hd__xor2_1 _5423_ (.A(_1874_),
    .B(_2306_),
    .X(_2307_));
 sky130_fd_sc_hd__mux2_1 _5424_ (.A0(_1808_),
    .A1(_1812_),
    .S(_1488_),
    .X(_2308_));
 sky130_fd_sc_hd__mux2_1 _5425_ (.A0(_2231_),
    .A1(_2308_),
    .S(_1829_),
    .X(_2309_));
 sky130_fd_sc_hd__mux2_1 _5426_ (.A0(_2158_),
    .A1(_2309_),
    .S(_1826_),
    .X(_2310_));
 sky130_fd_sc_hd__nor2_1 _5427_ (.A(_2230_),
    .B(_2310_),
    .Y(_2311_));
 sky130_fd_sc_hd__nor2_2 _5428_ (.A(_1419_),
    .B(_2160_),
    .Y(_2312_));
 sky130_fd_sc_hd__o22a_1 _5429_ (.A1(_1470_),
    .A2(_1485_),
    .B1(_1486_),
    .B2(_1501_),
    .X(_2313_));
 sky130_fd_sc_hd__nand2_1 _5430_ (.A(_2207_),
    .B(_2313_),
    .Y(_2314_));
 sky130_fd_sc_hd__o221a_1 _5431_ (.A1(_2269_),
    .A2(_2166_),
    .B1(_2312_),
    .B2(_1504_),
    .C1(_2314_),
    .X(_2315_));
 sky130_fd_sc_hd__a22o_1 _5432_ (.A1(_0846_),
    .A2(_1347_),
    .B1(_1446_),
    .B2(_1531_),
    .X(_2316_));
 sky130_fd_sc_hd__a221o_1 _5433_ (.A1(_0814_),
    .A2(_1945_),
    .B1(_1946_),
    .B2(_0832_),
    .C1(_2316_),
    .X(_2317_));
 sky130_fd_sc_hd__a221o_1 _5434_ (.A1(_0839_),
    .A2(_1936_),
    .B1(_2315_),
    .B2(_2116_),
    .C1(_2317_),
    .X(_2318_));
 sky130_fd_sc_hd__a211o_1 _5435_ (.A1(_0863_),
    .A2(_2307_),
    .B1(_2311_),
    .C1(_2318_),
    .X(_2319_));
 sky130_fd_sc_hd__a31o_2 _5436_ (.A1(_0780_),
    .A2(_2303_),
    .A3(_2305_),
    .B1(_2319_),
    .X(_2320_));
 sky130_fd_sc_hd__a21o_1 _5437_ (.A1(_0859_),
    .A2(\core_1.execute.alu_mul_div.mul_res[7] ),
    .B1(\core_1.execute.alu_mul_div.i_div ),
    .X(_2321_));
 sky130_fd_sc_hd__a21o_1 _5438_ (.A1(_1316_),
    .A2(_2320_),
    .B1(_2321_),
    .X(_2322_));
 sky130_fd_sc_hd__a22o_2 _5439_ (.A1(\core_1.execute.alu_mul_div.div_cur[7] ),
    .A2(\core_1.execute.alu_mul_div.i_mod ),
    .B1(_2302_),
    .B2(_2322_),
    .X(_2323_));
 sky130_fd_sc_hd__mux2_1 _5440_ (.A0(_2301_),
    .A1(_2323_),
    .S(_2078_),
    .X(_2324_));
 sky130_fd_sc_hd__mux2_1 _5441_ (.A0(net207),
    .A1(_2324_),
    .S(_2081_),
    .X(_2325_));
 sky130_fd_sc_hd__mux2_1 _5442_ (.A0(\core_1.ew_data[7] ),
    .A1(_2325_),
    .S(_2101_),
    .X(_2326_));
 sky130_fd_sc_hd__clkbuf_1 _5443_ (.A(_2326_),
    .X(_0236_));
 sky130_fd_sc_hd__or2b_1 _5444_ (.A(_2292_),
    .B_N(_2300_),
    .X(_2327_));
 sky130_fd_sc_hd__a22o_1 _5445_ (.A1(net15),
    .A2(_2257_),
    .B1(_2293_),
    .B2(\core_1.execute.sreg_scratch.o_d[8] ),
    .X(_2328_));
 sky130_fd_sc_hd__a221o_1 _5446_ (.A1(\core_1.execute.sreg_priv_control.o_d[8] ),
    .A2(_1145_),
    .B1(_2294_),
    .B2(\core_1.execute.sreg_irq_pc.o_d[8] ),
    .C1(_2328_),
    .X(_2329_));
 sky130_fd_sc_hd__a22oi_1 _5447_ (.A1(net86),
    .A2(_2256_),
    .B1(_2329_),
    .B2(_1138_),
    .Y(_2330_));
 sky130_fd_sc_hd__nand2_1 _5448_ (.A(\core_1.execute.sreg_irq_pc.o_d[8] ),
    .B(_1018_),
    .Y(_2331_));
 sky130_fd_sc_hd__o21ai_2 _5449_ (.A1(_1019_),
    .A2(_2330_),
    .B1(_2331_),
    .Y(_2332_));
 sky130_fd_sc_hd__xnor2_1 _5450_ (.A(_2327_),
    .B(_2332_),
    .Y(_2333_));
 sky130_fd_sc_hd__a21bo_1 _5451_ (.A1(\core_1.execute.alu_mul_div.div_res[8] ),
    .A2(_1312_),
    .B1_N(_0727_),
    .X(_2334_));
 sky130_fd_sc_hd__or2_1 _5452_ (.A(_1880_),
    .B(_1892_),
    .X(_2335_));
 sky130_fd_sc_hd__nand2_1 _5453_ (.A(_1904_),
    .B(_2335_),
    .Y(_2336_));
 sky130_fd_sc_hd__and2_1 _5454_ (.A(_0862_),
    .B(_2336_),
    .X(_2337_));
 sky130_fd_sc_hd__o21a_1 _5455_ (.A1(_1904_),
    .A2(_2335_),
    .B1(_2337_),
    .X(_2338_));
 sky130_fd_sc_hd__inv_2 _5456_ (.A(_2058_),
    .Y(_2339_));
 sky130_fd_sc_hd__nor2_4 _5457_ (.A(_1451_),
    .B(_1566_),
    .Y(_2340_));
 sky130_fd_sc_hd__and2_4 _5458_ (.A(\core_1.decode.oc_alu_mode[3] ),
    .B(_1531_),
    .X(_2341_));
 sky130_fd_sc_hd__a221o_1 _5459_ (.A1(_0846_),
    .A2(_1355_),
    .B1(_1900_),
    .B2(\core_1.decode.oc_alu_mode[9] ),
    .C1(_2341_),
    .X(_2342_));
 sky130_fd_sc_hd__a22o_1 _5460_ (.A1(_1445_),
    .A2(_1746_),
    .B1(_1899_),
    .B2(\core_1.decode.oc_alu_mode[2] ),
    .X(_2343_));
 sky130_fd_sc_hd__a211o_1 _5461_ (.A1(_0832_),
    .A2(_1901_),
    .B1(_2342_),
    .C1(_2343_),
    .X(_2344_));
 sky130_fd_sc_hd__and2_1 _5462_ (.A(\core_1.decode.oc_alu_mode[4] ),
    .B(_1957_),
    .X(_2345_));
 sky130_fd_sc_hd__o41a_1 _5463_ (.A1(_1901_),
    .A2(_1936_),
    .A3(_1948_),
    .A4(_1956_),
    .B1(_2345_),
    .X(_2346_));
 sky130_fd_sc_hd__a211o_1 _5464_ (.A1(_2339_),
    .A2(_2340_),
    .B1(_2344_),
    .C1(_2346_),
    .X(_2347_));
 sky130_fd_sc_hd__o32a_1 _5465_ (.A1(_1504_),
    .A2(_1419_),
    .A3(_1394_),
    .B1(_1421_),
    .B2(_1824_),
    .X(_2348_));
 sky130_fd_sc_hd__nor2_1 _5466_ (.A(_1417_),
    .B(_2348_),
    .Y(_2349_));
 sky130_fd_sc_hd__nor3_4 _5467_ (.A(_2338_),
    .B(_2347_),
    .C(_2349_),
    .Y(_2350_));
 sky130_fd_sc_hd__nor2_1 _5468_ (.A(_0859_),
    .B(_2350_),
    .Y(_2351_));
 sky130_fd_sc_hd__a211o_1 _5469_ (.A1(_2104_),
    .A2(\core_1.execute.alu_mul_div.mul_res[8] ),
    .B1(_2351_),
    .C1(_0831_),
    .X(_2352_));
 sky130_fd_sc_hd__a22o_2 _5470_ (.A1(\core_1.execute.alu_mul_div.div_cur[8] ),
    .A2(\core_1.execute.alu_mul_div.i_mod ),
    .B1(_2334_),
    .B2(_2352_),
    .X(_2353_));
 sky130_fd_sc_hd__mux2_1 _5471_ (.A0(_2333_),
    .A1(_2353_),
    .S(_2078_),
    .X(_2354_));
 sky130_fd_sc_hd__mux2_1 _5472_ (.A0(net208),
    .A1(_2354_),
    .S(_2081_),
    .X(_2355_));
 sky130_fd_sc_hd__mux2_1 _5473_ (.A0(\core_1.ew_data[8] ),
    .A1(_2355_),
    .S(_2101_),
    .X(_2356_));
 sky130_fd_sc_hd__clkbuf_1 _5474_ (.A(_2356_),
    .X(_0237_));
 sky130_fd_sc_hd__inv_2 _5475_ (.A(\core_1.ew_data[9] ),
    .Y(_2357_));
 sky130_fd_sc_hd__a21bo_1 _5476_ (.A1(\core_1.execute.alu_mul_div.div_res[9] ),
    .A2(_1313_),
    .B1_N(_1314_),
    .X(_2358_));
 sky130_fd_sc_hd__nand2_1 _5477_ (.A(_1896_),
    .B(_1898_),
    .Y(_2359_));
 sky130_fd_sc_hd__a21oi_1 _5478_ (.A1(_1902_),
    .A2(_2336_),
    .B1(_2359_),
    .Y(_2360_));
 sky130_fd_sc_hd__a31o_1 _5479_ (.A1(_2359_),
    .A2(_1902_),
    .A3(_2336_),
    .B1(_2047_),
    .X(_2361_));
 sky130_fd_sc_hd__inv_2 _5480_ (.A(_1895_),
    .Y(_2362_));
 sky130_fd_sc_hd__and2b_1 _5481_ (.A_N(_1899_),
    .B(_1957_),
    .X(_2363_));
 sky130_fd_sc_hd__xnor2_1 _5482_ (.A(_2362_),
    .B(_2363_),
    .Y(_2364_));
 sky130_fd_sc_hd__nand2_1 _5483_ (.A(_1421_),
    .B(_1826_),
    .Y(_2365_));
 sky130_fd_sc_hd__nand2_1 _5484_ (.A(_1823_),
    .B(_2232_),
    .Y(_2366_));
 sky130_fd_sc_hd__mux2_1 _5485_ (.A0(_1809_),
    .A1(_1836_),
    .S(_1406_),
    .X(_2367_));
 sky130_fd_sc_hd__and2_1 _5486_ (.A(_1828_),
    .B(_2367_),
    .X(_2368_));
 sky130_fd_sc_hd__a21oi_1 _5487_ (.A1(_1330_),
    .A2(_2308_),
    .B1(_2368_),
    .Y(_2369_));
 sky130_fd_sc_hd__o21a_1 _5488_ (.A1(_1823_),
    .A2(_2369_),
    .B1(_1845_),
    .X(_2370_));
 sky130_fd_sc_hd__a2bb2o_1 _5489_ (.A1_N(_1409_),
    .A2_N(_2365_),
    .B1(_2366_),
    .B2(_2370_),
    .X(_2371_));
 sky130_fd_sc_hd__inv_2 _5490_ (.A(_1503_),
    .Y(_2372_));
 sky130_fd_sc_hd__inv_2 _5491_ (.A(_1893_),
    .Y(_2373_));
 sky130_fd_sc_hd__a221o_1 _5492_ (.A1(\core_1.decode.oc_alu_mode[7] ),
    .A2(_1354_),
    .B1(_1445_),
    .B2(_1465_),
    .C1(_2341_),
    .X(_2374_));
 sky130_fd_sc_hd__a221o_1 _5493_ (.A1(\core_1.decode.oc_alu_mode[9] ),
    .A2(_2373_),
    .B1(_1894_),
    .B2(\core_1.decode.oc_alu_mode[2] ),
    .C1(_2374_),
    .X(_2375_));
 sky130_fd_sc_hd__a221o_1 _5494_ (.A1(\core_1.decode.oc_alu_mode[6] ),
    .A2(_2362_),
    .B1(_2340_),
    .B2(_2372_),
    .C1(_2375_),
    .X(_2376_));
 sky130_fd_sc_hd__a221o_1 _5495_ (.A1(_0780_),
    .A2(_2364_),
    .B1(_2371_),
    .B2(_2039_),
    .C1(_2376_),
    .X(_2377_));
 sky130_fd_sc_hd__o21ba_2 _5496_ (.A1(_2360_),
    .A2(_2361_),
    .B1_N(_2377_),
    .X(_2378_));
 sky130_fd_sc_hd__nor2_1 _5497_ (.A(_0860_),
    .B(_2378_),
    .Y(_2379_));
 sky130_fd_sc_hd__a211o_1 _5498_ (.A1(_0860_),
    .A2(\core_1.execute.alu_mul_div.mul_res[9] ),
    .B1(_2379_),
    .C1(_0831_),
    .X(_2380_));
 sky130_fd_sc_hd__a22o_4 _5499_ (.A1(\core_1.execute.alu_mul_div.div_cur[9] ),
    .A2(_0835_),
    .B1(_2358_),
    .B2(_2380_),
    .X(_2381_));
 sky130_fd_sc_hd__nand2_2 _5500_ (.A(\core_1.execute.sreg_irq_pc.o_d[9] ),
    .B(_1019_),
    .Y(_2382_));
 sky130_fd_sc_hd__a22o_1 _5501_ (.A1(net16),
    .A2(_2257_),
    .B1(_2293_),
    .B2(\core_1.execute.sreg_scratch.o_d[9] ),
    .X(_2383_));
 sky130_fd_sc_hd__a221o_1 _5502_ (.A1(\core_1.execute.sreg_priv_control.o_d[9] ),
    .A2(_1145_),
    .B1(_2294_),
    .B2(\core_1.execute.sreg_irq_pc.o_d[9] ),
    .C1(_2383_),
    .X(_2384_));
 sky130_fd_sc_hd__a22o_1 _5503_ (.A1(net87),
    .A2(_2256_),
    .B1(_2384_),
    .B2(_1138_),
    .X(_2385_));
 sky130_fd_sc_hd__nand2_1 _5504_ (.A(_1141_),
    .B(_2385_),
    .Y(_2386_));
 sky130_fd_sc_hd__or2b_1 _5505_ (.A(_2327_),
    .B_N(_2332_),
    .X(_2387_));
 sky130_fd_sc_hd__a21o_1 _5506_ (.A1(_2382_),
    .A2(_2386_),
    .B1(_2387_),
    .X(_2388_));
 sky130_fd_sc_hd__a31oi_2 _5507_ (.A1(_2387_),
    .A2(_2382_),
    .A3(_2386_),
    .B1(_2084_),
    .Y(_2389_));
 sky130_fd_sc_hd__a221oi_2 _5508_ (.A1(_2084_),
    .A2(_2381_),
    .B1(_2388_),
    .B2(_2389_),
    .C1(\core_1.dec_mem_access ),
    .Y(_2390_));
 sky130_fd_sc_hd__a211o_1 _5509_ (.A1(\core_1.dec_mem_access ),
    .A2(_0596_),
    .B1(_1796_),
    .C1(_2390_),
    .X(_2391_));
 sky130_fd_sc_hd__o21ai_1 _5510_ (.A1(_2357_),
    .A2(_1801_),
    .B1(_2391_),
    .Y(_0238_));
 sky130_fd_sc_hd__a22o_1 _5511_ (.A1(net2),
    .A2(_2257_),
    .B1(_2293_),
    .B2(\core_1.execute.sreg_scratch.o_d[10] ),
    .X(_2392_));
 sky130_fd_sc_hd__a221o_1 _5512_ (.A1(\core_1.execute.sreg_priv_control.o_d[10] ),
    .A2(_1145_),
    .B1(_2294_),
    .B2(\core_1.execute.sreg_irq_pc.o_d[10] ),
    .C1(_2392_),
    .X(_2393_));
 sky130_fd_sc_hd__a22o_1 _5513_ (.A1(net73),
    .A2(_2256_),
    .B1(_2393_),
    .B2(_1138_),
    .X(_2394_));
 sky130_fd_sc_hd__nand2_1 _5514_ (.A(\core_1.execute.sreg_irq_pc.o_d[10] ),
    .B(_1019_),
    .Y(_2395_));
 sky130_fd_sc_hd__a21bo_1 _5515_ (.A1(_1141_),
    .A2(_2394_),
    .B1_N(_2395_),
    .X(_2396_));
 sky130_fd_sc_hd__xnor2_1 _5516_ (.A(_2388_),
    .B(_2396_),
    .Y(_2397_));
 sky130_fd_sc_hd__a21bo_1 _5517_ (.A1(\core_1.execute.alu_mul_div.div_res[10] ),
    .A2(_1312_),
    .B1_N(_0727_),
    .X(_2398_));
 sky130_fd_sc_hd__a21oi_2 _5518_ (.A1(_1905_),
    .A2(_1906_),
    .B1(_1912_),
    .Y(_2399_));
 sky130_fd_sc_hd__and3_1 _5519_ (.A(_1905_),
    .B(_1906_),
    .C(_1912_),
    .X(_2400_));
 sky130_fd_sc_hd__nor2_1 _5520_ (.A(_2399_),
    .B(_2400_),
    .Y(_2401_));
 sky130_fd_sc_hd__inv_2 _5521_ (.A(_1909_),
    .Y(_2402_));
 sky130_fd_sc_hd__inv_2 _5522_ (.A(_1908_),
    .Y(_2403_));
 sky130_fd_sc_hd__a221o_1 _5523_ (.A1(_0846_),
    .A2(_1352_),
    .B1(_2403_),
    .B2(_0814_),
    .C1(_2341_),
    .X(_2404_));
 sky130_fd_sc_hd__a221o_1 _5524_ (.A1(_0839_),
    .A2(_1907_),
    .B1(_2402_),
    .B2(_0832_),
    .C1(_2404_),
    .X(_2405_));
 sky130_fd_sc_hd__a21o_1 _5525_ (.A1(_1935_),
    .A2(_1957_),
    .B1(_1893_),
    .X(_2406_));
 sky130_fd_sc_hd__nand2_1 _5526_ (.A(_1909_),
    .B(_2406_),
    .Y(_2407_));
 sky130_fd_sc_hd__nor2_1 _5527_ (.A(_2046_),
    .B(_1958_),
    .Y(_2408_));
 sky130_fd_sc_hd__a22o_1 _5528_ (.A1(_2110_),
    .A2(_2340_),
    .B1(_2407_),
    .B2(_2408_),
    .X(_2409_));
 sky130_fd_sc_hd__a211o_1 _5529_ (.A1(_0863_),
    .A2(_2401_),
    .B1(_2405_),
    .C1(_2409_),
    .X(_2410_));
 sky130_fd_sc_hd__mux2_1 _5530_ (.A0(_1810_),
    .A1(_1838_),
    .S(_1829_),
    .X(_2411_));
 sky130_fd_sc_hd__mux2_1 _5531_ (.A0(_2267_),
    .A1(_2411_),
    .S(_1826_),
    .X(_2412_));
 sky130_fd_sc_hd__or3_1 _5532_ (.A(_1845_),
    .B(_1823_),
    .C(_2266_),
    .X(_2413_));
 sky130_fd_sc_hd__o21a_1 _5533_ (.A1(_1421_),
    .A2(_2412_),
    .B1(_2413_),
    .X(_2414_));
 sky130_fd_sc_hd__nor2_1 _5534_ (.A(_1417_),
    .B(_2414_),
    .Y(_2415_));
 sky130_fd_sc_hd__a211o_2 _5535_ (.A1(_1445_),
    .A2(_1457_),
    .B1(_2410_),
    .C1(_2415_),
    .X(_2416_));
 sky130_fd_sc_hd__a21o_1 _5536_ (.A1(_0859_),
    .A2(\core_1.execute.alu_mul_div.mul_res[10] ),
    .B1(\core_1.execute.alu_mul_div.i_div ),
    .X(_2417_));
 sky130_fd_sc_hd__a21o_1 _5537_ (.A1(_1316_),
    .A2(_2416_),
    .B1(_2417_),
    .X(_2418_));
 sky130_fd_sc_hd__a22o_4 _5538_ (.A1(\core_1.execute.alu_mul_div.div_cur[10] ),
    .A2(\core_1.execute.alu_mul_div.i_mod ),
    .B1(_2398_),
    .B2(_2418_),
    .X(_2419_));
 sky130_fd_sc_hd__mux2_1 _5539_ (.A0(_2397_),
    .A1(_2419_),
    .S(_2078_),
    .X(_2420_));
 sky130_fd_sc_hd__mux2_1 _5540_ (.A0(net195),
    .A1(_2420_),
    .S(_2081_),
    .X(_2421_));
 sky130_fd_sc_hd__mux2_1 _5541_ (.A0(\core_1.ew_data[10] ),
    .A1(_2421_),
    .S(_2101_),
    .X(_2422_));
 sky130_fd_sc_hd__clkbuf_1 _5542_ (.A(_2422_),
    .X(_0239_));
 sky130_fd_sc_hd__a21bo_1 _5543_ (.A1(\core_1.execute.alu_mul_div.div_res[11] ),
    .A2(_1313_),
    .B1_N(_1314_),
    .X(_2423_));
 sky130_fd_sc_hd__o21ai_1 _5544_ (.A1(_1907_),
    .A2(_1958_),
    .B1(_1915_),
    .Y(_2424_));
 sky130_fd_sc_hd__o31a_1 _5545_ (.A1(_1915_),
    .A2(_1907_),
    .A3(_1958_),
    .B1(_0780_),
    .X(_2425_));
 sky130_fd_sc_hd__mux2_1 _5546_ (.A0(_1837_),
    .A1(_1839_),
    .S(_1406_),
    .X(_2426_));
 sky130_fd_sc_hd__mux2_1 _5547_ (.A0(_2367_),
    .A1(_2426_),
    .S(_1829_),
    .X(_2427_));
 sky130_fd_sc_hd__nand2_1 _5548_ (.A(_1826_),
    .B(_2427_),
    .Y(_2428_));
 sky130_fd_sc_hd__a21oi_1 _5549_ (.A1(_1823_),
    .A2(_2309_),
    .B1(_1421_),
    .Y(_2429_));
 sky130_fd_sc_hd__a2bb2o_1 _5550_ (.A1_N(_2158_),
    .A2_N(_2365_),
    .B1(_2428_),
    .B2(_2429_),
    .X(_2430_));
 sky130_fd_sc_hd__o21ai_1 _5551_ (.A1(_1505_),
    .A2(_2313_),
    .B1(_2161_),
    .Y(_2431_));
 sky130_fd_sc_hd__a221o_1 _5552_ (.A1(_0846_),
    .A2(_1353_),
    .B1(_1445_),
    .B2(_1734_),
    .C1(_2341_),
    .X(_2432_));
 sky130_fd_sc_hd__a221o_1 _5553_ (.A1(_0814_),
    .A2(_1959_),
    .B1(_1914_),
    .B2(_0839_),
    .C1(_2432_),
    .X(_2433_));
 sky130_fd_sc_hd__a221o_1 _5554_ (.A1(_0832_),
    .A2(_1915_),
    .B1(_2431_),
    .B2(_2340_),
    .C1(_2433_),
    .X(_2434_));
 sky130_fd_sc_hd__a21o_1 _5555_ (.A1(_2039_),
    .A2(_2430_),
    .B1(_2434_),
    .X(_2435_));
 sky130_fd_sc_hd__or3_1 _5556_ (.A(_1918_),
    .B(_1911_),
    .C(_2399_),
    .X(_2436_));
 sky130_fd_sc_hd__o21ai_1 _5557_ (.A1(_1911_),
    .A2(_2399_),
    .B1(_1918_),
    .Y(_2437_));
 sky130_fd_sc_hd__and3_1 _5558_ (.A(_0863_),
    .B(_2436_),
    .C(_2437_),
    .X(_2438_));
 sky130_fd_sc_hd__a211oi_4 _5559_ (.A1(_2424_),
    .A2(_2425_),
    .B1(_2435_),
    .C1(_2438_),
    .Y(_2439_));
 sky130_fd_sc_hd__nor2_1 _5560_ (.A(_2104_),
    .B(_2439_),
    .Y(_2440_));
 sky130_fd_sc_hd__a211o_1 _5561_ (.A1(_0860_),
    .A2(\core_1.execute.alu_mul_div.mul_res[11] ),
    .B1(_2440_),
    .C1(_0831_),
    .X(_2441_));
 sky130_fd_sc_hd__a22o_4 _5562_ (.A1(\core_1.execute.alu_mul_div.div_cur[11] ),
    .A2(_0835_),
    .B1(_2423_),
    .B2(_2441_),
    .X(_2442_));
 sky130_fd_sc_hd__nand2_1 _5563_ (.A(\core_1.execute.sreg_irq_pc.o_d[11] ),
    .B(_1019_),
    .Y(_2443_));
 sky130_fd_sc_hd__nand2_1 _5564_ (.A(net74),
    .B(_2256_),
    .Y(_2444_));
 sky130_fd_sc_hd__a22o_1 _5565_ (.A1(net3),
    .A2(_2257_),
    .B1(_2293_),
    .B2(\core_1.execute.sreg_scratch.o_d[11] ),
    .X(_2445_));
 sky130_fd_sc_hd__a221o_1 _5566_ (.A1(\core_1.execute.sreg_priv_control.o_d[11] ),
    .A2(_1145_),
    .B1(_2294_),
    .B2(\core_1.execute.sreg_irq_pc.o_d[11] ),
    .C1(_2445_),
    .X(_2446_));
 sky130_fd_sc_hd__nand2_1 _5567_ (.A(_1138_),
    .B(_2446_),
    .Y(_2447_));
 sky130_fd_sc_hd__a21o_1 _5568_ (.A1(_2444_),
    .A2(_2447_),
    .B1(_1019_),
    .X(_2448_));
 sky130_fd_sc_hd__or2b_1 _5569_ (.A(_2388_),
    .B_N(_2396_),
    .X(_2449_));
 sky130_fd_sc_hd__a21o_1 _5570_ (.A1(_2443_),
    .A2(_2448_),
    .B1(_2449_),
    .X(_2450_));
 sky130_fd_sc_hd__a31oi_1 _5571_ (.A1(_2449_),
    .A2(_2443_),
    .A3(_2448_),
    .B1(_2077_),
    .Y(_2451_));
 sky130_fd_sc_hd__a22o_1 _5572_ (.A1(_2084_),
    .A2(_2442_),
    .B1(_2450_),
    .B2(_2451_),
    .X(_2452_));
 sky130_fd_sc_hd__mux2_1 _5573_ (.A0(net196),
    .A1(_2452_),
    .S(_2080_),
    .X(_2453_));
 sky130_fd_sc_hd__mux2_1 _5574_ (.A0(\core_1.ew_data[11] ),
    .A1(_2453_),
    .S(_2101_),
    .X(_2454_));
 sky130_fd_sc_hd__clkbuf_1 _5575_ (.A(_2454_),
    .X(_0240_));
 sky130_fd_sc_hd__a22o_1 _5576_ (.A1(net4),
    .A2(_2257_),
    .B1(_2293_),
    .B2(\core_1.execute.sreg_scratch.o_d[12] ),
    .X(_2455_));
 sky130_fd_sc_hd__a221o_1 _5577_ (.A1(\core_1.execute.sreg_priv_control.o_d[12] ),
    .A2(_1145_),
    .B1(_2294_),
    .B2(\core_1.execute.sreg_irq_pc.o_d[12] ),
    .C1(_2455_),
    .X(_2456_));
 sky130_fd_sc_hd__a22o_1 _5578_ (.A1(net75),
    .A2(_2256_),
    .B1(_2456_),
    .B2(_1138_),
    .X(_2457_));
 sky130_fd_sc_hd__nand2_1 _5579_ (.A(\core_1.execute.sreg_irq_pc.o_d[12] ),
    .B(_1019_),
    .Y(_2458_));
 sky130_fd_sc_hd__a21bo_1 _5580_ (.A1(_1141_),
    .A2(_2457_),
    .B1_N(_2458_),
    .X(_2459_));
 sky130_fd_sc_hd__xnor2_1 _5581_ (.A(_2450_),
    .B(_2459_),
    .Y(_2460_));
 sky130_fd_sc_hd__a21bo_1 _5582_ (.A1(\core_1.execute.alu_mul_div.div_res[12] ),
    .A2(_1312_),
    .B1_N(_0727_),
    .X(_2461_));
 sky130_fd_sc_hd__a211o_1 _5583_ (.A1(_1918_),
    .A2(_2399_),
    .B1(_1921_),
    .C1(_1924_),
    .X(_2462_));
 sky130_fd_sc_hd__o31a_1 _5584_ (.A1(_1914_),
    .A2(_1907_),
    .A3(_1958_),
    .B1(_1959_),
    .X(_2463_));
 sky130_fd_sc_hd__nor2_1 _5585_ (.A(_1960_),
    .B(_2463_),
    .Y(_2464_));
 sky130_fd_sc_hd__nor2_1 _5586_ (.A(_1961_),
    .B(_2464_),
    .Y(_2465_));
 sky130_fd_sc_hd__nor2_1 _5587_ (.A(_2273_),
    .B(_1864_),
    .Y(_2466_));
 sky130_fd_sc_hd__inv_2 _5588_ (.A(_1863_),
    .Y(_2467_));
 sky130_fd_sc_hd__a221o_1 _5589_ (.A1(\core_1.decode.oc_alu_mode[7] ),
    .A2(_1373_),
    .B1(_1445_),
    .B2(_1477_),
    .C1(_2341_),
    .X(_2468_));
 sky130_fd_sc_hd__a221o_1 _5590_ (.A1(\core_1.decode.oc_alu_mode[2] ),
    .A2(_1862_),
    .B1(_2467_),
    .B2(\core_1.decode.oc_alu_mode[9] ),
    .C1(_2468_),
    .X(_2469_));
 sky130_fd_sc_hd__a211o_1 _5591_ (.A1(_2206_),
    .A2(_2340_),
    .B1(_2466_),
    .C1(_2469_),
    .X(_2470_));
 sky130_fd_sc_hd__mux4_1 _5592_ (.A0(_1810_),
    .A1(_1814_),
    .A2(_1841_),
    .A3(_1838_),
    .S0(_1330_),
    .S1(_1424_),
    .X(_2471_));
 sky130_fd_sc_hd__nand2_1 _5593_ (.A(_1845_),
    .B(_2471_),
    .Y(_2472_));
 sky130_fd_sc_hd__o211a_1 _5594_ (.A1(_1845_),
    .A2(_2199_),
    .B1(_2472_),
    .C1(_2039_),
    .X(_2473_));
 sky130_fd_sc_hd__a211o_1 _5595_ (.A1(_0780_),
    .A2(_2465_),
    .B1(_2470_),
    .C1(_2473_),
    .X(_2474_));
 sky130_fd_sc_hd__a31oi_4 _5596_ (.A1(_0863_),
    .A2(_1925_),
    .A3(_2462_),
    .B1(_2474_),
    .Y(_2475_));
 sky130_fd_sc_hd__nor2_1 _5597_ (.A(_0859_),
    .B(_2475_),
    .Y(_2476_));
 sky130_fd_sc_hd__a211o_1 _5598_ (.A1(_2104_),
    .A2(\core_1.execute.alu_mul_div.mul_res[12] ),
    .B1(_2476_),
    .C1(\core_1.execute.alu_mul_div.i_div ),
    .X(_2477_));
 sky130_fd_sc_hd__a22o_4 _5599_ (.A1(\core_1.execute.alu_mul_div.div_cur[12] ),
    .A2(\core_1.execute.alu_mul_div.i_mod ),
    .B1(_2461_),
    .B2(_2477_),
    .X(_2478_));
 sky130_fd_sc_hd__mux2_1 _5600_ (.A0(_2460_),
    .A1(_2478_),
    .S(_2078_),
    .X(_2479_));
 sky130_fd_sc_hd__mux2_1 _5601_ (.A0(net197),
    .A1(_2479_),
    .S(_2080_),
    .X(_2480_));
 sky130_fd_sc_hd__buf_6 _5602_ (.A(_1800_),
    .X(_2481_));
 sky130_fd_sc_hd__mux2_1 _5603_ (.A0(\core_1.ew_data[12] ),
    .A1(_2480_),
    .S(_2481_),
    .X(_2482_));
 sky130_fd_sc_hd__clkbuf_1 _5604_ (.A(_2482_),
    .X(_0241_));
 sky130_fd_sc_hd__a21bo_1 _5605_ (.A1(\core_1.execute.alu_mul_div.div_res[13] ),
    .A2(_1313_),
    .B1_N(_1314_),
    .X(_2483_));
 sky130_fd_sc_hd__inv_2 _5606_ (.A(_1861_),
    .Y(_2484_));
 sky130_fd_sc_hd__a211o_1 _5607_ (.A1(_1865_),
    .A2(_1925_),
    .B1(_2484_),
    .C1(_1926_),
    .X(_2485_));
 sky130_fd_sc_hd__o211ai_2 _5608_ (.A1(_2484_),
    .A2(_1926_),
    .B1(_1865_),
    .C1(_1925_),
    .Y(_2486_));
 sky130_fd_sc_hd__or2_1 _5609_ (.A(_1862_),
    .B(_1961_),
    .X(_2487_));
 sky130_fd_sc_hd__xnor2_1 _5610_ (.A(_1860_),
    .B(_2487_),
    .Y(_2488_));
 sky130_fd_sc_hd__mux2_1 _5611_ (.A0(_1840_),
    .A1(_1832_),
    .S(_1406_),
    .X(_2489_));
 sky130_fd_sc_hd__mux2_1 _5612_ (.A0(_2426_),
    .A1(_2489_),
    .S(_1828_),
    .X(_2490_));
 sky130_fd_sc_hd__clkinv_2 _5613_ (.A(_2490_),
    .Y(_2491_));
 sky130_fd_sc_hd__mux2_1 _5614_ (.A0(_2369_),
    .A1(_2491_),
    .S(_1826_),
    .X(_2492_));
 sky130_fd_sc_hd__nor2_1 _5615_ (.A(_2273_),
    .B(_1860_),
    .Y(_2493_));
 sky130_fd_sc_hd__a221o_1 _5616_ (.A1(\core_1.decode.oc_alu_mode[7] ),
    .A2(_1371_),
    .B1(_1445_),
    .B2(_1493_),
    .C1(_2341_),
    .X(_2494_));
 sky130_fd_sc_hd__a221o_1 _5617_ (.A1(\core_1.decode.oc_alu_mode[9] ),
    .A2(_1858_),
    .B1(_1934_),
    .B2(\core_1.decode.oc_alu_mode[2] ),
    .C1(_2494_),
    .X(_2495_));
 sky130_fd_sc_hd__a211oi_1 _5618_ (.A1(_2243_),
    .A2(_2340_),
    .B1(_2493_),
    .C1(_2495_),
    .Y(_2496_));
 sky130_fd_sc_hd__o31ai_1 _5619_ (.A1(_1417_),
    .A2(_1845_),
    .A3(_2233_),
    .B1(_2496_),
    .Y(_2497_));
 sky130_fd_sc_hd__a221o_1 _5620_ (.A1(_0780_),
    .A2(_2488_),
    .B1(_2492_),
    .B2(_1422_),
    .C1(_2497_),
    .X(_2498_));
 sky130_fd_sc_hd__a31oi_4 _5621_ (.A1(_0863_),
    .A2(_2485_),
    .A3(_2486_),
    .B1(_2498_),
    .Y(_2499_));
 sky130_fd_sc_hd__nor2_1 _5622_ (.A(_2104_),
    .B(_2499_),
    .Y(_2500_));
 sky130_fd_sc_hd__a211o_1 _5623_ (.A1(_0860_),
    .A2(\core_1.execute.alu_mul_div.mul_res[13] ),
    .B1(_2500_),
    .C1(_0831_),
    .X(_2501_));
 sky130_fd_sc_hd__a22o_4 _5624_ (.A1(\core_1.execute.alu_mul_div.div_cur[13] ),
    .A2(_0835_),
    .B1(_2483_),
    .B2(_2501_),
    .X(_2502_));
 sky130_fd_sc_hd__nor2b_1 _5625_ (.A(_2450_),
    .B_N(_2459_),
    .Y(_2503_));
 sky130_fd_sc_hd__a22o_1 _5626_ (.A1(\core_1.execute.sreg_priv_control.o_d[13] ),
    .A2(_1145_),
    .B1(_2257_),
    .B2(net5),
    .X(_2504_));
 sky130_fd_sc_hd__a221o_1 _5627_ (.A1(\core_1.execute.sreg_irq_pc.o_d[13] ),
    .A2(_2294_),
    .B1(_2293_),
    .B2(\core_1.execute.sreg_scratch.o_d[13] ),
    .C1(_2504_),
    .X(_2505_));
 sky130_fd_sc_hd__or2_1 _5628_ (.A(_2030_),
    .B(_2505_),
    .X(_2506_));
 sky130_fd_sc_hd__a22o_1 _5629_ (.A1(net76),
    .A2(_2256_),
    .B1(_2506_),
    .B2(_1138_),
    .X(_2507_));
 sky130_fd_sc_hd__mux2_2 _5630_ (.A0(\core_1.execute.sreg_irq_pc.o_d[13] ),
    .A1(_2507_),
    .S(_1141_),
    .X(_2508_));
 sky130_fd_sc_hd__xnor2_1 _5631_ (.A(_2503_),
    .B(_2508_),
    .Y(_2509_));
 sky130_fd_sc_hd__nor2_1 _5632_ (.A(_2084_),
    .B(_2509_),
    .Y(_2510_));
 sky130_fd_sc_hd__a21o_1 _5633_ (.A1(_2084_),
    .A2(_2502_),
    .B1(_2510_),
    .X(_2511_));
 sky130_fd_sc_hd__mux2_1 _5634_ (.A0(net198),
    .A1(_2511_),
    .S(_2080_),
    .X(_2512_));
 sky130_fd_sc_hd__mux2_1 _5635_ (.A0(\core_1.ew_data[13] ),
    .A1(_2512_),
    .S(_2481_),
    .X(_2513_));
 sky130_fd_sc_hd__clkbuf_1 _5636_ (.A(_2513_),
    .X(_0242_));
 sky130_fd_sc_hd__nand2_1 _5637_ (.A(_2503_),
    .B(_2508_),
    .Y(_2514_));
 sky130_fd_sc_hd__a22o_1 _5638_ (.A1(\core_1.execute.sreg_priv_control.o_d[14] ),
    .A2(_1145_),
    .B1(_2257_),
    .B2(net6),
    .X(_2515_));
 sky130_fd_sc_hd__a221o_1 _5639_ (.A1(\core_1.execute.sreg_irq_pc.o_d[14] ),
    .A2(_2294_),
    .B1(_2293_),
    .B2(\core_1.execute.sreg_scratch.o_d[14] ),
    .C1(_2515_),
    .X(_2516_));
 sky130_fd_sc_hd__nor2_1 _5640_ (.A(_2030_),
    .B(_2516_),
    .Y(_2517_));
 sky130_fd_sc_hd__o2bb2a_1 _5641_ (.A1_N(net77),
    .A2_N(_2256_),
    .B1(_2517_),
    .B2(\core_1.dec_sreg_jal_over ),
    .X(_2518_));
 sky130_fd_sc_hd__nand2_1 _5642_ (.A(\core_1.execute.sreg_irq_pc.o_d[14] ),
    .B(_1019_),
    .Y(_2519_));
 sky130_fd_sc_hd__o21ai_2 _5643_ (.A1(_1019_),
    .A2(_2518_),
    .B1(_2519_),
    .Y(_2520_));
 sky130_fd_sc_hd__xnor2_1 _5644_ (.A(_2514_),
    .B(_2520_),
    .Y(_2521_));
 sky130_fd_sc_hd__nor2_1 _5645_ (.A(_1855_),
    .B(_1962_),
    .Y(_2522_));
 sky130_fd_sc_hd__nor2_1 _5646_ (.A(_1963_),
    .B(_2522_),
    .Y(_2523_));
 sky130_fd_sc_hd__a221o_1 _5647_ (.A1(_0846_),
    .A2(_1351_),
    .B1(_1854_),
    .B2(_0814_),
    .C1(_2341_),
    .X(_2524_));
 sky130_fd_sc_hd__a221o_1 _5648_ (.A1(_0839_),
    .A2(_1853_),
    .B1(_1855_),
    .B2(_0832_),
    .C1(_2524_),
    .X(_2525_));
 sky130_fd_sc_hd__a31o_1 _5649_ (.A1(_1861_),
    .A2(_1865_),
    .A3(_1925_),
    .B1(_1926_),
    .X(_2526_));
 sky130_fd_sc_hd__nand2_1 _5650_ (.A(_1928_),
    .B(_2526_),
    .Y(_2527_));
 sky130_fd_sc_hd__and3b_1 _5651_ (.A_N(_2107_),
    .B(_2340_),
    .C(_1418_),
    .X(_2528_));
 sky130_fd_sc_hd__a31o_1 _5652_ (.A1(_0862_),
    .A2(_1929_),
    .A3(_2527_),
    .B1(_2528_),
    .X(_2529_));
 sky130_fd_sc_hd__mux2_1 _5653_ (.A0(_1841_),
    .A1(_1833_),
    .S(_1829_),
    .X(_2530_));
 sky130_fd_sc_hd__mux4_1 _5654_ (.A0(_2266_),
    .A1(_2267_),
    .A2(_2411_),
    .A3(_2530_),
    .S0(_1826_),
    .S1(_1845_),
    .X(_2531_));
 sky130_fd_sc_hd__nor2_1 _5655_ (.A(_1417_),
    .B(_2531_),
    .Y(_2532_));
 sky130_fd_sc_hd__a2111o_1 _5656_ (.A1(_1445_),
    .A2(_1745_),
    .B1(_2525_),
    .C1(_2529_),
    .D1(_2532_),
    .X(_2533_));
 sky130_fd_sc_hd__a21oi_2 _5657_ (.A1(_0780_),
    .A2(_2523_),
    .B1(_2533_),
    .Y(_2534_));
 sky130_fd_sc_hd__nor2_1 _5658_ (.A(_2104_),
    .B(_2534_),
    .Y(_2535_));
 sky130_fd_sc_hd__a211o_1 _5659_ (.A1(_0860_),
    .A2(\core_1.execute.alu_mul_div.mul_res[14] ),
    .B1(_2535_),
    .C1(_0831_),
    .X(_2536_));
 sky130_fd_sc_hd__a21bo_1 _5660_ (.A1(\core_1.execute.alu_mul_div.div_res[14] ),
    .A2(_1312_),
    .B1_N(_0727_),
    .X(_2537_));
 sky130_fd_sc_hd__a22o_4 _5661_ (.A1(\core_1.execute.alu_mul_div.div_cur[14] ),
    .A2(\core_1.execute.alu_mul_div.i_mod ),
    .B1(_2536_),
    .B2(_2537_),
    .X(_2538_));
 sky130_fd_sc_hd__mux2_1 _5662_ (.A0(_2521_),
    .A1(_2538_),
    .S(_2078_),
    .X(_2539_));
 sky130_fd_sc_hd__mux2_1 _5663_ (.A0(net199),
    .A1(_2539_),
    .S(_2080_),
    .X(_2540_));
 sky130_fd_sc_hd__mux2_1 _5664_ (.A0(\core_1.ew_data[14] ),
    .A1(_2540_),
    .S(_2481_),
    .X(_2541_));
 sky130_fd_sc_hd__clkbuf_1 _5665_ (.A(_2541_),
    .X(_0243_));
 sky130_fd_sc_hd__nand2_1 _5666_ (.A(_1827_),
    .B(_1831_),
    .Y(_2542_));
 sky130_fd_sc_hd__o21ai_1 _5667_ (.A1(_1827_),
    .A2(_1830_),
    .B1(_2542_),
    .Y(_2543_));
 sky130_fd_sc_hd__mux2_1 _5668_ (.A0(_2489_),
    .A1(_2543_),
    .S(_1829_),
    .X(_2544_));
 sky130_fd_sc_hd__mux4_1 _5669_ (.A0(_2158_),
    .A1(_2309_),
    .A2(_2427_),
    .A3(_2544_),
    .S0(_1826_),
    .S1(_1845_),
    .X(_2545_));
 sky130_fd_sc_hd__inv_2 _5670_ (.A(_2545_),
    .Y(_2546_));
 sky130_fd_sc_hd__a211oi_1 _5671_ (.A1(_1857_),
    .A2(_1929_),
    .B1(_1932_),
    .C1(_1852_),
    .Y(_2547_));
 sky130_fd_sc_hd__o211a_1 _5672_ (.A1(_1852_),
    .A2(_1932_),
    .B1(_1929_),
    .C1(_1857_),
    .X(_2548_));
 sky130_fd_sc_hd__nor2_1 _5673_ (.A(_2547_),
    .B(_2548_),
    .Y(_2549_));
 sky130_fd_sc_hd__nor2_2 _5674_ (.A(_1849_),
    .B(_1850_),
    .Y(_2550_));
 sky130_fd_sc_hd__o21ai_1 _5675_ (.A1(_1853_),
    .A2(_1963_),
    .B1(_2550_),
    .Y(_2551_));
 sky130_fd_sc_hd__o31a_1 _5676_ (.A1(_2550_),
    .A2(_1853_),
    .A3(_1963_),
    .B1(\core_1.decode.oc_alu_mode[4] ),
    .X(_2552_));
 sky130_fd_sc_hd__a22o_1 _5677_ (.A1(_0862_),
    .A2(_2549_),
    .B1(_2551_),
    .B2(_2552_),
    .X(_2553_));
 sky130_fd_sc_hd__a221o_1 _5678_ (.A1(_0846_),
    .A2(_1804_),
    .B1(_1964_),
    .B2(_0814_),
    .C1(_2341_),
    .X(_2554_));
 sky130_fd_sc_hd__a21o_1 _5679_ (.A1(_0839_),
    .A2(_1850_),
    .B1(_2554_),
    .X(_2555_));
 sky130_fd_sc_hd__a221o_1 _5680_ (.A1(_0832_),
    .A2(_2550_),
    .B1(_2312_),
    .B2(_2340_),
    .C1(_2555_),
    .X(_2556_));
 sky130_fd_sc_hd__a211o_1 _5681_ (.A1(_2039_),
    .A2(_2546_),
    .B1(_2553_),
    .C1(_2556_),
    .X(_2557_));
 sky130_fd_sc_hd__a21o_2 _5682_ (.A1(_1733_),
    .A2(_1445_),
    .B1(_2557_),
    .X(_2558_));
 sky130_fd_sc_hd__a21o_1 _5683_ (.A1(_0859_),
    .A2(\core_1.execute.alu_mul_div.mul_res[15] ),
    .B1(\core_1.execute.alu_mul_div.i_div ),
    .X(_2559_));
 sky130_fd_sc_hd__a21o_1 _5684_ (.A1(_1316_),
    .A2(_2558_),
    .B1(_2559_),
    .X(_2560_));
 sky130_fd_sc_hd__a21bo_1 _5685_ (.A1(\core_1.execute.alu_mul_div.div_res[15] ),
    .A2(_1313_),
    .B1_N(_1314_),
    .X(_2561_));
 sky130_fd_sc_hd__a22o_4 _5686_ (.A1(\core_1.execute.alu_mul_div.div_cur[15] ),
    .A2(_0835_),
    .B1(_2560_),
    .B2(_2561_),
    .X(_2562_));
 sky130_fd_sc_hd__and3_1 _5687_ (.A(_2503_),
    .B(_2508_),
    .C(_2520_),
    .X(_2563_));
 sky130_fd_sc_hd__a221o_1 _5688_ (.A1(net7),
    .A2(_2257_),
    .B1(_2293_),
    .B2(\core_1.execute.sreg_scratch.o_d[15] ),
    .C1(_2030_),
    .X(_2564_));
 sky130_fd_sc_hd__a221o_1 _5689_ (.A1(\core_1.execute.sreg_priv_control.o_d[15] ),
    .A2(_1145_),
    .B1(_2294_),
    .B2(\core_1.execute.sreg_irq_pc.o_d[15] ),
    .C1(_2564_),
    .X(_2565_));
 sky130_fd_sc_hd__a22o_1 _5690_ (.A1(net78),
    .A2(_2256_),
    .B1(_2565_),
    .B2(_1138_),
    .X(_2566_));
 sky130_fd_sc_hd__mux2_1 _5691_ (.A0(\core_1.execute.sreg_irq_pc.o_d[15] ),
    .A1(_2566_),
    .S(_1141_),
    .X(_2567_));
 sky130_fd_sc_hd__or2_1 _5692_ (.A(_2563_),
    .B(_2567_),
    .X(_2568_));
 sky130_fd_sc_hd__a21oi_1 _5693_ (.A1(_2563_),
    .A2(_2567_),
    .B1(_2078_),
    .Y(_2569_));
 sky130_fd_sc_hd__a22o_1 _5694_ (.A1(_2084_),
    .A2(_2562_),
    .B1(_2568_),
    .B2(_2569_),
    .X(_2570_));
 sky130_fd_sc_hd__mux2_1 _5695_ (.A0(net200),
    .A1(_2570_),
    .S(_2080_),
    .X(_2571_));
 sky130_fd_sc_hd__mux2_1 _5696_ (.A0(\core_1.ew_data[15] ),
    .A1(_2571_),
    .S(_2481_),
    .X(_2572_));
 sky130_fd_sc_hd__clkbuf_1 _5697_ (.A(_2572_),
    .X(_0244_));
 sky130_fd_sc_hd__mux2_1 _5698_ (.A0(\core_1.ew_addr[0] ),
    .A1(_2076_),
    .S(_2481_),
    .X(_2573_));
 sky130_fd_sc_hd__clkbuf_1 _5699_ (.A(_2573_),
    .X(_0245_));
 sky130_fd_sc_hd__mux2_1 _5700_ (.A0(net116),
    .A1(_1573_),
    .S(_2481_),
    .X(_2574_));
 sky130_fd_sc_hd__clkbuf_1 _5701_ (.A(_2574_),
    .X(_0246_));
 sky130_fd_sc_hd__mux2_1 _5702_ (.A0(net123),
    .A1(_2131_),
    .S(_2481_),
    .X(_2575_));
 sky130_fd_sc_hd__clkbuf_1 _5703_ (.A(_2575_),
    .X(_0247_));
 sky130_fd_sc_hd__mux2_1 _5704_ (.A0(net124),
    .A1(_2180_),
    .S(_2481_),
    .X(_2576_));
 sky130_fd_sc_hd__clkbuf_1 _5705_ (.A(_2576_),
    .X(_0248_));
 sky130_fd_sc_hd__mux2_1 _5706_ (.A0(net125),
    .A1(_2216_),
    .S(_2481_),
    .X(_2577_));
 sky130_fd_sc_hd__clkbuf_1 _5707_ (.A(_2577_),
    .X(_0249_));
 sky130_fd_sc_hd__mux2_1 _5708_ (.A0(net126),
    .A1(_2252_),
    .S(_2481_),
    .X(_2578_));
 sky130_fd_sc_hd__clkbuf_1 _5709_ (.A(_2578_),
    .X(_0250_));
 sky130_fd_sc_hd__buf_4 _5710_ (.A(_1800_),
    .X(_2579_));
 sky130_fd_sc_hd__mux2_1 _5711_ (.A0(net127),
    .A1(_2288_),
    .S(_2579_),
    .X(_2580_));
 sky130_fd_sc_hd__clkbuf_1 _5712_ (.A(_2580_),
    .X(_0251_));
 sky130_fd_sc_hd__mux2_1 _5713_ (.A0(net128),
    .A1(_2323_),
    .S(_2579_),
    .X(_2581_));
 sky130_fd_sc_hd__clkbuf_1 _5714_ (.A(_2581_),
    .X(_0252_));
 sky130_fd_sc_hd__mux2_1 _5715_ (.A0(net129),
    .A1(_2353_),
    .S(_2579_),
    .X(_2582_));
 sky130_fd_sc_hd__clkbuf_1 _5716_ (.A(_2582_),
    .X(_0253_));
 sky130_fd_sc_hd__mux2_1 _5717_ (.A0(net130),
    .A1(_2381_),
    .S(_2579_),
    .X(_2583_));
 sky130_fd_sc_hd__clkbuf_1 _5718_ (.A(_2583_),
    .X(_0254_));
 sky130_fd_sc_hd__mux2_1 _5719_ (.A0(net131),
    .A1(_2419_),
    .S(_2579_),
    .X(_2584_));
 sky130_fd_sc_hd__clkbuf_1 _5720_ (.A(_2584_),
    .X(_0255_));
 sky130_fd_sc_hd__mux2_1 _5721_ (.A0(net117),
    .A1(_2442_),
    .S(_2579_),
    .X(_2585_));
 sky130_fd_sc_hd__clkbuf_1 _5722_ (.A(_2585_),
    .X(_0256_));
 sky130_fd_sc_hd__mux2_1 _5723_ (.A0(net118),
    .A1(_2478_),
    .S(_2579_),
    .X(_2586_));
 sky130_fd_sc_hd__clkbuf_1 _5724_ (.A(_2586_),
    .X(_0257_));
 sky130_fd_sc_hd__mux2_1 _5725_ (.A0(net119),
    .A1(_2502_),
    .S(_2579_),
    .X(_2587_));
 sky130_fd_sc_hd__clkbuf_1 _5726_ (.A(_2587_),
    .X(_0258_));
 sky130_fd_sc_hd__mux2_1 _5727_ (.A0(net120),
    .A1(_2538_),
    .S(_2579_),
    .X(_2588_));
 sky130_fd_sc_hd__clkbuf_1 _5728_ (.A(_2588_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_1 _5729_ (.A0(net121),
    .A1(_2562_),
    .S(_2579_),
    .X(_2589_));
 sky130_fd_sc_hd__clkbuf_1 _5730_ (.A(_2589_),
    .X(_0260_));
 sky130_fd_sc_hd__buf_4 _5731_ (.A(_1800_),
    .X(_2590_));
 sky130_fd_sc_hd__mux2_1 _5732_ (.A0(\core_1.ew_reg_ie[0] ),
    .A1(\core_1.dec_rf_ie[0] ),
    .S(_2590_),
    .X(_2591_));
 sky130_fd_sc_hd__clkbuf_1 _5733_ (.A(_2591_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_1 _5734_ (.A0(\core_1.ew_reg_ie[1] ),
    .A1(\core_1.dec_rf_ie[1] ),
    .S(_2590_),
    .X(_2592_));
 sky130_fd_sc_hd__clkbuf_1 _5735_ (.A(_2592_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_1 _5736_ (.A0(\core_1.ew_reg_ie[2] ),
    .A1(\core_1.dec_rf_ie[2] ),
    .S(_2590_),
    .X(_2593_));
 sky130_fd_sc_hd__clkbuf_1 _5737_ (.A(_2593_),
    .X(_0263_));
 sky130_fd_sc_hd__mux2_1 _5738_ (.A0(\core_1.ew_reg_ie[3] ),
    .A1(\core_1.dec_rf_ie[3] ),
    .S(_2590_),
    .X(_2594_));
 sky130_fd_sc_hd__clkbuf_1 _5739_ (.A(_2594_),
    .X(_0264_));
 sky130_fd_sc_hd__mux2_1 _5740_ (.A0(\core_1.ew_reg_ie[4] ),
    .A1(\core_1.dec_rf_ie[4] ),
    .S(_2590_),
    .X(_2595_));
 sky130_fd_sc_hd__clkbuf_1 _5741_ (.A(_2595_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_1 _5742_ (.A0(\core_1.ew_reg_ie[5] ),
    .A1(\core_1.dec_rf_ie[5] ),
    .S(_2590_),
    .X(_2596_));
 sky130_fd_sc_hd__clkbuf_1 _5743_ (.A(_2596_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_1 _5744_ (.A0(\core_1.ew_reg_ie[6] ),
    .A1(\core_1.dec_rf_ie[6] ),
    .S(_2590_),
    .X(_2597_));
 sky130_fd_sc_hd__clkbuf_1 _5745_ (.A(_2597_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_1 _5746_ (.A0(\core_1.ew_reg_ie[7] ),
    .A1(\core_1.dec_rf_ie[7] ),
    .S(_2590_),
    .X(_2598_));
 sky130_fd_sc_hd__clkbuf_1 _5747_ (.A(_2598_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_1 _5748_ (.A0(_1300_),
    .A1(\core_1.dec_mem_access ),
    .S(_2590_),
    .X(_2599_));
 sky130_fd_sc_hd__clkbuf_1 _5749_ (.A(_2599_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_1 _5750_ (.A0(\core_1.ew_mem_width ),
    .A1(\core_1.dec_mem_width ),
    .S(_2590_),
    .X(_2600_));
 sky130_fd_sc_hd__clkbuf_1 _5751_ (.A(_2600_),
    .X(_0270_));
 sky130_fd_sc_hd__mux2_1 _5752_ (.A0(net155),
    .A1(_0707_),
    .S(_1800_),
    .X(_2601_));
 sky130_fd_sc_hd__clkbuf_1 _5753_ (.A(_2601_),
    .X(_0271_));
 sky130_fd_sc_hd__nor2_1 _5754_ (.A(_1165_),
    .B(_0735_),
    .Y(_0272_));
 sky130_fd_sc_hd__mux2_4 _5755_ (.A0(\core_1.ew_submit ),
    .A1(net20),
    .S(\core_1.ew_mem_access ),
    .X(_2602_));
 sky130_fd_sc_hd__buf_6 _5756_ (.A(_2602_),
    .X(_2603_));
 sky130_fd_sc_hd__nand2_4 _5757_ (.A(\core_1.ew_reg_ie[7] ),
    .B(_2603_),
    .Y(_2604_));
 sky130_fd_sc_hd__mux2_1 _5758_ (.A0(net35),
    .A1(net21),
    .S(_0983_),
    .X(_2605_));
 sky130_fd_sc_hd__mux2_1 _5759_ (.A0(\core_1.ew_data[0] ),
    .A1(_2605_),
    .S(_1299_),
    .X(_2606_));
 sky130_fd_sc_hd__clkbuf_8 _5760_ (.A(_2606_),
    .X(_2607_));
 sky130_fd_sc_hd__and2_2 _5761_ (.A(\core_1.ew_reg_ie[7] ),
    .B(_2602_),
    .X(_2608_));
 sky130_fd_sc_hd__clkbuf_4 _5762_ (.A(_2608_),
    .X(_2609_));
 sky130_fd_sc_hd__or2_1 _5763_ (.A(\core_1.execute.rf.reg_outputs[7][0] ),
    .B(_2609_),
    .X(_2610_));
 sky130_fd_sc_hd__o211a_1 _5764_ (.A1(_2604_),
    .A2(_2607_),
    .B1(_2610_),
    .C1(_1789_),
    .X(_0273_));
 sky130_fd_sc_hd__mux2_1 _5765_ (.A0(net36),
    .A1(net28),
    .S(_0983_),
    .X(_2611_));
 sky130_fd_sc_hd__mux2_1 _5766_ (.A0(\core_1.ew_data[1] ),
    .A1(_2611_),
    .S(_1299_),
    .X(_2612_));
 sky130_fd_sc_hd__clkbuf_8 _5767_ (.A(_2612_),
    .X(_2613_));
 sky130_fd_sc_hd__or2_1 _5768_ (.A(\core_1.execute.rf.reg_outputs[7][1] ),
    .B(_2609_),
    .X(_2614_));
 sky130_fd_sc_hd__o211a_1 _5769_ (.A1(_2604_),
    .A2(_2613_),
    .B1(_2614_),
    .C1(_1789_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_1 _5770_ (.A0(net22),
    .A1(net29),
    .S(_0982_),
    .X(_2615_));
 sky130_fd_sc_hd__mux2_1 _5771_ (.A0(\core_1.ew_data[2] ),
    .A1(_2615_),
    .S(_1299_),
    .X(_2616_));
 sky130_fd_sc_hd__buf_4 _5772_ (.A(_2616_),
    .X(_2617_));
 sky130_fd_sc_hd__or2_1 _5773_ (.A(\core_1.execute.rf.reg_outputs[7][2] ),
    .B(_2609_),
    .X(_2618_));
 sky130_fd_sc_hd__o211a_1 _5774_ (.A1(_2604_),
    .A2(_2617_),
    .B1(_2618_),
    .C1(_1789_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_1 _5775_ (.A0(net23),
    .A1(net30),
    .S(_0982_),
    .X(_2619_));
 sky130_fd_sc_hd__mux2_1 _5776_ (.A0(\core_1.ew_data[3] ),
    .A1(_2619_),
    .S(_1299_),
    .X(_2620_));
 sky130_fd_sc_hd__buf_6 _5777_ (.A(_2620_),
    .X(_2621_));
 sky130_fd_sc_hd__or2_1 _5778_ (.A(\core_1.execute.rf.reg_outputs[7][3] ),
    .B(_2609_),
    .X(_2622_));
 sky130_fd_sc_hd__clkbuf_4 _5779_ (.A(_1788_),
    .X(_2623_));
 sky130_fd_sc_hd__o211a_1 _5780_ (.A1(_2604_),
    .A2(_2621_),
    .B1(_2622_),
    .C1(_2623_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_1 _5781_ (.A0(net24),
    .A1(net31),
    .S(_0982_),
    .X(_2624_));
 sky130_fd_sc_hd__mux2_1 _5782_ (.A0(\core_1.ew_data[4] ),
    .A1(_2624_),
    .S(_1299_),
    .X(_2625_));
 sky130_fd_sc_hd__buf_6 _5783_ (.A(_2625_),
    .X(_2626_));
 sky130_fd_sc_hd__or2_1 _5784_ (.A(\core_1.execute.rf.reg_outputs[7][4] ),
    .B(_2608_),
    .X(_2627_));
 sky130_fd_sc_hd__o211a_1 _5785_ (.A1(_2604_),
    .A2(_2626_),
    .B1(_2627_),
    .C1(_2623_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_1 _5786_ (.A0(net25),
    .A1(net32),
    .S(_0982_),
    .X(_2628_));
 sky130_fd_sc_hd__mux2_1 _5787_ (.A0(\core_1.ew_data[5] ),
    .A1(_2628_),
    .S(_1299_),
    .X(_2629_));
 sky130_fd_sc_hd__buf_4 _5788_ (.A(_2629_),
    .X(_2630_));
 sky130_fd_sc_hd__or2_1 _5789_ (.A(\core_1.execute.rf.reg_outputs[7][5] ),
    .B(_2608_),
    .X(_2631_));
 sky130_fd_sc_hd__o211a_1 _5790_ (.A1(_2604_),
    .A2(_2630_),
    .B1(_2631_),
    .C1(_2623_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_1 _5791_ (.A0(net26),
    .A1(net33),
    .S(_0982_),
    .X(_2632_));
 sky130_fd_sc_hd__mux2_1 _5792_ (.A0(\core_1.ew_data[6] ),
    .A1(_2632_),
    .S(_1299_),
    .X(_2633_));
 sky130_fd_sc_hd__buf_4 _5793_ (.A(_2633_),
    .X(_2634_));
 sky130_fd_sc_hd__or2_1 _5794_ (.A(\core_1.execute.rf.reg_outputs[7][6] ),
    .B(_2608_),
    .X(_2635_));
 sky130_fd_sc_hd__o211a_1 _5795_ (.A1(_2604_),
    .A2(_2634_),
    .B1(_2635_),
    .C1(_2623_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_1 _5796_ (.A0(net27),
    .A1(net34),
    .S(_0982_),
    .X(_2636_));
 sky130_fd_sc_hd__mux2_1 _5797_ (.A0(\core_1.ew_data[7] ),
    .A1(_2636_),
    .S(_1299_),
    .X(_2637_));
 sky130_fd_sc_hd__buf_4 _5798_ (.A(_2637_),
    .X(_2638_));
 sky130_fd_sc_hd__or2_1 _5799_ (.A(\core_1.execute.rf.reg_outputs[7][7] ),
    .B(_2608_),
    .X(_2639_));
 sky130_fd_sc_hd__o211a_1 _5800_ (.A1(_2604_),
    .A2(_2638_),
    .B1(_2639_),
    .C1(_2623_),
    .X(_0280_));
 sky130_fd_sc_hd__buf_2 _5801_ (.A(_2608_),
    .X(_2640_));
 sky130_fd_sc_hd__and2b_1 _5802_ (.A_N(\core_1.ew_mem_width ),
    .B(_1299_),
    .X(_2641_));
 sky130_fd_sc_hd__buf_4 _5803_ (.A(_2641_),
    .X(_2642_));
 sky130_fd_sc_hd__inv_2 _5804_ (.A(\core_1.ew_data[8] ),
    .Y(_2643_));
 sky130_fd_sc_hd__o2bb2a_4 _5805_ (.A1_N(net35),
    .A2_N(_2642_),
    .B1(_2643_),
    .B2(_1300_),
    .X(_2644_));
 sky130_fd_sc_hd__nand2_1 _5806_ (.A(_2640_),
    .B(_2644_),
    .Y(_2645_));
 sky130_fd_sc_hd__o211a_1 _5807_ (.A1(\core_1.execute.rf.reg_outputs[7][8] ),
    .A2(_2640_),
    .B1(_2645_),
    .C1(_2623_),
    .X(_0281_));
 sky130_fd_sc_hd__o2bb2a_4 _5808_ (.A1_N(net36),
    .A2_N(_2642_),
    .B1(_2357_),
    .B2(_1300_),
    .X(_2646_));
 sky130_fd_sc_hd__nand2_1 _5809_ (.A(_2640_),
    .B(_2646_),
    .Y(_2647_));
 sky130_fd_sc_hd__o211a_1 _5810_ (.A1(\core_1.execute.rf.reg_outputs[7][9] ),
    .A2(_2640_),
    .B1(_2647_),
    .C1(_2623_),
    .X(_0282_));
 sky130_fd_sc_hd__inv_2 _5811_ (.A(\core_1.ew_data[10] ),
    .Y(_2648_));
 sky130_fd_sc_hd__o2bb2a_4 _5812_ (.A1_N(net22),
    .A2_N(_2642_),
    .B1(_2648_),
    .B2(_1300_),
    .X(_2649_));
 sky130_fd_sc_hd__nand2_1 _5813_ (.A(_2609_),
    .B(_2649_),
    .Y(_2650_));
 sky130_fd_sc_hd__o211a_1 _5814_ (.A1(\core_1.execute.rf.reg_outputs[7][10] ),
    .A2(_2640_),
    .B1(_2650_),
    .C1(_2623_),
    .X(_0283_));
 sky130_fd_sc_hd__inv_2 _5815_ (.A(\core_1.ew_data[11] ),
    .Y(_2651_));
 sky130_fd_sc_hd__o2bb2a_4 _5816_ (.A1_N(net23),
    .A2_N(_2642_),
    .B1(_2651_),
    .B2(_1300_),
    .X(_2652_));
 sky130_fd_sc_hd__nand2_1 _5817_ (.A(_2609_),
    .B(_2652_),
    .Y(_2653_));
 sky130_fd_sc_hd__o211a_1 _5818_ (.A1(\core_1.execute.rf.reg_outputs[7][11] ),
    .A2(_2640_),
    .B1(_2653_),
    .C1(_2623_),
    .X(_0284_));
 sky130_fd_sc_hd__inv_2 _5819_ (.A(\core_1.ew_data[12] ),
    .Y(_2654_));
 sky130_fd_sc_hd__o2bb2a_4 _5820_ (.A1_N(net24),
    .A2_N(_2642_),
    .B1(_2654_),
    .B2(_1300_),
    .X(_2655_));
 sky130_fd_sc_hd__nand2_1 _5821_ (.A(_2609_),
    .B(_2655_),
    .Y(_2656_));
 sky130_fd_sc_hd__o211a_1 _5822_ (.A1(\core_1.execute.rf.reg_outputs[7][12] ),
    .A2(_2640_),
    .B1(_2656_),
    .C1(_2623_),
    .X(_0285_));
 sky130_fd_sc_hd__inv_2 _5823_ (.A(\core_1.ew_data[13] ),
    .Y(_2657_));
 sky130_fd_sc_hd__o2bb2a_4 _5824_ (.A1_N(net25),
    .A2_N(_2642_),
    .B1(_2657_),
    .B2(_1300_),
    .X(_2658_));
 sky130_fd_sc_hd__nand2_1 _5825_ (.A(_2609_),
    .B(_2658_),
    .Y(_2659_));
 sky130_fd_sc_hd__clkbuf_4 _5826_ (.A(_1788_),
    .X(_2660_));
 sky130_fd_sc_hd__o211a_1 _5827_ (.A1(\core_1.execute.rf.reg_outputs[7][13] ),
    .A2(_2640_),
    .B1(_2659_),
    .C1(_2660_),
    .X(_0286_));
 sky130_fd_sc_hd__inv_2 _5828_ (.A(\core_1.ew_data[14] ),
    .Y(_2661_));
 sky130_fd_sc_hd__o2bb2a_4 _5829_ (.A1_N(net26),
    .A2_N(_2642_),
    .B1(_2661_),
    .B2(_1300_),
    .X(_2662_));
 sky130_fd_sc_hd__nand2_1 _5830_ (.A(_2609_),
    .B(_2662_),
    .Y(_2663_));
 sky130_fd_sc_hd__o211a_1 _5831_ (.A1(\core_1.execute.rf.reg_outputs[7][14] ),
    .A2(_2640_),
    .B1(_2663_),
    .C1(_2660_),
    .X(_0287_));
 sky130_fd_sc_hd__inv_2 _5832_ (.A(\core_1.ew_data[15] ),
    .Y(_2664_));
 sky130_fd_sc_hd__o2bb2a_4 _5833_ (.A1_N(net27),
    .A2_N(_2642_),
    .B1(_2664_),
    .B2(_1300_),
    .X(_2665_));
 sky130_fd_sc_hd__nand2_1 _5834_ (.A(_2609_),
    .B(_2665_),
    .Y(_2666_));
 sky130_fd_sc_hd__o211a_1 _5835_ (.A1(\core_1.execute.rf.reg_outputs[7][15] ),
    .A2(_2640_),
    .B1(_2666_),
    .C1(_2660_),
    .X(_0288_));
 sky130_fd_sc_hd__nand2_2 _5836_ (.A(\core_1.ew_reg_ie[6] ),
    .B(_2603_),
    .Y(_2667_));
 sky130_fd_sc_hd__and2_1 _5837_ (.A(\core_1.ew_reg_ie[6] ),
    .B(_2603_),
    .X(_2668_));
 sky130_fd_sc_hd__buf_2 _5838_ (.A(_2668_),
    .X(_2669_));
 sky130_fd_sc_hd__or2_1 _5839_ (.A(\core_1.execute.rf.reg_outputs[6][0] ),
    .B(_2669_),
    .X(_2670_));
 sky130_fd_sc_hd__o211a_1 _5840_ (.A1(_2607_),
    .A2(_2667_),
    .B1(_2670_),
    .C1(_2660_),
    .X(_0289_));
 sky130_fd_sc_hd__or2_1 _5841_ (.A(\core_1.execute.rf.reg_outputs[6][1] ),
    .B(_2669_),
    .X(_2671_));
 sky130_fd_sc_hd__o211a_1 _5842_ (.A1(_2613_),
    .A2(_2667_),
    .B1(_2671_),
    .C1(_2660_),
    .X(_0290_));
 sky130_fd_sc_hd__or2_1 _5843_ (.A(\core_1.execute.rf.reg_outputs[6][2] ),
    .B(_2669_),
    .X(_2672_));
 sky130_fd_sc_hd__o211a_1 _5844_ (.A1(_2617_),
    .A2(_2667_),
    .B1(_2672_),
    .C1(_2660_),
    .X(_0291_));
 sky130_fd_sc_hd__or2_1 _5845_ (.A(\core_1.execute.rf.reg_outputs[6][3] ),
    .B(_2669_),
    .X(_2673_));
 sky130_fd_sc_hd__o211a_1 _5846_ (.A1(_2621_),
    .A2(_2667_),
    .B1(_2673_),
    .C1(_2660_),
    .X(_0292_));
 sky130_fd_sc_hd__or2_1 _5847_ (.A(\core_1.execute.rf.reg_outputs[6][4] ),
    .B(_2668_),
    .X(_2674_));
 sky130_fd_sc_hd__o211a_1 _5848_ (.A1(_2626_),
    .A2(_2667_),
    .B1(_2674_),
    .C1(_2660_),
    .X(_0293_));
 sky130_fd_sc_hd__or2_1 _5849_ (.A(\core_1.execute.rf.reg_outputs[6][5] ),
    .B(_2668_),
    .X(_2675_));
 sky130_fd_sc_hd__o211a_1 _5850_ (.A1(_2630_),
    .A2(_2667_),
    .B1(_2675_),
    .C1(_2660_),
    .X(_0294_));
 sky130_fd_sc_hd__or2_1 _5851_ (.A(\core_1.execute.rf.reg_outputs[6][6] ),
    .B(_2668_),
    .X(_2676_));
 sky130_fd_sc_hd__o211a_1 _5852_ (.A1(_2634_),
    .A2(_2667_),
    .B1(_2676_),
    .C1(_2660_),
    .X(_0295_));
 sky130_fd_sc_hd__or2_1 _5853_ (.A(\core_1.execute.rf.reg_outputs[6][7] ),
    .B(_2668_),
    .X(_2677_));
 sky130_fd_sc_hd__clkbuf_4 _5854_ (.A(_1788_),
    .X(_2678_));
 sky130_fd_sc_hd__o211a_1 _5855_ (.A1(_2638_),
    .A2(_2667_),
    .B1(_2677_),
    .C1(_2678_),
    .X(_0296_));
 sky130_fd_sc_hd__clkbuf_4 _5856_ (.A(_2668_),
    .X(_2679_));
 sky130_fd_sc_hd__nand2_1 _5857_ (.A(_2644_),
    .B(_2679_),
    .Y(_2680_));
 sky130_fd_sc_hd__o211a_1 _5858_ (.A1(\core_1.execute.rf.reg_outputs[6][8] ),
    .A2(_2679_),
    .B1(_2680_),
    .C1(_2678_),
    .X(_0297_));
 sky130_fd_sc_hd__nand2_1 _5859_ (.A(_2646_),
    .B(_2679_),
    .Y(_2681_));
 sky130_fd_sc_hd__o211a_1 _5860_ (.A1(\core_1.execute.rf.reg_outputs[6][9] ),
    .A2(_2679_),
    .B1(_2681_),
    .C1(_2678_),
    .X(_0298_));
 sky130_fd_sc_hd__nand2_1 _5861_ (.A(_2649_),
    .B(_2669_),
    .Y(_2682_));
 sky130_fd_sc_hd__o211a_1 _5862_ (.A1(\core_1.execute.rf.reg_outputs[6][10] ),
    .A2(_2679_),
    .B1(_2682_),
    .C1(_2678_),
    .X(_0299_));
 sky130_fd_sc_hd__nand2_1 _5863_ (.A(_2652_),
    .B(_2669_),
    .Y(_2683_));
 sky130_fd_sc_hd__o211a_1 _5864_ (.A1(\core_1.execute.rf.reg_outputs[6][11] ),
    .A2(_2679_),
    .B1(_2683_),
    .C1(_2678_),
    .X(_0300_));
 sky130_fd_sc_hd__nand2_1 _5865_ (.A(_2655_),
    .B(_2669_),
    .Y(_2684_));
 sky130_fd_sc_hd__o211a_1 _5866_ (.A1(\core_1.execute.rf.reg_outputs[6][12] ),
    .A2(_2679_),
    .B1(_2684_),
    .C1(_2678_),
    .X(_0301_));
 sky130_fd_sc_hd__nand2_1 _5867_ (.A(_2658_),
    .B(_2669_),
    .Y(_2685_));
 sky130_fd_sc_hd__o211a_1 _5868_ (.A1(\core_1.execute.rf.reg_outputs[6][13] ),
    .A2(_2679_),
    .B1(_2685_),
    .C1(_2678_),
    .X(_0302_));
 sky130_fd_sc_hd__nand2_1 _5869_ (.A(_2662_),
    .B(_2669_),
    .Y(_2686_));
 sky130_fd_sc_hd__o211a_1 _5870_ (.A1(\core_1.execute.rf.reg_outputs[6][14] ),
    .A2(_2679_),
    .B1(_2686_),
    .C1(_2678_),
    .X(_0303_));
 sky130_fd_sc_hd__nand2_1 _5871_ (.A(_2665_),
    .B(_2669_),
    .Y(_2687_));
 sky130_fd_sc_hd__o211a_1 _5872_ (.A1(\core_1.execute.rf.reg_outputs[6][15] ),
    .A2(_2679_),
    .B1(_2687_),
    .C1(_2678_),
    .X(_0304_));
 sky130_fd_sc_hd__nand2_2 _5873_ (.A(\core_1.ew_reg_ie[5] ),
    .B(_2603_),
    .Y(_2688_));
 sky130_fd_sc_hd__and2_1 _5874_ (.A(\core_1.ew_reg_ie[5] ),
    .B(_2603_),
    .X(_2689_));
 sky130_fd_sc_hd__clkbuf_4 _5875_ (.A(_2689_),
    .X(_2690_));
 sky130_fd_sc_hd__or2_1 _5876_ (.A(\core_1.execute.rf.reg_outputs[5][0] ),
    .B(_2690_),
    .X(_2691_));
 sky130_fd_sc_hd__o211a_1 _5877_ (.A1(_2607_),
    .A2(_2688_),
    .B1(_2691_),
    .C1(_2678_),
    .X(_0305_));
 sky130_fd_sc_hd__or2_1 _5878_ (.A(\core_1.execute.rf.reg_outputs[5][1] ),
    .B(_2690_),
    .X(_2692_));
 sky130_fd_sc_hd__clkbuf_4 _5879_ (.A(_1788_),
    .X(_2693_));
 sky130_fd_sc_hd__o211a_1 _5880_ (.A1(_2613_),
    .A2(_2688_),
    .B1(_2692_),
    .C1(_2693_),
    .X(_0306_));
 sky130_fd_sc_hd__or2_1 _5881_ (.A(\core_1.execute.rf.reg_outputs[5][2] ),
    .B(_2690_),
    .X(_2694_));
 sky130_fd_sc_hd__o211a_1 _5882_ (.A1(_2617_),
    .A2(_2688_),
    .B1(_2694_),
    .C1(_2693_),
    .X(_0307_));
 sky130_fd_sc_hd__or2_1 _5883_ (.A(\core_1.execute.rf.reg_outputs[5][3] ),
    .B(_2690_),
    .X(_2695_));
 sky130_fd_sc_hd__o211a_1 _5884_ (.A1(_2621_),
    .A2(_2688_),
    .B1(_2695_),
    .C1(_2693_),
    .X(_0308_));
 sky130_fd_sc_hd__or2_1 _5885_ (.A(\core_1.execute.rf.reg_outputs[5][4] ),
    .B(_2689_),
    .X(_2696_));
 sky130_fd_sc_hd__o211a_1 _5886_ (.A1(_2626_),
    .A2(_2688_),
    .B1(_2696_),
    .C1(_2693_),
    .X(_0309_));
 sky130_fd_sc_hd__or2_1 _5887_ (.A(\core_1.execute.rf.reg_outputs[5][5] ),
    .B(_2689_),
    .X(_2697_));
 sky130_fd_sc_hd__o211a_1 _5888_ (.A1(_2630_),
    .A2(_2688_),
    .B1(_2697_),
    .C1(_2693_),
    .X(_0310_));
 sky130_fd_sc_hd__or2_1 _5889_ (.A(\core_1.execute.rf.reg_outputs[5][6] ),
    .B(_2689_),
    .X(_2698_));
 sky130_fd_sc_hd__o211a_1 _5890_ (.A1(_2634_),
    .A2(_2688_),
    .B1(_2698_),
    .C1(_2693_),
    .X(_0311_));
 sky130_fd_sc_hd__or2_1 _5891_ (.A(\core_1.execute.rf.reg_outputs[5][7] ),
    .B(_2689_),
    .X(_2699_));
 sky130_fd_sc_hd__o211a_1 _5892_ (.A1(_2638_),
    .A2(_2688_),
    .B1(_2699_),
    .C1(_2693_),
    .X(_0312_));
 sky130_fd_sc_hd__buf_2 _5893_ (.A(_2689_),
    .X(_2700_));
 sky130_fd_sc_hd__nand2_1 _5894_ (.A(_2644_),
    .B(_2700_),
    .Y(_2701_));
 sky130_fd_sc_hd__o211a_1 _5895_ (.A1(\core_1.execute.rf.reg_outputs[5][8] ),
    .A2(_2700_),
    .B1(_2701_),
    .C1(_2693_),
    .X(_0313_));
 sky130_fd_sc_hd__nand2_1 _5896_ (.A(_2646_),
    .B(_2700_),
    .Y(_2702_));
 sky130_fd_sc_hd__o211a_1 _5897_ (.A1(\core_1.execute.rf.reg_outputs[5][9] ),
    .A2(_2700_),
    .B1(_2702_),
    .C1(_2693_),
    .X(_0314_));
 sky130_fd_sc_hd__nand2_1 _5898_ (.A(_2649_),
    .B(_2690_),
    .Y(_2703_));
 sky130_fd_sc_hd__o211a_1 _5899_ (.A1(\core_1.execute.rf.reg_outputs[5][10] ),
    .A2(_2700_),
    .B1(_2703_),
    .C1(_2693_),
    .X(_0315_));
 sky130_fd_sc_hd__nand2_1 _5900_ (.A(_2652_),
    .B(_2690_),
    .Y(_2704_));
 sky130_fd_sc_hd__clkbuf_4 _5901_ (.A(_1788_),
    .X(_2705_));
 sky130_fd_sc_hd__o211a_1 _5902_ (.A1(\core_1.execute.rf.reg_outputs[5][11] ),
    .A2(_2700_),
    .B1(_2704_),
    .C1(_2705_),
    .X(_0316_));
 sky130_fd_sc_hd__nand2_1 _5903_ (.A(_2655_),
    .B(_2690_),
    .Y(_2706_));
 sky130_fd_sc_hd__o211a_1 _5904_ (.A1(\core_1.execute.rf.reg_outputs[5][12] ),
    .A2(_2700_),
    .B1(_2706_),
    .C1(_2705_),
    .X(_0317_));
 sky130_fd_sc_hd__nand2_1 _5905_ (.A(_2658_),
    .B(_2690_),
    .Y(_2707_));
 sky130_fd_sc_hd__o211a_1 _5906_ (.A1(\core_1.execute.rf.reg_outputs[5][13] ),
    .A2(_2700_),
    .B1(_2707_),
    .C1(_2705_),
    .X(_0318_));
 sky130_fd_sc_hd__nand2_1 _5907_ (.A(_2662_),
    .B(_2690_),
    .Y(_2708_));
 sky130_fd_sc_hd__o211a_1 _5908_ (.A1(\core_1.execute.rf.reg_outputs[5][14] ),
    .A2(_2700_),
    .B1(_2708_),
    .C1(_2705_),
    .X(_0319_));
 sky130_fd_sc_hd__nand2_1 _5909_ (.A(_2665_),
    .B(_2690_),
    .Y(_2709_));
 sky130_fd_sc_hd__o211a_1 _5910_ (.A1(\core_1.execute.rf.reg_outputs[5][15] ),
    .A2(_2700_),
    .B1(_2709_),
    .C1(_2705_),
    .X(_0320_));
 sky130_fd_sc_hd__nand2_4 _5911_ (.A(\core_1.ew_reg_ie[4] ),
    .B(_2603_),
    .Y(_2710_));
 sky130_fd_sc_hd__and2_1 _5912_ (.A(\core_1.ew_reg_ie[4] ),
    .B(_2602_),
    .X(_2711_));
 sky130_fd_sc_hd__clkbuf_4 _5913_ (.A(_2711_),
    .X(_2712_));
 sky130_fd_sc_hd__or2_1 _5914_ (.A(\core_1.execute.rf.reg_outputs[4][0] ),
    .B(_2712_),
    .X(_2713_));
 sky130_fd_sc_hd__o211a_1 _5915_ (.A1(_2607_),
    .A2(_2710_),
    .B1(_2713_),
    .C1(_2705_),
    .X(_0321_));
 sky130_fd_sc_hd__or2_1 _5916_ (.A(\core_1.execute.rf.reg_outputs[4][1] ),
    .B(_2712_),
    .X(_2714_));
 sky130_fd_sc_hd__o211a_1 _5917_ (.A1(_2613_),
    .A2(_2710_),
    .B1(_2714_),
    .C1(_2705_),
    .X(_0322_));
 sky130_fd_sc_hd__or2_1 _5918_ (.A(\core_1.execute.rf.reg_outputs[4][2] ),
    .B(_2712_),
    .X(_2715_));
 sky130_fd_sc_hd__o211a_1 _5919_ (.A1(_2617_),
    .A2(_2710_),
    .B1(_2715_),
    .C1(_2705_),
    .X(_0323_));
 sky130_fd_sc_hd__or2_1 _5920_ (.A(\core_1.execute.rf.reg_outputs[4][3] ),
    .B(_2712_),
    .X(_2716_));
 sky130_fd_sc_hd__o211a_1 _5921_ (.A1(_2621_),
    .A2(_2710_),
    .B1(_2716_),
    .C1(_2705_),
    .X(_0324_));
 sky130_fd_sc_hd__or2_1 _5922_ (.A(\core_1.execute.rf.reg_outputs[4][4] ),
    .B(_2711_),
    .X(_2717_));
 sky130_fd_sc_hd__o211a_1 _5923_ (.A1(_2626_),
    .A2(_2710_),
    .B1(_2717_),
    .C1(_2705_),
    .X(_0325_));
 sky130_fd_sc_hd__or2_1 _5924_ (.A(\core_1.execute.rf.reg_outputs[4][5] ),
    .B(_2711_),
    .X(_2718_));
 sky130_fd_sc_hd__clkbuf_4 _5925_ (.A(_1788_),
    .X(_2719_));
 sky130_fd_sc_hd__o211a_1 _5926_ (.A1(_2630_),
    .A2(_2710_),
    .B1(_2718_),
    .C1(_2719_),
    .X(_0326_));
 sky130_fd_sc_hd__or2_1 _5927_ (.A(\core_1.execute.rf.reg_outputs[4][6] ),
    .B(_2711_),
    .X(_2720_));
 sky130_fd_sc_hd__o211a_1 _5928_ (.A1(_2634_),
    .A2(_2710_),
    .B1(_2720_),
    .C1(_2719_),
    .X(_0327_));
 sky130_fd_sc_hd__or2_1 _5929_ (.A(\core_1.execute.rf.reg_outputs[4][7] ),
    .B(_2711_),
    .X(_2721_));
 sky130_fd_sc_hd__o211a_1 _5930_ (.A1(_2638_),
    .A2(_2710_),
    .B1(_2721_),
    .C1(_2719_),
    .X(_0328_));
 sky130_fd_sc_hd__clkbuf_4 _5931_ (.A(_2711_),
    .X(_2722_));
 sky130_fd_sc_hd__nand2_1 _5932_ (.A(_2644_),
    .B(_2722_),
    .Y(_2723_));
 sky130_fd_sc_hd__o211a_1 _5933_ (.A1(\core_1.execute.rf.reg_outputs[4][8] ),
    .A2(_2722_),
    .B1(_2723_),
    .C1(_2719_),
    .X(_0329_));
 sky130_fd_sc_hd__nand2_1 _5934_ (.A(_2646_),
    .B(_2722_),
    .Y(_2724_));
 sky130_fd_sc_hd__o211a_1 _5935_ (.A1(\core_1.execute.rf.reg_outputs[4][9] ),
    .A2(_2722_),
    .B1(_2724_),
    .C1(_2719_),
    .X(_0330_));
 sky130_fd_sc_hd__nand2_1 _5936_ (.A(_2649_),
    .B(_2712_),
    .Y(_2725_));
 sky130_fd_sc_hd__o211a_1 _5937_ (.A1(\core_1.execute.rf.reg_outputs[4][10] ),
    .A2(_2722_),
    .B1(_2725_),
    .C1(_2719_),
    .X(_0331_));
 sky130_fd_sc_hd__nand2_1 _5938_ (.A(_2652_),
    .B(_2712_),
    .Y(_2726_));
 sky130_fd_sc_hd__o211a_1 _5939_ (.A1(\core_1.execute.rf.reg_outputs[4][11] ),
    .A2(_2722_),
    .B1(_2726_),
    .C1(_2719_),
    .X(_0332_));
 sky130_fd_sc_hd__nand2_1 _5940_ (.A(_2655_),
    .B(_2712_),
    .Y(_2727_));
 sky130_fd_sc_hd__o211a_1 _5941_ (.A1(\core_1.execute.rf.reg_outputs[4][12] ),
    .A2(_2722_),
    .B1(_2727_),
    .C1(_2719_),
    .X(_0333_));
 sky130_fd_sc_hd__nand2_1 _5942_ (.A(_2658_),
    .B(_2712_),
    .Y(_2728_));
 sky130_fd_sc_hd__o211a_1 _5943_ (.A1(\core_1.execute.rf.reg_outputs[4][13] ),
    .A2(_2722_),
    .B1(_2728_),
    .C1(_2719_),
    .X(_0334_));
 sky130_fd_sc_hd__nand2_1 _5944_ (.A(_2662_),
    .B(_2712_),
    .Y(_2729_));
 sky130_fd_sc_hd__o211a_1 _5945_ (.A1(\core_1.execute.rf.reg_outputs[4][14] ),
    .A2(_2722_),
    .B1(_2729_),
    .C1(_2719_),
    .X(_0335_));
 sky130_fd_sc_hd__nand2_1 _5946_ (.A(_2665_),
    .B(_2712_),
    .Y(_2730_));
 sky130_fd_sc_hd__buf_4 _5947_ (.A(_1788_),
    .X(_2731_));
 sky130_fd_sc_hd__o211a_1 _5948_ (.A1(\core_1.execute.rf.reg_outputs[4][15] ),
    .A2(_2722_),
    .B1(_2730_),
    .C1(_2731_),
    .X(_0336_));
 sky130_fd_sc_hd__nand2_4 _5949_ (.A(\core_1.ew_reg_ie[3] ),
    .B(_2603_),
    .Y(_2732_));
 sky130_fd_sc_hd__and2_2 _5950_ (.A(\core_1.ew_reg_ie[3] ),
    .B(_2602_),
    .X(_2733_));
 sky130_fd_sc_hd__buf_4 _5951_ (.A(_2733_),
    .X(_2734_));
 sky130_fd_sc_hd__or2_1 _5952_ (.A(\core_1.execute.rf.reg_outputs[3][0] ),
    .B(_2734_),
    .X(_2735_));
 sky130_fd_sc_hd__o211a_1 _5953_ (.A1(_2607_),
    .A2(_2732_),
    .B1(_2735_),
    .C1(_2731_),
    .X(_0337_));
 sky130_fd_sc_hd__or2_1 _5954_ (.A(\core_1.execute.rf.reg_outputs[3][1] ),
    .B(_2734_),
    .X(_2736_));
 sky130_fd_sc_hd__o211a_1 _5955_ (.A1(_2613_),
    .A2(_2732_),
    .B1(_2736_),
    .C1(_2731_),
    .X(_0338_));
 sky130_fd_sc_hd__or2_1 _5956_ (.A(\core_1.execute.rf.reg_outputs[3][2] ),
    .B(_2734_),
    .X(_2737_));
 sky130_fd_sc_hd__o211a_1 _5957_ (.A1(_2617_),
    .A2(_2732_),
    .B1(_2737_),
    .C1(_2731_),
    .X(_0339_));
 sky130_fd_sc_hd__or2_1 _5958_ (.A(\core_1.execute.rf.reg_outputs[3][3] ),
    .B(_2734_),
    .X(_2738_));
 sky130_fd_sc_hd__o211a_1 _5959_ (.A1(_2621_),
    .A2(_2732_),
    .B1(_2738_),
    .C1(_2731_),
    .X(_0340_));
 sky130_fd_sc_hd__or2_1 _5960_ (.A(\core_1.execute.rf.reg_outputs[3][4] ),
    .B(_2733_),
    .X(_2739_));
 sky130_fd_sc_hd__o211a_1 _5961_ (.A1(_2626_),
    .A2(_2732_),
    .B1(_2739_),
    .C1(_2731_),
    .X(_0341_));
 sky130_fd_sc_hd__or2_1 _5962_ (.A(\core_1.execute.rf.reg_outputs[3][5] ),
    .B(_2733_),
    .X(_2740_));
 sky130_fd_sc_hd__o211a_1 _5963_ (.A1(_2630_),
    .A2(_2732_),
    .B1(_2740_),
    .C1(_2731_),
    .X(_0342_));
 sky130_fd_sc_hd__or2_1 _5964_ (.A(\core_1.execute.rf.reg_outputs[3][6] ),
    .B(_2733_),
    .X(_2741_));
 sky130_fd_sc_hd__o211a_1 _5965_ (.A1(_2634_),
    .A2(_2732_),
    .B1(_2741_),
    .C1(_2731_),
    .X(_0343_));
 sky130_fd_sc_hd__or2_1 _5966_ (.A(\core_1.execute.rf.reg_outputs[3][7] ),
    .B(_2733_),
    .X(_2742_));
 sky130_fd_sc_hd__o211a_1 _5967_ (.A1(_2638_),
    .A2(_2732_),
    .B1(_2742_),
    .C1(_2731_),
    .X(_0344_));
 sky130_fd_sc_hd__clkbuf_4 _5968_ (.A(_2733_),
    .X(_2743_));
 sky130_fd_sc_hd__nand2_1 _5969_ (.A(_2644_),
    .B(_2743_),
    .Y(_2744_));
 sky130_fd_sc_hd__o211a_1 _5970_ (.A1(\core_1.execute.rf.reg_outputs[3][8] ),
    .A2(_2743_),
    .B1(_2744_),
    .C1(_2731_),
    .X(_0345_));
 sky130_fd_sc_hd__nand2_1 _5971_ (.A(_2646_),
    .B(_2743_),
    .Y(_2745_));
 sky130_fd_sc_hd__clkbuf_4 _5972_ (.A(_1788_),
    .X(_2746_));
 sky130_fd_sc_hd__o211a_1 _5973_ (.A1(\core_1.execute.rf.reg_outputs[3][9] ),
    .A2(_2743_),
    .B1(_2745_),
    .C1(_2746_),
    .X(_0346_));
 sky130_fd_sc_hd__nand2_1 _5974_ (.A(_2649_),
    .B(_2734_),
    .Y(_2747_));
 sky130_fd_sc_hd__o211a_1 _5975_ (.A1(\core_1.execute.rf.reg_outputs[3][10] ),
    .A2(_2743_),
    .B1(_2747_),
    .C1(_2746_),
    .X(_0347_));
 sky130_fd_sc_hd__nand2_1 _5976_ (.A(_2652_),
    .B(_2734_),
    .Y(_2748_));
 sky130_fd_sc_hd__o211a_1 _5977_ (.A1(\core_1.execute.rf.reg_outputs[3][11] ),
    .A2(_2743_),
    .B1(_2748_),
    .C1(_2746_),
    .X(_0348_));
 sky130_fd_sc_hd__nand2_1 _5978_ (.A(_2655_),
    .B(_2734_),
    .Y(_2749_));
 sky130_fd_sc_hd__o211a_1 _5979_ (.A1(\core_1.execute.rf.reg_outputs[3][12] ),
    .A2(_2743_),
    .B1(_2749_),
    .C1(_2746_),
    .X(_0349_));
 sky130_fd_sc_hd__nand2_1 _5980_ (.A(_2658_),
    .B(_2734_),
    .Y(_2750_));
 sky130_fd_sc_hd__o211a_1 _5981_ (.A1(\core_1.execute.rf.reg_outputs[3][13] ),
    .A2(_2743_),
    .B1(_2750_),
    .C1(_2746_),
    .X(_0350_));
 sky130_fd_sc_hd__nand2_1 _5982_ (.A(_2662_),
    .B(_2734_),
    .Y(_2751_));
 sky130_fd_sc_hd__o211a_1 _5983_ (.A1(\core_1.execute.rf.reg_outputs[3][14] ),
    .A2(_2743_),
    .B1(_2751_),
    .C1(_2746_),
    .X(_0351_));
 sky130_fd_sc_hd__nand2_1 _5984_ (.A(_2665_),
    .B(_2734_),
    .Y(_2752_));
 sky130_fd_sc_hd__o211a_1 _5985_ (.A1(\core_1.execute.rf.reg_outputs[3][15] ),
    .A2(_2743_),
    .B1(_2752_),
    .C1(_2746_),
    .X(_0352_));
 sky130_fd_sc_hd__nand2_2 _5986_ (.A(\core_1.ew_reg_ie[2] ),
    .B(_2603_),
    .Y(_2753_));
 sky130_fd_sc_hd__and2_1 _5987_ (.A(\core_1.ew_reg_ie[2] ),
    .B(_2602_),
    .X(_2754_));
 sky130_fd_sc_hd__buf_2 _5988_ (.A(_2754_),
    .X(_2755_));
 sky130_fd_sc_hd__or2_1 _5989_ (.A(\core_1.execute.rf.reg_outputs[2][0] ),
    .B(_2755_),
    .X(_2756_));
 sky130_fd_sc_hd__o211a_1 _5990_ (.A1(_2607_),
    .A2(_2753_),
    .B1(_2756_),
    .C1(_2746_),
    .X(_0353_));
 sky130_fd_sc_hd__or2_1 _5991_ (.A(\core_1.execute.rf.reg_outputs[2][1] ),
    .B(_2755_),
    .X(_2757_));
 sky130_fd_sc_hd__o211a_1 _5992_ (.A1(_2613_),
    .A2(_2753_),
    .B1(_2757_),
    .C1(_2746_),
    .X(_0354_));
 sky130_fd_sc_hd__or2_1 _5993_ (.A(\core_1.execute.rf.reg_outputs[2][2] ),
    .B(_2755_),
    .X(_2758_));
 sky130_fd_sc_hd__o211a_1 _5994_ (.A1(_2617_),
    .A2(_2753_),
    .B1(_2758_),
    .C1(_2746_),
    .X(_0355_));
 sky130_fd_sc_hd__or2_1 _5995_ (.A(\core_1.execute.rf.reg_outputs[2][3] ),
    .B(_2755_),
    .X(_2759_));
 sky130_fd_sc_hd__clkbuf_4 _5996_ (.A(_1788_),
    .X(_2760_));
 sky130_fd_sc_hd__o211a_1 _5997_ (.A1(_2621_),
    .A2(_2753_),
    .B1(_2759_),
    .C1(_2760_),
    .X(_0356_));
 sky130_fd_sc_hd__or2_1 _5998_ (.A(\core_1.execute.rf.reg_outputs[2][4] ),
    .B(_2754_),
    .X(_2761_));
 sky130_fd_sc_hd__o211a_1 _5999_ (.A1(_2626_),
    .A2(_2753_),
    .B1(_2761_),
    .C1(_2760_),
    .X(_0357_));
 sky130_fd_sc_hd__or2_1 _6000_ (.A(\core_1.execute.rf.reg_outputs[2][5] ),
    .B(_2754_),
    .X(_2762_));
 sky130_fd_sc_hd__o211a_1 _6001_ (.A1(_2630_),
    .A2(_2753_),
    .B1(_2762_),
    .C1(_2760_),
    .X(_0358_));
 sky130_fd_sc_hd__or2_1 _6002_ (.A(\core_1.execute.rf.reg_outputs[2][6] ),
    .B(_2754_),
    .X(_2763_));
 sky130_fd_sc_hd__o211a_1 _6003_ (.A1(_2634_),
    .A2(_2753_),
    .B1(_2763_),
    .C1(_2760_),
    .X(_0359_));
 sky130_fd_sc_hd__or2_1 _6004_ (.A(\core_1.execute.rf.reg_outputs[2][7] ),
    .B(_2754_),
    .X(_2764_));
 sky130_fd_sc_hd__o211a_1 _6005_ (.A1(_2638_),
    .A2(_2753_),
    .B1(_2764_),
    .C1(_2760_),
    .X(_0360_));
 sky130_fd_sc_hd__buf_2 _6006_ (.A(_2754_),
    .X(_2765_));
 sky130_fd_sc_hd__nand2_1 _6007_ (.A(_2644_),
    .B(_2765_),
    .Y(_2766_));
 sky130_fd_sc_hd__o211a_1 _6008_ (.A1(\core_1.execute.rf.reg_outputs[2][8] ),
    .A2(_2765_),
    .B1(_2766_),
    .C1(_2760_),
    .X(_0361_));
 sky130_fd_sc_hd__nand2_1 _6009_ (.A(_2646_),
    .B(_2765_),
    .Y(_2767_));
 sky130_fd_sc_hd__o211a_1 _6010_ (.A1(\core_1.execute.rf.reg_outputs[2][9] ),
    .A2(_2765_),
    .B1(_2767_),
    .C1(_2760_),
    .X(_0362_));
 sky130_fd_sc_hd__nand2_1 _6011_ (.A(_2649_),
    .B(_2755_),
    .Y(_2768_));
 sky130_fd_sc_hd__o211a_1 _6012_ (.A1(\core_1.execute.rf.reg_outputs[2][10] ),
    .A2(_2765_),
    .B1(_2768_),
    .C1(_2760_),
    .X(_0363_));
 sky130_fd_sc_hd__nand2_1 _6013_ (.A(_2652_),
    .B(_2755_),
    .Y(_2769_));
 sky130_fd_sc_hd__o211a_1 _6014_ (.A1(\core_1.execute.rf.reg_outputs[2][11] ),
    .A2(_2765_),
    .B1(_2769_),
    .C1(_2760_),
    .X(_0364_));
 sky130_fd_sc_hd__nand2_1 _6015_ (.A(_2655_),
    .B(_2755_),
    .Y(_2770_));
 sky130_fd_sc_hd__o211a_1 _6016_ (.A1(\core_1.execute.rf.reg_outputs[2][12] ),
    .A2(_2765_),
    .B1(_2770_),
    .C1(_2760_),
    .X(_0365_));
 sky130_fd_sc_hd__nand2_1 _6017_ (.A(_2658_),
    .B(_2755_),
    .Y(_2771_));
 sky130_fd_sc_hd__buf_4 _6018_ (.A(_1155_),
    .X(_2772_));
 sky130_fd_sc_hd__o211a_1 _6019_ (.A1(\core_1.execute.rf.reg_outputs[2][13] ),
    .A2(_2765_),
    .B1(_2771_),
    .C1(_2772_),
    .X(_0366_));
 sky130_fd_sc_hd__nand2_1 _6020_ (.A(_2662_),
    .B(_2755_),
    .Y(_2773_));
 sky130_fd_sc_hd__o211a_1 _6021_ (.A1(\core_1.execute.rf.reg_outputs[2][14] ),
    .A2(_2765_),
    .B1(_2773_),
    .C1(_2772_),
    .X(_0367_));
 sky130_fd_sc_hd__nand2_1 _6022_ (.A(_2665_),
    .B(_2755_),
    .Y(_2774_));
 sky130_fd_sc_hd__o211a_1 _6023_ (.A1(\core_1.execute.rf.reg_outputs[2][15] ),
    .A2(_2765_),
    .B1(_2774_),
    .C1(_2772_),
    .X(_0368_));
 sky130_fd_sc_hd__nand2_2 _6024_ (.A(\core_1.ew_reg_ie[1] ),
    .B(_2603_),
    .Y(_2775_));
 sky130_fd_sc_hd__and2_2 _6025_ (.A(\core_1.ew_reg_ie[1] ),
    .B(_2602_),
    .X(_2776_));
 sky130_fd_sc_hd__clkbuf_4 _6026_ (.A(_2776_),
    .X(_2777_));
 sky130_fd_sc_hd__or2_1 _6027_ (.A(\core_1.execute.rf.reg_outputs[1][0] ),
    .B(_2777_),
    .X(_2778_));
 sky130_fd_sc_hd__o211a_1 _6028_ (.A1(_2607_),
    .A2(_2775_),
    .B1(_2778_),
    .C1(_2772_),
    .X(_0369_));
 sky130_fd_sc_hd__or2_1 _6029_ (.A(\core_1.execute.rf.reg_outputs[1][1] ),
    .B(_2777_),
    .X(_2779_));
 sky130_fd_sc_hd__o211a_1 _6030_ (.A1(_2613_),
    .A2(_2775_),
    .B1(_2779_),
    .C1(_2772_),
    .X(_0370_));
 sky130_fd_sc_hd__or2_1 _6031_ (.A(\core_1.execute.rf.reg_outputs[1][2] ),
    .B(_2777_),
    .X(_2780_));
 sky130_fd_sc_hd__o211a_1 _6032_ (.A1(_2617_),
    .A2(_2775_),
    .B1(_2780_),
    .C1(_2772_),
    .X(_0371_));
 sky130_fd_sc_hd__or2_1 _6033_ (.A(\core_1.execute.rf.reg_outputs[1][3] ),
    .B(_2777_),
    .X(_2781_));
 sky130_fd_sc_hd__o211a_1 _6034_ (.A1(_2621_),
    .A2(_2775_),
    .B1(_2781_),
    .C1(_2772_),
    .X(_0372_));
 sky130_fd_sc_hd__or2_1 _6035_ (.A(\core_1.execute.rf.reg_outputs[1][4] ),
    .B(_2776_),
    .X(_2782_));
 sky130_fd_sc_hd__o211a_1 _6036_ (.A1(_2626_),
    .A2(_2775_),
    .B1(_2782_),
    .C1(_2772_),
    .X(_0373_));
 sky130_fd_sc_hd__or2_1 _6037_ (.A(\core_1.execute.rf.reg_outputs[1][5] ),
    .B(_2776_),
    .X(_2783_));
 sky130_fd_sc_hd__o211a_1 _6038_ (.A1(_2630_),
    .A2(_2775_),
    .B1(_2783_),
    .C1(_2772_),
    .X(_0374_));
 sky130_fd_sc_hd__or2_1 _6039_ (.A(\core_1.execute.rf.reg_outputs[1][6] ),
    .B(_2776_),
    .X(_2784_));
 sky130_fd_sc_hd__o211a_1 _6040_ (.A1(_2634_),
    .A2(_2775_),
    .B1(_2784_),
    .C1(_2772_),
    .X(_0375_));
 sky130_fd_sc_hd__or2_1 _6041_ (.A(\core_1.execute.rf.reg_outputs[1][7] ),
    .B(_2776_),
    .X(_2785_));
 sky130_fd_sc_hd__clkbuf_4 _6042_ (.A(_1155_),
    .X(_2786_));
 sky130_fd_sc_hd__o211a_1 _6043_ (.A1(_2638_),
    .A2(_2775_),
    .B1(_2785_),
    .C1(_2786_),
    .X(_0376_));
 sky130_fd_sc_hd__clkbuf_4 _6044_ (.A(_2776_),
    .X(_2787_));
 sky130_fd_sc_hd__nand2_1 _6045_ (.A(_2644_),
    .B(_2787_),
    .Y(_2788_));
 sky130_fd_sc_hd__o211a_1 _6046_ (.A1(\core_1.execute.rf.reg_outputs[1][8] ),
    .A2(_2787_),
    .B1(_2788_),
    .C1(_2786_),
    .X(_0377_));
 sky130_fd_sc_hd__nand2_1 _6047_ (.A(_2646_),
    .B(_2787_),
    .Y(_2789_));
 sky130_fd_sc_hd__o211a_1 _6048_ (.A1(\core_1.execute.rf.reg_outputs[1][9] ),
    .A2(_2787_),
    .B1(_2789_),
    .C1(_2786_),
    .X(_0378_));
 sky130_fd_sc_hd__nand2_1 _6049_ (.A(_2649_),
    .B(_2777_),
    .Y(_2790_));
 sky130_fd_sc_hd__o211a_1 _6050_ (.A1(\core_1.execute.rf.reg_outputs[1][10] ),
    .A2(_2787_),
    .B1(_2790_),
    .C1(_2786_),
    .X(_0379_));
 sky130_fd_sc_hd__nand2_1 _6051_ (.A(_2652_),
    .B(_2777_),
    .Y(_2791_));
 sky130_fd_sc_hd__o211a_1 _6052_ (.A1(\core_1.execute.rf.reg_outputs[1][11] ),
    .A2(_2787_),
    .B1(_2791_),
    .C1(_2786_),
    .X(_0380_));
 sky130_fd_sc_hd__nand2_1 _6053_ (.A(_2655_),
    .B(_2777_),
    .Y(_2792_));
 sky130_fd_sc_hd__o211a_1 _6054_ (.A1(\core_1.execute.rf.reg_outputs[1][12] ),
    .A2(_2787_),
    .B1(_2792_),
    .C1(_2786_),
    .X(_0381_));
 sky130_fd_sc_hd__nand2_1 _6055_ (.A(_2658_),
    .B(_2777_),
    .Y(_2793_));
 sky130_fd_sc_hd__o211a_1 _6056_ (.A1(\core_1.execute.rf.reg_outputs[1][13] ),
    .A2(_2787_),
    .B1(_2793_),
    .C1(_2786_),
    .X(_0382_));
 sky130_fd_sc_hd__nand2_1 _6057_ (.A(_2662_),
    .B(_2777_),
    .Y(_2794_));
 sky130_fd_sc_hd__o211a_1 _6058_ (.A1(\core_1.execute.rf.reg_outputs[1][14] ),
    .A2(_2787_),
    .B1(_2794_),
    .C1(_2786_),
    .X(_0383_));
 sky130_fd_sc_hd__nand2_1 _6059_ (.A(_2665_),
    .B(_2777_),
    .Y(_2795_));
 sky130_fd_sc_hd__o211a_1 _6060_ (.A1(\core_1.execute.rf.reg_outputs[1][15] ),
    .A2(_2787_),
    .B1(_2795_),
    .C1(_2786_),
    .X(_0384_));
 sky130_fd_sc_hd__nand2_2 _6061_ (.A(\core_1.ew_reg_ie[0] ),
    .B(_2603_),
    .Y(_2796_));
 sky130_fd_sc_hd__and2_1 _6062_ (.A(\core_1.ew_reg_ie[0] ),
    .B(_2602_),
    .X(_2797_));
 sky130_fd_sc_hd__buf_2 _6063_ (.A(_2797_),
    .X(_2798_));
 sky130_fd_sc_hd__or2_1 _6064_ (.A(net88),
    .B(_2798_),
    .X(_2799_));
 sky130_fd_sc_hd__o211a_1 _6065_ (.A1(_2607_),
    .A2(_2796_),
    .B1(_2799_),
    .C1(_2786_),
    .X(_0385_));
 sky130_fd_sc_hd__or2_1 _6066_ (.A(net95),
    .B(_2798_),
    .X(_2800_));
 sky130_fd_sc_hd__clkbuf_4 _6067_ (.A(_1155_),
    .X(_2801_));
 sky130_fd_sc_hd__o211a_1 _6068_ (.A1(_2613_),
    .A2(_2796_),
    .B1(_2800_),
    .C1(_2801_),
    .X(_0386_));
 sky130_fd_sc_hd__or2_1 _6069_ (.A(net96),
    .B(_2798_),
    .X(_2802_));
 sky130_fd_sc_hd__o211a_1 _6070_ (.A1(_2617_),
    .A2(_2796_),
    .B1(_2802_),
    .C1(_2801_),
    .X(_0387_));
 sky130_fd_sc_hd__or2_1 _6071_ (.A(net97),
    .B(_2798_),
    .X(_2803_));
 sky130_fd_sc_hd__o211a_1 _6072_ (.A1(_2621_),
    .A2(_2796_),
    .B1(_2803_),
    .C1(_2801_),
    .X(_0388_));
 sky130_fd_sc_hd__or2_1 _6073_ (.A(net98),
    .B(_2797_),
    .X(_2804_));
 sky130_fd_sc_hd__o211a_1 _6074_ (.A1(_2626_),
    .A2(_2796_),
    .B1(_2804_),
    .C1(_2801_),
    .X(_0389_));
 sky130_fd_sc_hd__or2_1 _6075_ (.A(net99),
    .B(_2797_),
    .X(_2805_));
 sky130_fd_sc_hd__o211a_1 _6076_ (.A1(_2630_),
    .A2(_2796_),
    .B1(_2805_),
    .C1(_2801_),
    .X(_0390_));
 sky130_fd_sc_hd__or2_1 _6077_ (.A(net100),
    .B(_2797_),
    .X(_2806_));
 sky130_fd_sc_hd__o211a_1 _6078_ (.A1(_2634_),
    .A2(_2796_),
    .B1(_2806_),
    .C1(_2801_),
    .X(_0391_));
 sky130_fd_sc_hd__or2_1 _6079_ (.A(net101),
    .B(_2797_),
    .X(_2807_));
 sky130_fd_sc_hd__o211a_1 _6080_ (.A1(_2638_),
    .A2(_2796_),
    .B1(_2807_),
    .C1(_2801_),
    .X(_0392_));
 sky130_fd_sc_hd__buf_2 _6081_ (.A(_2797_),
    .X(_2808_));
 sky130_fd_sc_hd__nand2_1 _6082_ (.A(_2644_),
    .B(_2808_),
    .Y(_2809_));
 sky130_fd_sc_hd__o211a_1 _6083_ (.A1(net102),
    .A2(_2808_),
    .B1(_2809_),
    .C1(_2801_),
    .X(_0393_));
 sky130_fd_sc_hd__nand2_1 _6084_ (.A(_2646_),
    .B(_2808_),
    .Y(_2810_));
 sky130_fd_sc_hd__o211a_1 _6085_ (.A1(net103),
    .A2(_2808_),
    .B1(_2810_),
    .C1(_2801_),
    .X(_0394_));
 sky130_fd_sc_hd__nand2_1 _6086_ (.A(_2649_),
    .B(_2798_),
    .Y(_2811_));
 sky130_fd_sc_hd__o211a_1 _6087_ (.A1(net89),
    .A2(_2808_),
    .B1(_2811_),
    .C1(_2801_),
    .X(_0395_));
 sky130_fd_sc_hd__nand2_1 _6088_ (.A(_2652_),
    .B(_2798_),
    .Y(_2812_));
 sky130_fd_sc_hd__buf_6 _6089_ (.A(_1155_),
    .X(_2813_));
 sky130_fd_sc_hd__o211a_1 _6090_ (.A1(net90),
    .A2(_2808_),
    .B1(_2812_),
    .C1(_2813_),
    .X(_0396_));
 sky130_fd_sc_hd__nand2_1 _6091_ (.A(_2655_),
    .B(_2798_),
    .Y(_2814_));
 sky130_fd_sc_hd__o211a_1 _6092_ (.A1(net91),
    .A2(_2808_),
    .B1(_2814_),
    .C1(_2813_),
    .X(_0397_));
 sky130_fd_sc_hd__nand2_1 _6093_ (.A(_2658_),
    .B(_2798_),
    .Y(_2815_));
 sky130_fd_sc_hd__o211a_1 _6094_ (.A1(net92),
    .A2(_2808_),
    .B1(_2815_),
    .C1(_2813_),
    .X(_0398_));
 sky130_fd_sc_hd__nand2_1 _6095_ (.A(_2662_),
    .B(_2798_),
    .Y(_2816_));
 sky130_fd_sc_hd__o211a_1 _6096_ (.A1(net93),
    .A2(_2808_),
    .B1(_2816_),
    .C1(_2813_),
    .X(_0399_));
 sky130_fd_sc_hd__nand2_1 _6097_ (.A(_2665_),
    .B(_2798_),
    .Y(_2817_));
 sky130_fd_sc_hd__o211a_1 _6098_ (.A1(net94),
    .A2(_2808_),
    .B1(_2817_),
    .C1(_2813_),
    .X(_0400_));
 sky130_fd_sc_hd__and4_1 _6099_ (.A(_1141_),
    .B(_0643_),
    .C(_1006_),
    .D(_1147_),
    .X(_2818_));
 sky130_fd_sc_hd__nor2_4 _6100_ (.A(_0659_),
    .B(_0667_),
    .Y(_2819_));
 sky130_fd_sc_hd__a21o_1 _6101_ (.A1(_1006_),
    .A2(_1147_),
    .B1(\core_1.execute.irq_en ),
    .X(_2820_));
 sky130_fd_sc_hd__and3b_1 _6102_ (.A_N(_2818_),
    .B(_2819_),
    .C(_2820_),
    .X(_2821_));
 sky130_fd_sc_hd__clkbuf_1 _6103_ (.A(_2821_),
    .X(_0401_));
 sky130_fd_sc_hd__and2_2 _6104_ (.A(\core_1.decode.o_submit ),
    .B(_0860_),
    .X(_2822_));
 sky130_fd_sc_hd__a21o_1 _6105_ (.A1(_1737_),
    .A2(_0728_),
    .B1(_2822_),
    .X(_2823_));
 sky130_fd_sc_hd__mux2_1 _6106_ (.A0(_2823_),
    .A1(_1192_),
    .S(_1760_),
    .X(_2824_));
 sky130_fd_sc_hd__clkbuf_1 _6107_ (.A(_2824_),
    .X(_0402_));
 sky130_fd_sc_hd__nand2_1 _6108_ (.A(_1737_),
    .B(_1193_),
    .Y(_2825_));
 sky130_fd_sc_hd__nand2_1 _6109_ (.A(_1192_),
    .B(_1764_),
    .Y(_2826_));
 sky130_fd_sc_hd__nand2_1 _6110_ (.A(_1765_),
    .B(_1589_),
    .Y(_2827_));
 sky130_fd_sc_hd__o221a_1 _6111_ (.A1(_1743_),
    .A2(_1355_),
    .B1(_2826_),
    .B2(_1354_),
    .C1(_2827_),
    .X(_2828_));
 sky130_fd_sc_hd__o211a_1 _6112_ (.A1(_1352_),
    .A2(_2825_),
    .B1(_2828_),
    .C1(_1191_),
    .X(_2829_));
 sky130_fd_sc_hd__or2_1 _6113_ (.A(_1743_),
    .B(_1373_),
    .X(_2830_));
 sky130_fd_sc_hd__o221a_1 _6114_ (.A1(_1371_),
    .A2(_2826_),
    .B1(_2825_),
    .B2(_1351_),
    .C1(_2830_),
    .X(_2831_));
 sky130_fd_sc_hd__o211a_1 _6115_ (.A1(_1194_),
    .A2(_1804_),
    .B1(_2831_),
    .C1(_1741_),
    .X(_2832_));
 sky130_fd_sc_hd__nand2_1 _6116_ (.A(_1555_),
    .B(_1738_),
    .Y(_2833_));
 sky130_fd_sc_hd__o221a_1 _6117_ (.A1(_1743_),
    .A2(_1827_),
    .B1(_1451_),
    .B2(_1194_),
    .C1(_2833_),
    .X(_2834_));
 sky130_fd_sc_hd__o211a_1 _6118_ (.A1(_1505_),
    .A2(_2825_),
    .B1(_2834_),
    .C1(_1191_),
    .X(_2835_));
 sky130_fd_sc_hd__or2_1 _6119_ (.A(_1599_),
    .B(_2825_),
    .X(_2836_));
 sky130_fd_sc_hd__o221a_1 _6120_ (.A1(_1743_),
    .A2(_1410_),
    .B1(_2826_),
    .B2(_1468_),
    .C1(_2836_),
    .X(_2837_));
 sky130_fd_sc_hd__o211a_1 _6121_ (.A1(_1194_),
    .A2(_1347_),
    .B1(_2837_),
    .C1(_1741_),
    .X(_2838_));
 sky130_fd_sc_hd__or3_1 _6122_ (.A(_1188_),
    .B(_2835_),
    .C(_2838_),
    .X(_2839_));
 sky130_fd_sc_hd__o311a_1 _6123_ (.A1(_1769_),
    .A2(_2829_),
    .A3(_2832_),
    .B1(_2839_),
    .C1(_0860_),
    .X(_2840_));
 sky130_fd_sc_hd__nand2_2 _6124_ (.A(\core_1.execute.alu_mul_div.comp ),
    .B(_2840_),
    .Y(_2841_));
 sky130_fd_sc_hd__and2_2 _6125_ (.A(_0729_),
    .B(_2841_),
    .X(_2842_));
 sky130_fd_sc_hd__clkbuf_4 _6126_ (.A(_2842_),
    .X(_2843_));
 sky130_fd_sc_hd__nor2_2 _6127_ (.A(_0729_),
    .B(_1407_),
    .Y(_2844_));
 sky130_fd_sc_hd__clkbuf_4 _6128_ (.A(_2844_),
    .X(_2845_));
 sky130_fd_sc_hd__nor2_4 _6129_ (.A(\core_1.decode.o_submit ),
    .B(_2841_),
    .Y(_2846_));
 sky130_fd_sc_hd__nor2_1 _6130_ (.A(\core_1.execute.alu_mul_div.cbit[0] ),
    .B(\core_1.execute.alu_mul_div.cbit[1] ),
    .Y(_2847_));
 sky130_fd_sc_hd__nand2_1 _6131_ (.A(_1189_),
    .B(_2847_),
    .Y(_2848_));
 sky130_fd_sc_hd__or4_1 _6132_ (.A(\core_1.execute.alu_mul_div.cbit[3] ),
    .B(_2073_),
    .C(_2848_),
    .D(_2041_),
    .X(_2849_));
 sky130_fd_sc_hd__a31o_1 _6133_ (.A1(_1769_),
    .A2(_1744_),
    .A3(_1346_),
    .B1(\core_1.execute.alu_mul_div.mul_res[0] ),
    .X(_2850_));
 sky130_fd_sc_hd__and3_1 _6134_ (.A(_2846_),
    .B(_2849_),
    .C(_2850_),
    .X(_2851_));
 sky130_fd_sc_hd__a221o_1 _6135_ (.A1(\core_1.execute.alu_mul_div.mul_res[0] ),
    .A2(_2843_),
    .B1(_2845_),
    .B2(_1346_),
    .C1(_2851_),
    .X(_0403_));
 sky130_fd_sc_hd__and3_1 _6136_ (.A(\core_1.execute.alu_mul_div.cbit[0] ),
    .B(_1343_),
    .C(_1345_),
    .X(_2852_));
 sky130_fd_sc_hd__o211a_4 _6137_ (.A1(net95),
    .A2(_1377_),
    .B1(_1402_),
    .C1(_1736_),
    .X(_2853_));
 sky130_fd_sc_hd__o2111a_1 _6138_ (.A1(_2852_),
    .A2(_2853_),
    .B1(_1768_),
    .C1(_1189_),
    .D1(_1751_),
    .X(_2854_));
 sky130_fd_sc_hd__xnor2_1 _6139_ (.A(\core_1.execute.alu_mul_div.mul_res[1] ),
    .B(_2854_),
    .Y(_2855_));
 sky130_fd_sc_hd__nand2_1 _6140_ (.A(_2849_),
    .B(_2855_),
    .Y(_2856_));
 sky130_fd_sc_hd__or2_1 _6141_ (.A(_2849_),
    .B(_2855_),
    .X(_2857_));
 sky130_fd_sc_hd__a32o_1 _6142_ (.A1(_2846_),
    .A2(_2856_),
    .A3(_2857_),
    .B1(_2843_),
    .B2(\core_1.execute.alu_mul_div.mul_res[1] ),
    .X(_2858_));
 sky130_fd_sc_hd__a21o_1 _6143_ (.A1(_1404_),
    .A2(_2845_),
    .B1(_2858_),
    .X(_0404_));
 sky130_fd_sc_hd__clkinv_2 _6144_ (.A(_2843_),
    .Y(_2859_));
 sky130_fd_sc_hd__and4_1 _6145_ (.A(_1768_),
    .B(_1189_),
    .C(\core_1.execute.alu_mul_div.mul_res[2] ),
    .D(_1753_),
    .X(_2860_));
 sky130_fd_sc_hd__a31oi_1 _6146_ (.A1(_1768_),
    .A2(_1190_),
    .A3(_1753_),
    .B1(\core_1.execute.alu_mul_div.mul_res[2] ),
    .Y(_2861_));
 sky130_fd_sc_hd__nand2_1 _6147_ (.A(\core_1.execute.alu_mul_div.mul_res[1] ),
    .B(_2854_),
    .Y(_2862_));
 sky130_fd_sc_hd__o211ai_1 _6148_ (.A1(_2860_),
    .A2(_2861_),
    .B1(_2862_),
    .C1(_2857_),
    .Y(_2863_));
 sky130_fd_sc_hd__a211o_1 _6149_ (.A1(_2862_),
    .A2(_2857_),
    .B1(_2860_),
    .C1(_2861_),
    .X(_2864_));
 sky130_fd_sc_hd__and3_1 _6150_ (.A(_0729_),
    .B(_2863_),
    .C(_2864_),
    .X(_2865_));
 sky130_fd_sc_hd__a211o_1 _6151_ (.A1(_1820_),
    .A2(_2844_),
    .B1(_2865_),
    .C1(_2843_),
    .X(_2866_));
 sky130_fd_sc_hd__o21a_1 _6152_ (.A1(\core_1.execute.alu_mul_div.mul_res[2] ),
    .A2(_2859_),
    .B1(_2866_),
    .X(_0405_));
 sky130_fd_sc_hd__nand2_1 _6153_ (.A(_1190_),
    .B(_1753_),
    .Y(_2867_));
 sky130_fd_sc_hd__or3b_1 _6154_ (.A(_2867_),
    .B(_1187_),
    .C_N(\core_1.execute.alu_mul_div.mul_res[2] ),
    .X(_2868_));
 sky130_fd_sc_hd__mux4_1 _6155_ (.A0(_2041_),
    .A1(_1403_),
    .A2(_1562_),
    .A3(_1553_),
    .S0(_1737_),
    .S1(_1751_),
    .X(_2869_));
 sky130_fd_sc_hd__or2_1 _6156_ (.A(\core_1.execute.alu_mul_div.cbit[2] ),
    .B(_2869_),
    .X(_2870_));
 sky130_fd_sc_hd__or3b_1 _6157_ (.A(_2870_),
    .B(_1187_),
    .C_N(\core_1.execute.alu_mul_div.mul_res[3] ),
    .X(_2871_));
 sky130_fd_sc_hd__o21bai_1 _6158_ (.A1(_1187_),
    .A2(_2870_),
    .B1_N(\core_1.execute.alu_mul_div.mul_res[3] ),
    .Y(_2872_));
 sky130_fd_sc_hd__nand2_1 _6159_ (.A(_2871_),
    .B(_2872_),
    .Y(_2873_));
 sky130_fd_sc_hd__a31o_1 _6160_ (.A1(_2868_),
    .A2(_2864_),
    .A3(_2873_),
    .B1(_2822_),
    .X(_2874_));
 sky130_fd_sc_hd__a21o_1 _6161_ (.A1(_2868_),
    .A2(_2864_),
    .B1(_2873_),
    .X(_2875_));
 sky130_fd_sc_hd__and2b_1 _6162_ (.A_N(_2874_),
    .B(_2875_),
    .X(_2876_));
 sky130_fd_sc_hd__a31o_1 _6163_ (.A1(_2822_),
    .A2(_1827_),
    .A3(_1817_),
    .B1(_2842_),
    .X(_2877_));
 sky130_fd_sc_hd__o22a_1 _6164_ (.A1(\core_1.execute.alu_mul_div.mul_res[3] ),
    .A2(_2859_),
    .B1(_2876_),
    .B2(_2877_),
    .X(_0406_));
 sky130_fd_sc_hd__nor2_1 _6165_ (.A(_1189_),
    .B(_1743_),
    .Y(_2878_));
 sky130_fd_sc_hd__mux4_1 _6166_ (.A0(_1404_),
    .A1(_1817_),
    .A2(_1820_),
    .A3(_1815_),
    .S0(_1764_),
    .S1(_1737_),
    .X(_2879_));
 sky130_fd_sc_hd__a22o_1 _6167_ (.A1(_1346_),
    .A2(_2878_),
    .B1(_2879_),
    .B2(_1190_),
    .X(_2880_));
 sky130_fd_sc_hd__and3_1 _6168_ (.A(_1768_),
    .B(\core_1.execute.alu_mul_div.mul_res[4] ),
    .C(_2880_),
    .X(_2881_));
 sky130_fd_sc_hd__a21oi_1 _6169_ (.A1(_1768_),
    .A2(_2880_),
    .B1(\core_1.execute.alu_mul_div.mul_res[4] ),
    .Y(_2882_));
 sky130_fd_sc_hd__or2_1 _6170_ (.A(_2881_),
    .B(_2882_),
    .X(_2883_));
 sky130_fd_sc_hd__a21oi_1 _6171_ (.A1(_2871_),
    .A2(_2875_),
    .B1(_2883_),
    .Y(_2884_));
 sky130_fd_sc_hd__a31o_1 _6172_ (.A1(_2871_),
    .A2(_2875_),
    .A3(_2883_),
    .B1(_2822_),
    .X(_2885_));
 sky130_fd_sc_hd__nor2_1 _6173_ (.A(_2884_),
    .B(_2885_),
    .Y(_2886_));
 sky130_fd_sc_hd__a211o_1 _6174_ (.A1(_1815_),
    .A2(_2844_),
    .B1(_2886_),
    .C1(_2843_),
    .X(_2887_));
 sky130_fd_sc_hd__o21a_1 _6175_ (.A1(\core_1.execute.alu_mul_div.mul_res[4] ),
    .A2(_2859_),
    .B1(_2887_),
    .X(_0407_));
 sky130_fd_sc_hd__o21ai_1 _6176_ (.A1(_2852_),
    .A2(_2853_),
    .B1(_1764_),
    .Y(_2888_));
 sky130_fd_sc_hd__mux4_1 _6177_ (.A0(_1523_),
    .A1(_1547_),
    .A2(_1553_),
    .A3(_1562_),
    .S0(\core_1.execute.alu_mul_div.cbit[0] ),
    .S1(_1193_),
    .X(_2889_));
 sky130_fd_sc_hd__mux2_1 _6178_ (.A0(_2888_),
    .A1(_2889_),
    .S(_1190_),
    .X(_2890_));
 sky130_fd_sc_hd__nor2_1 _6179_ (.A(_1187_),
    .B(_2890_),
    .Y(_2891_));
 sky130_fd_sc_hd__xnor2_1 _6180_ (.A(\core_1.execute.alu_mul_div.mul_res[5] ),
    .B(_2891_),
    .Y(_2892_));
 sky130_fd_sc_hd__or3b_1 _6181_ (.A(_2881_),
    .B(_2884_),
    .C_N(_2892_),
    .X(_2893_));
 sky130_fd_sc_hd__o21bai_1 _6182_ (.A1(_2881_),
    .A2(_2884_),
    .B1_N(_2892_),
    .Y(_2894_));
 sky130_fd_sc_hd__a22o_1 _6183_ (.A1(\core_1.execute.alu_mul_div.mul_res[5] ),
    .A2(_2842_),
    .B1(_2845_),
    .B2(_1522_),
    .X(_2895_));
 sky130_fd_sc_hd__a31o_1 _6184_ (.A1(_2846_),
    .A2(_2893_),
    .A3(_2894_),
    .B1(_2895_),
    .X(_0408_));
 sky130_fd_sc_hd__nand2_1 _6185_ (.A(\core_1.execute.alu_mul_div.mul_res[5] ),
    .B(_2891_),
    .Y(_2896_));
 sky130_fd_sc_hd__nor2_1 _6186_ (.A(_1187_),
    .B(_1755_),
    .Y(_2897_));
 sky130_fd_sc_hd__xnor2_1 _6187_ (.A(\core_1.execute.alu_mul_div.mul_res[6] ),
    .B(_2897_),
    .Y(_2898_));
 sky130_fd_sc_hd__nand3_1 _6188_ (.A(_2896_),
    .B(_2894_),
    .C(_2898_),
    .Y(_2899_));
 sky130_fd_sc_hd__a21o_1 _6189_ (.A1(_2896_),
    .A2(_2894_),
    .B1(_2898_),
    .X(_2900_));
 sky130_fd_sc_hd__a22o_1 _6190_ (.A1(\core_1.execute.alu_mul_div.mul_res[6] ),
    .A2(_2842_),
    .B1(_2845_),
    .B2(_1811_),
    .X(_2901_));
 sky130_fd_sc_hd__a31o_1 _6191_ (.A1(_2846_),
    .A2(_2899_),
    .A3(_2900_),
    .B1(_2901_),
    .X(_0409_));
 sky130_fd_sc_hd__nand2_1 _6192_ (.A(\core_1.execute.alu_mul_div.mul_res[6] ),
    .B(_2897_),
    .Y(_2902_));
 sky130_fd_sc_hd__mux2_1 _6193_ (.A0(_1523_),
    .A1(_1547_),
    .S(_1192_),
    .X(_2903_));
 sky130_fd_sc_hd__mux2_1 _6194_ (.A0(_1811_),
    .A1(_1531_),
    .S(_1737_),
    .X(_2904_));
 sky130_fd_sc_hd__clkinv_2 _6195_ (.A(_2904_),
    .Y(_2905_));
 sky130_fd_sc_hd__mux2_1 _6196_ (.A0(_2903_),
    .A1(_2905_),
    .S(_1764_),
    .X(_2906_));
 sky130_fd_sc_hd__mux2_1 _6197_ (.A0(_2869_),
    .A1(_2906_),
    .S(_1190_),
    .X(_2907_));
 sky130_fd_sc_hd__or3b_1 _6198_ (.A(_2907_),
    .B(_1187_),
    .C_N(\core_1.execute.alu_mul_div.mul_res[7] ),
    .X(_2908_));
 sky130_fd_sc_hd__o21bai_1 _6199_ (.A1(_1187_),
    .A2(_2907_),
    .B1_N(\core_1.execute.alu_mul_div.mul_res[7] ),
    .Y(_2909_));
 sky130_fd_sc_hd__nand2_1 _6200_ (.A(_2908_),
    .B(_2909_),
    .Y(_2910_));
 sky130_fd_sc_hd__nand3_1 _6201_ (.A(_2902_),
    .B(_2900_),
    .C(_2910_),
    .Y(_2911_));
 sky130_fd_sc_hd__a21o_1 _6202_ (.A1(_2902_),
    .A2(_2900_),
    .B1(_2910_),
    .X(_2912_));
 sky130_fd_sc_hd__a22o_1 _6203_ (.A1(\core_1.execute.alu_mul_div.mul_res[7] ),
    .A2(_2842_),
    .B1(_2844_),
    .B2(_1531_),
    .X(_2913_));
 sky130_fd_sc_hd__a31o_1 _6204_ (.A1(_2846_),
    .A2(_2911_),
    .A3(_2912_),
    .B1(_2913_),
    .X(_0410_));
 sky130_fd_sc_hd__mux4_1 _6205_ (.A0(_1811_),
    .A1(_1522_),
    .A2(_1746_),
    .A3(_1531_),
    .S0(_1192_),
    .S1(_1764_),
    .X(_2914_));
 sky130_fd_sc_hd__or2_1 _6206_ (.A(\core_1.execute.alu_mul_div.cbit[2] ),
    .B(_2914_),
    .X(_2915_));
 sky130_fd_sc_hd__o211a_1 _6207_ (.A1(_1190_),
    .A2(_2879_),
    .B1(_2915_),
    .C1(_1769_),
    .X(_2916_));
 sky130_fd_sc_hd__a31o_1 _6208_ (.A1(_1187_),
    .A2(_1744_),
    .A3(_1346_),
    .B1(_2916_),
    .X(_2917_));
 sky130_fd_sc_hd__and2_1 _6209_ (.A(\core_1.execute.alu_mul_div.mul_res[8] ),
    .B(_2917_),
    .X(_2918_));
 sky130_fd_sc_hd__nor2_1 _6210_ (.A(\core_1.execute.alu_mul_div.mul_res[8] ),
    .B(_2917_),
    .Y(_2919_));
 sky130_fd_sc_hd__or2_1 _6211_ (.A(_2918_),
    .B(_2919_),
    .X(_2920_));
 sky130_fd_sc_hd__and3_1 _6212_ (.A(_2908_),
    .B(_2912_),
    .C(_2920_),
    .X(_2921_));
 sky130_fd_sc_hd__a21oi_1 _6213_ (.A1(_2908_),
    .A2(_2912_),
    .B1(_2920_),
    .Y(_2922_));
 sky130_fd_sc_hd__nor2_1 _6214_ (.A(_2921_),
    .B(_2922_),
    .Y(_2923_));
 sky130_fd_sc_hd__a22o_1 _6215_ (.A1(\core_1.execute.alu_mul_div.mul_res[8] ),
    .A2(_2843_),
    .B1(_2845_),
    .B2(_1746_),
    .X(_2924_));
 sky130_fd_sc_hd__a21o_1 _6216_ (.A1(_2846_),
    .A2(_2923_),
    .B1(_2924_),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_1 _6217_ (.A0(_1465_),
    .A1(_1746_),
    .S(_1192_),
    .X(_2925_));
 sky130_fd_sc_hd__mux2_1 _6218_ (.A0(_2904_),
    .A1(_2925_),
    .S(_1764_),
    .X(_2926_));
 sky130_fd_sc_hd__nor2_1 _6219_ (.A(_1741_),
    .B(_2926_),
    .Y(_2927_));
 sky130_fd_sc_hd__a211o_1 _6220_ (.A1(_1741_),
    .A2(_2889_),
    .B1(_2927_),
    .C1(_1187_),
    .X(_2928_));
 sky130_fd_sc_hd__o31ai_1 _6221_ (.A1(_1769_),
    .A2(_1741_),
    .A3(_2888_),
    .B1(_2928_),
    .Y(_2929_));
 sky130_fd_sc_hd__and2_1 _6222_ (.A(\core_1.execute.alu_mul_div.mul_res[9] ),
    .B(_2929_),
    .X(_2930_));
 sky130_fd_sc_hd__nor2_1 _6223_ (.A(\core_1.execute.alu_mul_div.mul_res[9] ),
    .B(_2929_),
    .Y(_2931_));
 sky130_fd_sc_hd__nor2_1 _6224_ (.A(_2930_),
    .B(_2931_),
    .Y(_2932_));
 sky130_fd_sc_hd__nor3_1 _6225_ (.A(_2918_),
    .B(_2922_),
    .C(_2932_),
    .Y(_2933_));
 sky130_fd_sc_hd__o21a_1 _6226_ (.A1(_2918_),
    .A2(_2922_),
    .B1(_2932_),
    .X(_2934_));
 sky130_fd_sc_hd__nor2_1 _6227_ (.A(_2933_),
    .B(_2934_),
    .Y(_2935_));
 sky130_fd_sc_hd__a22o_1 _6228_ (.A1(\core_1.execute.alu_mul_div.mul_res[9] ),
    .A2(_2843_),
    .B1(_2845_),
    .B2(_1465_),
    .X(_2936_));
 sky130_fd_sc_hd__a21o_1 _6229_ (.A1(_2846_),
    .A2(_2935_),
    .B1(_2936_),
    .X(_0412_));
 sky130_fd_sc_hd__nor2_1 _6230_ (.A(_1190_),
    .B(_1749_),
    .Y(_2937_));
 sky130_fd_sc_hd__a211o_1 _6231_ (.A1(_1190_),
    .A2(_1747_),
    .B1(_2937_),
    .C1(_1188_),
    .X(_2938_));
 sky130_fd_sc_hd__nand2_1 _6232_ (.A(_1188_),
    .B(_2867_),
    .Y(_2939_));
 sky130_fd_sc_hd__and3_1 _6233_ (.A(\core_1.execute.alu_mul_div.mul_res[10] ),
    .B(_2938_),
    .C(_2939_),
    .X(_2940_));
 sky130_fd_sc_hd__a21oi_1 _6234_ (.A1(_2938_),
    .A2(_2939_),
    .B1(\core_1.execute.alu_mul_div.mul_res[10] ),
    .Y(_2941_));
 sky130_fd_sc_hd__nor2_1 _6235_ (.A(_2940_),
    .B(_2941_),
    .Y(_2942_));
 sky130_fd_sc_hd__nor3_1 _6236_ (.A(_2930_),
    .B(_2934_),
    .C(_2942_),
    .Y(_2943_));
 sky130_fd_sc_hd__o21a_1 _6237_ (.A1(_2930_),
    .A2(_2934_),
    .B1(_2942_),
    .X(_2944_));
 sky130_fd_sc_hd__nor2_1 _6238_ (.A(_2943_),
    .B(_2944_),
    .Y(_2945_));
 sky130_fd_sc_hd__a22o_1 _6239_ (.A1(\core_1.execute.alu_mul_div.mul_res[10] ),
    .A2(_2842_),
    .B1(_2845_),
    .B2(_1457_),
    .X(_2946_));
 sky130_fd_sc_hd__a21o_1 _6240_ (.A1(_2846_),
    .A2(_2945_),
    .B1(_2946_),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_1 _6241_ (.A0(_1457_),
    .A1(_1734_),
    .S(_1737_),
    .X(_2947_));
 sky130_fd_sc_hd__or2_1 _6242_ (.A(_1764_),
    .B(_2925_),
    .X(_2948_));
 sky130_fd_sc_hd__o21ai_1 _6243_ (.A1(_1193_),
    .A2(_2947_),
    .B1(_2948_),
    .Y(_2949_));
 sky130_fd_sc_hd__mux2_1 _6244_ (.A0(_2906_),
    .A1(_2949_),
    .S(_1190_),
    .X(_2950_));
 sky130_fd_sc_hd__and2_1 _6245_ (.A(_1188_),
    .B(_2870_),
    .X(_2951_));
 sky130_fd_sc_hd__a21oi_1 _6246_ (.A1(_1769_),
    .A2(_2950_),
    .B1(_2951_),
    .Y(_2952_));
 sky130_fd_sc_hd__and2_1 _6247_ (.A(\core_1.execute.alu_mul_div.mul_res[11] ),
    .B(_2952_),
    .X(_2953_));
 sky130_fd_sc_hd__nor2_1 _6248_ (.A(\core_1.execute.alu_mul_div.mul_res[11] ),
    .B(_2952_),
    .Y(_2954_));
 sky130_fd_sc_hd__or2_1 _6249_ (.A(_2953_),
    .B(_2954_),
    .X(_2955_));
 sky130_fd_sc_hd__or3b_1 _6250_ (.A(_2940_),
    .B(_2944_),
    .C_N(_2955_),
    .X(_2956_));
 sky130_fd_sc_hd__o21ba_1 _6251_ (.A1(_2940_),
    .A2(_2944_),
    .B1_N(_2955_),
    .X(_2957_));
 sky130_fd_sc_hd__and2b_1 _6252_ (.A_N(_2957_),
    .B(_2846_),
    .X(_2958_));
 sky130_fd_sc_hd__a22o_1 _6253_ (.A1(\core_1.execute.alu_mul_div.mul_res[11] ),
    .A2(_2842_),
    .B1(_2845_),
    .B2(_1734_),
    .X(_2959_));
 sky130_fd_sc_hd__a21o_1 _6254_ (.A1(_2956_),
    .A2(_2958_),
    .B1(_2959_),
    .X(_0414_));
 sky130_fd_sc_hd__mux4_1 _6255_ (.A0(_1457_),
    .A1(_1465_),
    .A2(_1477_),
    .A3(_1734_),
    .S0(_1192_),
    .S1(_1764_),
    .X(_2960_));
 sky130_fd_sc_hd__mux2_1 _6256_ (.A0(_2914_),
    .A1(_2960_),
    .S(_1191_),
    .X(_2961_));
 sky130_fd_sc_hd__mux2_1 _6257_ (.A0(_2880_),
    .A1(_2961_),
    .S(_1769_),
    .X(_2962_));
 sky130_fd_sc_hd__nand2_1 _6258_ (.A(\core_1.execute.alu_mul_div.mul_res[12] ),
    .B(_2962_),
    .Y(_2963_));
 sky130_fd_sc_hd__or2_1 _6259_ (.A(\core_1.execute.alu_mul_div.mul_res[12] ),
    .B(_2962_),
    .X(_2964_));
 sky130_fd_sc_hd__nand2_1 _6260_ (.A(_2963_),
    .B(_2964_),
    .Y(_2965_));
 sky130_fd_sc_hd__o21bai_1 _6261_ (.A1(_2953_),
    .A2(_2957_),
    .B1_N(_2965_),
    .Y(_2966_));
 sky130_fd_sc_hd__or3b_1 _6262_ (.A(_2953_),
    .B(_2957_),
    .C_N(_2965_),
    .X(_2967_));
 sky130_fd_sc_hd__a32o_1 _6263_ (.A1(_0729_),
    .A2(_2966_),
    .A3(_2967_),
    .B1(_1477_),
    .B2(_2844_),
    .X(_2968_));
 sky130_fd_sc_hd__and3_1 _6264_ (.A(\core_1.execute.alu_mul_div.mul_res[12] ),
    .B(_0729_),
    .C(_2841_),
    .X(_2969_));
 sky130_fd_sc_hd__a21o_1 _6265_ (.A1(_2859_),
    .A2(_2968_),
    .B1(_2969_),
    .X(_0415_));
 sky130_fd_sc_hd__clkinv_2 _6266_ (.A(_2890_),
    .Y(_2970_));
 sky130_fd_sc_hd__mux2_1 _6267_ (.A0(_1477_),
    .A1(_1493_),
    .S(_1737_),
    .X(_2971_));
 sky130_fd_sc_hd__mux4_1 _6268_ (.A0(_2904_),
    .A1(_2925_),
    .A2(_2947_),
    .A3(_2971_),
    .S0(_1764_),
    .S1(_1191_),
    .X(_2972_));
 sky130_fd_sc_hd__mux2_1 _6269_ (.A0(_2970_),
    .A1(_2972_),
    .S(_1769_),
    .X(_2973_));
 sky130_fd_sc_hd__nand2_1 _6270_ (.A(\core_1.execute.alu_mul_div.mul_res[13] ),
    .B(_2973_),
    .Y(_2974_));
 sky130_fd_sc_hd__or2_1 _6271_ (.A(\core_1.execute.alu_mul_div.mul_res[13] ),
    .B(_2973_),
    .X(_2975_));
 sky130_fd_sc_hd__nand2_1 _6272_ (.A(_2974_),
    .B(_2975_),
    .Y(_2976_));
 sky130_fd_sc_hd__nand3_1 _6273_ (.A(_2963_),
    .B(_2966_),
    .C(_2976_),
    .Y(_2977_));
 sky130_fd_sc_hd__a21o_1 _6274_ (.A1(_2963_),
    .A2(_2966_),
    .B1(_2976_),
    .X(_2978_));
 sky130_fd_sc_hd__and3_1 _6275_ (.A(_2846_),
    .B(_2977_),
    .C(_2978_),
    .X(_2979_));
 sky130_fd_sc_hd__a221o_1 _6276_ (.A1(\core_1.execute.alu_mul_div.mul_res[13] ),
    .A2(_2843_),
    .B1(_2845_),
    .B2(_1493_),
    .C1(_2979_),
    .X(_0416_));
 sky130_fd_sc_hd__inv_2 _6277_ (.A(\core_1.execute.alu_mul_div.mul_res[14] ),
    .Y(_2980_));
 sky130_fd_sc_hd__or2_1 _6278_ (.A(_2980_),
    .B(_1756_),
    .X(_2981_));
 sky130_fd_sc_hd__nand2_1 _6279_ (.A(_2980_),
    .B(_1756_),
    .Y(_2982_));
 sky130_fd_sc_hd__nand2_1 _6280_ (.A(_2981_),
    .B(_2982_),
    .Y(_2983_));
 sky130_fd_sc_hd__a31o_1 _6281_ (.A1(_2974_),
    .A2(_2978_),
    .A3(_2983_),
    .B1(_2822_),
    .X(_2984_));
 sky130_fd_sc_hd__a21o_1 _6282_ (.A1(_2974_),
    .A2(_2978_),
    .B1(_2983_),
    .X(_2985_));
 sky130_fd_sc_hd__and2b_1 _6283_ (.A_N(_2984_),
    .B(_2985_),
    .X(_2986_));
 sky130_fd_sc_hd__a21o_1 _6284_ (.A1(_1745_),
    .A2(_2844_),
    .B1(_2843_),
    .X(_2987_));
 sky130_fd_sc_hd__o22a_1 _6285_ (.A1(\core_1.execute.alu_mul_div.mul_res[14] ),
    .A2(_2859_),
    .B1(_2986_),
    .B2(_2987_),
    .X(_0417_));
 sky130_fd_sc_hd__o22a_1 _6286_ (.A1(_1743_),
    .A2(_1389_),
    .B1(_1500_),
    .B2(_2826_),
    .X(_2988_));
 sky130_fd_sc_hd__a21oi_1 _6287_ (.A1(_1193_),
    .A2(_2971_),
    .B1(_1741_),
    .Y(_2989_));
 sky130_fd_sc_hd__a22o_1 _6288_ (.A1(_1741_),
    .A2(_2949_),
    .B1(_2988_),
    .B2(_2989_),
    .X(_2990_));
 sky130_fd_sc_hd__mux2_1 _6289_ (.A0(_2907_),
    .A1(_2990_),
    .S(_1769_),
    .X(_2991_));
 sky130_fd_sc_hd__xor2_1 _6290_ (.A(\core_1.execute.alu_mul_div.mul_res[15] ),
    .B(_2991_),
    .X(_2992_));
 sky130_fd_sc_hd__a21oi_1 _6291_ (.A1(_2981_),
    .A2(_2985_),
    .B1(_2992_),
    .Y(_2993_));
 sky130_fd_sc_hd__a311o_1 _6292_ (.A1(_2981_),
    .A2(_2985_),
    .A3(_2992_),
    .B1(_2841_),
    .C1(\core_1.decode.o_submit ),
    .X(_2994_));
 sky130_fd_sc_hd__a22oi_1 _6293_ (.A1(\core_1.execute.alu_mul_div.mul_res[15] ),
    .A2(_2843_),
    .B1(_2845_),
    .B2(_1733_),
    .Y(_2995_));
 sky130_fd_sc_hd__o21ai_1 _6294_ (.A1(_2993_),
    .A2(_2994_),
    .B1(_2995_),
    .Y(_0418_));
 sky130_fd_sc_hd__nor2_1 _6295_ (.A(_1056_),
    .B(_0726_),
    .Y(_0419_));
 sky130_fd_sc_hd__nand2_1 _6296_ (.A(_1637_),
    .B(_1638_),
    .Y(_2996_));
 sky130_fd_sc_hd__nor2_1 _6297_ (.A(_1197_),
    .B(_2996_),
    .Y(_2997_));
 sky130_fd_sc_hd__o21a_1 _6298_ (.A1(\core_1.execute.alu_mul_div.div_res[0] ),
    .A2(_2997_),
    .B1(_1654_),
    .X(_0420_));
 sky130_fd_sc_hd__nor2_2 _6299_ (.A(_1769_),
    .B(_2996_),
    .Y(_2998_));
 sky130_fd_sc_hd__a31o_1 _6300_ (.A1(_1763_),
    .A2(_1752_),
    .A3(_2998_),
    .B1(\core_1.execute.alu_mul_div.div_res[1] ),
    .X(_2999_));
 sky130_fd_sc_hd__and2_1 _6301_ (.A(_1653_),
    .B(_2999_),
    .X(_3000_));
 sky130_fd_sc_hd__clkbuf_1 _6302_ (.A(_3000_),
    .X(_0421_));
 sky130_fd_sc_hd__a31o_1 _6303_ (.A1(_1763_),
    .A2(_1738_),
    .A3(_2998_),
    .B1(\core_1.execute.alu_mul_div.div_res[2] ),
    .X(_3001_));
 sky130_fd_sc_hd__and2_1 _6304_ (.A(_1653_),
    .B(_3001_),
    .X(_3002_));
 sky130_fd_sc_hd__clkbuf_1 _6305_ (.A(_3002_),
    .X(_0422_));
 sky130_fd_sc_hd__a31o_1 _6306_ (.A1(_1763_),
    .A2(_2847_),
    .A3(_2998_),
    .B1(\core_1.execute.alu_mul_div.div_res[3] ),
    .X(_3003_));
 sky130_fd_sc_hd__and2_1 _6307_ (.A(_1653_),
    .B(_3003_),
    .X(_3004_));
 sky130_fd_sc_hd__clkbuf_1 _6308_ (.A(_3004_),
    .X(_0423_));
 sky130_fd_sc_hd__and2_1 _6309_ (.A(\core_1.decode.o_submit ),
    .B(_1314_),
    .X(_3005_));
 sky130_fd_sc_hd__nor2_1 _6310_ (.A(_1763_),
    .B(_1194_),
    .Y(_3006_));
 sky130_fd_sc_hd__a21oi_1 _6311_ (.A1(_2998_),
    .A2(_3006_),
    .B1(\core_1.execute.alu_mul_div.div_res[4] ),
    .Y(_3007_));
 sky130_fd_sc_hd__nor2_1 _6312_ (.A(_3005_),
    .B(_3007_),
    .Y(_0424_));
 sky130_fd_sc_hd__and3_1 _6313_ (.A(_1191_),
    .B(_1752_),
    .C(_2998_),
    .X(_3008_));
 sky130_fd_sc_hd__o21a_1 _6314_ (.A1(\core_1.execute.alu_mul_div.div_res[5] ),
    .A2(_3008_),
    .B1(_1654_),
    .X(_0425_));
 sky130_fd_sc_hd__and3_1 _6315_ (.A(_1191_),
    .B(_1738_),
    .C(_2998_),
    .X(_3009_));
 sky130_fd_sc_hd__o21a_1 _6316_ (.A1(\core_1.execute.alu_mul_div.div_res[6] ),
    .A2(_3009_),
    .B1(_1654_),
    .X(_0426_));
 sky130_fd_sc_hd__a21oi_1 _6317_ (.A1(_1744_),
    .A2(_2998_),
    .B1(\core_1.execute.alu_mul_div.div_res[7] ),
    .Y(_3010_));
 sky130_fd_sc_hd__nor2_1 _6318_ (.A(_3005_),
    .B(_3010_),
    .Y(_0427_));
 sky130_fd_sc_hd__nor2_2 _6319_ (.A(_1188_),
    .B(_2996_),
    .Y(_3011_));
 sky130_fd_sc_hd__a31o_1 _6320_ (.A1(_1763_),
    .A2(_1765_),
    .A3(_3011_),
    .B1(\core_1.execute.alu_mul_div.div_res[8] ),
    .X(_3012_));
 sky130_fd_sc_hd__and2_1 _6321_ (.A(_1653_),
    .B(_3012_),
    .X(_3013_));
 sky130_fd_sc_hd__clkbuf_1 _6322_ (.A(_3013_),
    .X(_0428_));
 sky130_fd_sc_hd__a31o_1 _6323_ (.A1(_1763_),
    .A2(_1752_),
    .A3(_3011_),
    .B1(\core_1.execute.alu_mul_div.div_res[9] ),
    .X(_3014_));
 sky130_fd_sc_hd__and2_1 _6324_ (.A(_1653_),
    .B(_3014_),
    .X(_3015_));
 sky130_fd_sc_hd__clkbuf_1 _6325_ (.A(_3015_),
    .X(_0429_));
 sky130_fd_sc_hd__a31o_1 _6326_ (.A1(_1763_),
    .A2(_1738_),
    .A3(_3011_),
    .B1(\core_1.execute.alu_mul_div.div_res[10] ),
    .X(_3016_));
 sky130_fd_sc_hd__and2_1 _6327_ (.A(_1653_),
    .B(_3016_),
    .X(_3017_));
 sky130_fd_sc_hd__clkbuf_1 _6328_ (.A(_3017_),
    .X(_0430_));
 sky130_fd_sc_hd__a31o_1 _6329_ (.A1(_1763_),
    .A2(_2847_),
    .A3(_3011_),
    .B1(\core_1.execute.alu_mul_div.div_res[11] ),
    .X(_3018_));
 sky130_fd_sc_hd__and2_1 _6330_ (.A(_1653_),
    .B(_3018_),
    .X(_3019_));
 sky130_fd_sc_hd__clkbuf_1 _6331_ (.A(_3019_),
    .X(_0431_));
 sky130_fd_sc_hd__a21oi_1 _6332_ (.A1(_3006_),
    .A2(_3011_),
    .B1(\core_1.execute.alu_mul_div.div_res[12] ),
    .Y(_3020_));
 sky130_fd_sc_hd__nor2_1 _6333_ (.A(_3005_),
    .B(_3020_),
    .Y(_0432_));
 sky130_fd_sc_hd__and3_1 _6334_ (.A(_1191_),
    .B(_1752_),
    .C(_3011_),
    .X(_3021_));
 sky130_fd_sc_hd__o21a_1 _6335_ (.A1(\core_1.execute.alu_mul_div.div_res[13] ),
    .A2(_3021_),
    .B1(_1654_),
    .X(_0433_));
 sky130_fd_sc_hd__and3_1 _6336_ (.A(_1191_),
    .B(_1738_),
    .C(_3011_),
    .X(_3022_));
 sky130_fd_sc_hd__o21a_1 _6337_ (.A1(\core_1.execute.alu_mul_div.div_res[14] ),
    .A2(_3022_),
    .B1(_1654_),
    .X(_0434_));
 sky130_fd_sc_hd__a21oi_1 _6338_ (.A1(_1744_),
    .A2(_3011_),
    .B1(\core_1.execute.alu_mul_div.div_res[15] ),
    .Y(_3023_));
 sky130_fd_sc_hd__nor2_1 _6339_ (.A(_3005_),
    .B(_3023_),
    .Y(_0435_));
 sky130_fd_sc_hd__or2_1 _6340_ (.A(_1146_),
    .B(_1057_),
    .X(_3024_));
 sky130_fd_sc_hd__o221a_1 _6341_ (.A1(net194),
    .A2(_1309_),
    .B1(_2076_),
    .B2(_3024_),
    .C1(_2036_),
    .X(_3025_));
 sky130_fd_sc_hd__and2_2 _6342_ (.A(_1774_),
    .B(_1576_),
    .X(_3026_));
 sky130_fd_sc_hd__nor2_1 _6343_ (.A(net72),
    .B(_3026_),
    .Y(_3027_));
 sky130_fd_sc_hd__o21ai_1 _6344_ (.A1(_1577_),
    .A2(_3027_),
    .B1(_1307_),
    .Y(_3028_));
 sky130_fd_sc_hd__clkbuf_4 _6345_ (.A(_2819_),
    .X(_3029_));
 sky130_fd_sc_hd__o211a_1 _6346_ (.A1(_1307_),
    .A2(_3025_),
    .B1(_3028_),
    .C1(_3029_),
    .X(_0436_));
 sky130_fd_sc_hd__nor2_1 _6347_ (.A(net80),
    .B(_1578_),
    .Y(_3030_));
 sky130_fd_sc_hd__and3_1 _6348_ (.A(net80),
    .B(net79),
    .C(_1577_),
    .X(_3031_));
 sky130_fd_sc_hd__or3_1 _6349_ (.A(_1580_),
    .B(_3030_),
    .C(_3031_),
    .X(_3032_));
 sky130_fd_sc_hd__and2_1 _6350_ (.A(_1141_),
    .B(\core_1.dec_sreg_store ),
    .X(_3033_));
 sky130_fd_sc_hd__nand2_1 _6351_ (.A(_0643_),
    .B(_3033_),
    .Y(_3034_));
 sky130_fd_sc_hd__o2111ai_1 _6352_ (.A1(_3024_),
    .A2(_2131_),
    .B1(_2139_),
    .C1(_3034_),
    .D1(_1580_),
    .Y(_3035_));
 sky130_fd_sc_hd__a21oi_1 _6353_ (.A1(_3032_),
    .A2(_3035_),
    .B1(_1151_),
    .Y(_0437_));
 sky130_fd_sc_hd__clkbuf_4 _6354_ (.A(_1311_),
    .X(_3036_));
 sky130_fd_sc_hd__o21ai_1 _6355_ (.A1(_0635_),
    .A2(_1309_),
    .B1(_2153_),
    .Y(_3037_));
 sky130_fd_sc_hd__clkbuf_4 _6356_ (.A(_1306_),
    .X(_3038_));
 sky130_fd_sc_hd__a211o_1 _6357_ (.A1(_3036_),
    .A2(_2180_),
    .B1(_3037_),
    .C1(_3038_),
    .X(_3039_));
 sky130_fd_sc_hd__nor2_1 _6358_ (.A(net81),
    .B(_3031_),
    .Y(_3040_));
 sky130_fd_sc_hd__and3_1 _6359_ (.A(net80),
    .B(net72),
    .C(net79),
    .X(_3041_));
 sky130_fd_sc_hd__and3_1 _6360_ (.A(net81),
    .B(_3026_),
    .C(_3041_),
    .X(_3042_));
 sky130_fd_sc_hd__o21ai_1 _6361_ (.A1(_3040_),
    .A2(_3042_),
    .B1(_1307_),
    .Y(_3043_));
 sky130_fd_sc_hd__and3_1 _6362_ (.A(_3029_),
    .B(_3039_),
    .C(_3043_),
    .X(_3044_));
 sky130_fd_sc_hd__clkbuf_1 _6363_ (.A(_3044_),
    .X(_0438_));
 sky130_fd_sc_hd__o21ai_1 _6364_ (.A1(_0629_),
    .A2(_1309_),
    .B1(_2190_),
    .Y(_3045_));
 sky130_fd_sc_hd__a211o_1 _6365_ (.A1(_3036_),
    .A2(_2216_),
    .B1(_3045_),
    .C1(_3038_),
    .X(_3046_));
 sky130_fd_sc_hd__inv_2 _6366_ (.A(net82),
    .Y(_3047_));
 sky130_fd_sc_hd__o22ai_1 _6367_ (.A1(_1043_),
    .A2(_1305_),
    .B1(_3042_),
    .B2(_3047_),
    .Y(_3048_));
 sky130_fd_sc_hd__a21o_1 _6368_ (.A1(_3047_),
    .A2(_3042_),
    .B1(_3048_),
    .X(_3049_));
 sky130_fd_sc_hd__and3_1 _6369_ (.A(_3029_),
    .B(_3046_),
    .C(_3049_),
    .X(_3050_));
 sky130_fd_sc_hd__clkbuf_1 _6370_ (.A(_3050_),
    .X(_0439_));
 sky130_fd_sc_hd__a21oi_1 _6371_ (.A1(net82),
    .A2(_3042_),
    .B1(net83),
    .Y(_3051_));
 sky130_fd_sc_hd__and3_1 _6372_ (.A(net83),
    .B(net82),
    .C(_3042_),
    .X(_3052_));
 sky130_fd_sc_hd__o21ai_1 _6373_ (.A1(_3051_),
    .A2(_3052_),
    .B1(_1307_),
    .Y(_3053_));
 sky130_fd_sc_hd__o21ai_1 _6374_ (.A1(_0623_),
    .A2(_1308_),
    .B1(_2224_),
    .Y(_3054_));
 sky130_fd_sc_hd__a211o_1 _6375_ (.A1(_1311_),
    .A2(_2252_),
    .B1(_3054_),
    .C1(_1306_),
    .X(_3055_));
 sky130_fd_sc_hd__and3_1 _6376_ (.A(_3029_),
    .B(_3053_),
    .C(_3055_),
    .X(_3056_));
 sky130_fd_sc_hd__clkbuf_1 _6377_ (.A(_3056_),
    .X(_0440_));
 sky130_fd_sc_hd__o21ai_1 _6378_ (.A1(_0617_),
    .A2(_1309_),
    .B1(_2262_),
    .Y(_3057_));
 sky130_fd_sc_hd__a211o_1 _6379_ (.A1(_3036_),
    .A2(_2288_),
    .B1(_3057_),
    .C1(_3038_),
    .X(_3058_));
 sky130_fd_sc_hd__nor2_1 _6380_ (.A(net84),
    .B(_3052_),
    .Y(_3059_));
 sky130_fd_sc_hd__and2_1 _6381_ (.A(net84),
    .B(_3052_),
    .X(_3060_));
 sky130_fd_sc_hd__o21ai_1 _6382_ (.A1(_3059_),
    .A2(_3060_),
    .B1(_1307_),
    .Y(_3061_));
 sky130_fd_sc_hd__and3_1 _6383_ (.A(_3029_),
    .B(_3058_),
    .C(_3061_),
    .X(_3062_));
 sky130_fd_sc_hd__clkbuf_1 _6384_ (.A(_3062_),
    .X(_0441_));
 sky130_fd_sc_hd__o21ai_1 _6385_ (.A1(_0611_),
    .A2(_1309_),
    .B1(_2299_),
    .Y(_3063_));
 sky130_fd_sc_hd__a211o_1 _6386_ (.A1(_3036_),
    .A2(_2323_),
    .B1(_3063_),
    .C1(_3038_),
    .X(_3064_));
 sky130_fd_sc_hd__nor2_1 _6387_ (.A(net85),
    .B(_3060_),
    .Y(_3065_));
 sky130_fd_sc_hd__and3_2 _6388_ (.A(net85),
    .B(net84),
    .C(_3052_),
    .X(_3066_));
 sky130_fd_sc_hd__o21ai_1 _6389_ (.A1(_3065_),
    .A2(_3066_),
    .B1(_1307_),
    .Y(_3067_));
 sky130_fd_sc_hd__and3_1 _6390_ (.A(_3029_),
    .B(_3064_),
    .C(_3067_),
    .X(_3068_));
 sky130_fd_sc_hd__clkbuf_1 _6391_ (.A(_3068_),
    .X(_0442_));
 sky130_fd_sc_hd__o21ai_1 _6392_ (.A1(_0603_),
    .A2(_1309_),
    .B1(_2331_),
    .Y(_3069_));
 sky130_fd_sc_hd__a211o_1 _6393_ (.A1(_3036_),
    .A2(_2353_),
    .B1(_3069_),
    .C1(_3038_),
    .X(_3070_));
 sky130_fd_sc_hd__or2_1 _6394_ (.A(net86),
    .B(_3066_),
    .X(_3071_));
 sky130_fd_sc_hd__nand2_1 _6395_ (.A(net86),
    .B(_3066_),
    .Y(_3072_));
 sky130_fd_sc_hd__a21o_1 _6396_ (.A1(_3071_),
    .A2(_3072_),
    .B1(_1580_),
    .X(_3073_));
 sky130_fd_sc_hd__and3_1 _6397_ (.A(_2819_),
    .B(_3070_),
    .C(_3073_),
    .X(_3074_));
 sky130_fd_sc_hd__clkbuf_1 _6398_ (.A(_3074_),
    .X(_0443_));
 sky130_fd_sc_hd__o21ai_1 _6399_ (.A1(_0596_),
    .A2(_1309_),
    .B1(_2382_),
    .Y(_3075_));
 sky130_fd_sc_hd__a211o_1 _6400_ (.A1(_3036_),
    .A2(_2381_),
    .B1(_3075_),
    .C1(_3038_),
    .X(_3076_));
 sky130_fd_sc_hd__xor2_1 _6401_ (.A(net87),
    .B(_3072_),
    .X(_3077_));
 sky130_fd_sc_hd__nand2_1 _6402_ (.A(_1307_),
    .B(_3077_),
    .Y(_3078_));
 sky130_fd_sc_hd__and3_1 _6403_ (.A(_2819_),
    .B(_3076_),
    .C(_3078_),
    .X(_3079_));
 sky130_fd_sc_hd__clkbuf_1 _6404_ (.A(_3079_),
    .X(_0444_));
 sky130_fd_sc_hd__o21ai_1 _6405_ (.A1(_0588_),
    .A2(_1309_),
    .B1(_2395_),
    .Y(_3080_));
 sky130_fd_sc_hd__a211o_1 _6406_ (.A1(_3036_),
    .A2(_2419_),
    .B1(_3080_),
    .C1(_3038_),
    .X(_3081_));
 sky130_fd_sc_hd__a31oi_1 _6407_ (.A1(net87),
    .A2(net86),
    .A3(_3066_),
    .B1(net73),
    .Y(_3082_));
 sky130_fd_sc_hd__and4_1 _6408_ (.A(net73),
    .B(net87),
    .C(net86),
    .D(_3066_),
    .X(_3083_));
 sky130_fd_sc_hd__o21ai_1 _6409_ (.A1(_3082_),
    .A2(_3083_),
    .B1(_1307_),
    .Y(_3084_));
 sky130_fd_sc_hd__and3_1 _6410_ (.A(_2819_),
    .B(_3081_),
    .C(_3084_),
    .X(_3085_));
 sky130_fd_sc_hd__clkbuf_1 _6411_ (.A(_3085_),
    .X(_0445_));
 sky130_fd_sc_hd__o21ai_1 _6412_ (.A1(_0582_),
    .A2(_1309_),
    .B1(_2443_),
    .Y(_3086_));
 sky130_fd_sc_hd__a211o_1 _6413_ (.A1(_3036_),
    .A2(_2442_),
    .B1(_3086_),
    .C1(_3038_),
    .X(_3087_));
 sky130_fd_sc_hd__or2_1 _6414_ (.A(net74),
    .B(_3083_),
    .X(_3088_));
 sky130_fd_sc_hd__nand2_1 _6415_ (.A(net74),
    .B(_3083_),
    .Y(_3089_));
 sky130_fd_sc_hd__a21o_1 _6416_ (.A1(_3088_),
    .A2(_3089_),
    .B1(_1580_),
    .X(_3090_));
 sky130_fd_sc_hd__and3_1 _6417_ (.A(_2819_),
    .B(_3087_),
    .C(_3090_),
    .X(_3091_));
 sky130_fd_sc_hd__clkbuf_1 _6418_ (.A(_3091_),
    .X(_0446_));
 sky130_fd_sc_hd__o21ai_1 _6419_ (.A1(_0575_),
    .A2(_1308_),
    .B1(_2458_),
    .Y(_3092_));
 sky130_fd_sc_hd__a211o_1 _6420_ (.A1(_1311_),
    .A2(_2478_),
    .B1(_3092_),
    .C1(_3038_),
    .X(_3093_));
 sky130_fd_sc_hd__o22ai_1 _6421_ (.A1(_1043_),
    .A2(_1305_),
    .B1(_3089_),
    .B2(net75),
    .Y(_3094_));
 sky130_fd_sc_hd__a21o_1 _6422_ (.A1(net75),
    .A2(_3089_),
    .B1(_3094_),
    .X(_3095_));
 sky130_fd_sc_hd__and3_1 _6423_ (.A(_2819_),
    .B(_3093_),
    .C(_3095_),
    .X(_3096_));
 sky130_fd_sc_hd__clkbuf_1 _6424_ (.A(_3096_),
    .X(_0447_));
 sky130_fd_sc_hd__and3_1 _6425_ (.A(net82),
    .B(net81),
    .C(_3041_),
    .X(_3097_));
 sky130_fd_sc_hd__and3_1 _6426_ (.A(net86),
    .B(net85),
    .C(net84),
    .X(_3098_));
 sky130_fd_sc_hd__and3_1 _6427_ (.A(net75),
    .B(net74),
    .C(net83),
    .X(_3099_));
 sky130_fd_sc_hd__and4_1 _6428_ (.A(net73),
    .B(net87),
    .C(_3098_),
    .D(_3099_),
    .X(_3100_));
 sky130_fd_sc_hd__and3_1 _6429_ (.A(_3026_),
    .B(_3097_),
    .C(_3100_),
    .X(_3101_));
 sky130_fd_sc_hd__nor2_1 _6430_ (.A(net76),
    .B(_3101_),
    .Y(_3102_));
 sky130_fd_sc_hd__and2_1 _6431_ (.A(net76),
    .B(_3101_),
    .X(_3103_));
 sky130_fd_sc_hd__o21ai_1 _6432_ (.A1(_3102_),
    .A2(_3103_),
    .B1(_1307_),
    .Y(_3104_));
 sky130_fd_sc_hd__a221o_1 _6433_ (.A1(\core_1.execute.sreg_irq_pc.o_d[13] ),
    .A2(_1146_),
    .B1(net198),
    .B2(_3033_),
    .C1(_1306_),
    .X(_3105_));
 sky130_fd_sc_hd__a21o_1 _6434_ (.A1(_3036_),
    .A2(_2502_),
    .B1(_3105_),
    .X(_3106_));
 sky130_fd_sc_hd__and3_1 _6435_ (.A(_2819_),
    .B(_3104_),
    .C(_3106_),
    .X(_3107_));
 sky130_fd_sc_hd__clkbuf_1 _6436_ (.A(_3107_),
    .X(_0448_));
 sky130_fd_sc_hd__o21ai_1 _6437_ (.A1(_0553_),
    .A2(_1308_),
    .B1(_2519_),
    .Y(_3108_));
 sky130_fd_sc_hd__a211o_1 _6438_ (.A1(_1311_),
    .A2(_2538_),
    .B1(_3108_),
    .C1(_3038_),
    .X(_3109_));
 sky130_fd_sc_hd__or2_1 _6439_ (.A(net77),
    .B(_3103_),
    .X(_3110_));
 sky130_fd_sc_hd__nand2_1 _6440_ (.A(net77),
    .B(_3103_),
    .Y(_3111_));
 sky130_fd_sc_hd__a21o_1 _6441_ (.A1(_3110_),
    .A2(_3111_),
    .B1(_1580_),
    .X(_3112_));
 sky130_fd_sc_hd__and3_1 _6442_ (.A(_2819_),
    .B(_3109_),
    .C(_3112_),
    .X(_3113_));
 sky130_fd_sc_hd__clkbuf_1 _6443_ (.A(_3113_),
    .X(_0449_));
 sky130_fd_sc_hd__a21oi_1 _6444_ (.A1(net78),
    .A2(_3111_),
    .B1(_1580_),
    .Y(_3114_));
 sky130_fd_sc_hd__o21ai_1 _6445_ (.A1(net78),
    .A2(_3111_),
    .B1(_3114_),
    .Y(_3115_));
 sky130_fd_sc_hd__a221o_1 _6446_ (.A1(\core_1.execute.sreg_irq_pc.o_d[15] ),
    .A2(_1146_),
    .B1(net200),
    .B2(_3033_),
    .C1(_1306_),
    .X(_3116_));
 sky130_fd_sc_hd__a21o_1 _6447_ (.A1(_3036_),
    .A2(_2562_),
    .B1(_3116_),
    .X(_3117_));
 sky130_fd_sc_hd__and3_1 _6448_ (.A(_2819_),
    .B(_3115_),
    .C(_3117_),
    .X(_3118_));
 sky130_fd_sc_hd__clkbuf_1 _6449_ (.A(_3118_),
    .X(_0450_));
 sky130_fd_sc_hd__and2_2 _6450_ (.A(\core_1.dec_sreg_store ),
    .B(_2013_),
    .X(_3119_));
 sky130_fd_sc_hd__o21a_1 _6451_ (.A1(\core_1.dec_alu_flags_ie ),
    .A2(_3119_),
    .B1(_0734_),
    .X(_3120_));
 sky130_fd_sc_hd__buf_2 _6452_ (.A(_3120_),
    .X(_3121_));
 sky130_fd_sc_hd__nand2_2 _6453_ (.A(_1057_),
    .B(_2013_),
    .Y(_3122_));
 sky130_fd_sc_hd__a211o_1 _6454_ (.A1(_0780_),
    .A2(_2523_),
    .B1(_2533_),
    .C1(_2558_),
    .X(_3123_));
 sky130_fd_sc_hd__nand2_1 _6455_ (.A(_2475_),
    .B(_2499_),
    .Y(_3124_));
 sky130_fd_sc_hd__clkinv_2 _6456_ (.A(_2285_),
    .Y(_3125_));
 sky130_fd_sc_hd__nand2_1 _6457_ (.A(_2128_),
    .B(_2177_),
    .Y(_3126_));
 sky130_fd_sc_hd__or4_1 _6458_ (.A(_1570_),
    .B(_2071_),
    .C(_3126_),
    .D(_3119_),
    .X(_3127_));
 sky130_fd_sc_hd__inv_2 _6459_ (.A(_2249_),
    .Y(_3128_));
 sky130_fd_sc_hd__nand2_1 _6460_ (.A(_2213_),
    .B(_3128_),
    .Y(_3129_));
 sky130_fd_sc_hd__or4_1 _6461_ (.A(_3125_),
    .B(_2320_),
    .C(_3127_),
    .D(_3129_),
    .X(_3130_));
 sky130_fd_sc_hd__and2b_1 _6462_ (.A_N(_2416_),
    .B(_2439_),
    .X(_3131_));
 sky130_fd_sc_hd__and3_1 _6463_ (.A(_2350_),
    .B(_2378_),
    .C(_3131_),
    .X(_3132_));
 sky130_fd_sc_hd__or4b_1 _6464_ (.A(_3123_),
    .B(_3124_),
    .C(_3130_),
    .D_N(_3132_),
    .X(_3133_));
 sky130_fd_sc_hd__o211ai_1 _6465_ (.A1(_0658_),
    .A2(_3122_),
    .B1(_3133_),
    .C1(_3121_),
    .Y(_3134_));
 sky130_fd_sc_hd__o211a_1 _6466_ (.A1(\core_1.execute.alu_flag_reg.o_d[0] ),
    .A2(_3121_),
    .B1(_3134_),
    .C1(_2813_),
    .X(_0451_));
 sky130_fd_sc_hd__o21ai_1 _6467_ (.A1(_0650_),
    .A2(_3122_),
    .B1(_3121_),
    .Y(_3135_));
 sky130_fd_sc_hd__a21o_1 _6468_ (.A1(_1966_),
    .A2(_3122_),
    .B1(_3135_),
    .X(_3136_));
 sky130_fd_sc_hd__o211a_1 _6469_ (.A1(\core_1.execute.alu_flag_reg.o_d[1] ),
    .A2(_3121_),
    .B1(_3136_),
    .C1(_2813_),
    .X(_0452_));
 sky130_fd_sc_hd__o21ai_1 _6470_ (.A1(_0643_),
    .A2(_3122_),
    .B1(_3121_),
    .Y(_3137_));
 sky130_fd_sc_hd__a21o_1 _6471_ (.A1(_2558_),
    .A2(_3122_),
    .B1(_3137_),
    .X(_3138_));
 sky130_fd_sc_hd__o211a_1 _6472_ (.A1(\core_1.execute.alu_flag_reg.o_d[2] ),
    .A2(_3121_),
    .B1(_3138_),
    .C1(_2813_),
    .X(_0453_));
 sky130_fd_sc_hd__nand2_1 _6473_ (.A(_1733_),
    .B(_2558_),
    .Y(_3139_));
 sky130_fd_sc_hd__a21oi_1 _6474_ (.A1(_0863_),
    .A2(_2550_),
    .B1(_3119_),
    .Y(_3140_));
 sky130_fd_sc_hd__o221a_1 _6475_ (.A1(_0863_),
    .A2(_2550_),
    .B1(_2557_),
    .B2(_1733_),
    .C1(_3140_),
    .X(_3141_));
 sky130_fd_sc_hd__o21ai_1 _6476_ (.A1(_0635_),
    .A2(_3122_),
    .B1(_3121_),
    .Y(_3142_));
 sky130_fd_sc_hd__a21o_1 _6477_ (.A1(_3139_),
    .A2(_3141_),
    .B1(_3142_),
    .X(_3143_));
 sky130_fd_sc_hd__o211a_1 _6478_ (.A1(\core_1.execute.alu_flag_reg.o_d[3] ),
    .A2(_3121_),
    .B1(_3143_),
    .C1(_2813_),
    .X(_0454_));
 sky130_fd_sc_hd__o21ai_1 _6479_ (.A1(\core_1.execute.alu_flag_reg.o_d[4] ),
    .A2(_3121_),
    .B1(_1156_),
    .Y(_3144_));
 sky130_fd_sc_hd__or2_1 _6480_ (.A(_2128_),
    .B(_2177_),
    .X(_3145_));
 sky130_fd_sc_hd__and2_1 _6481_ (.A(_3126_),
    .B(_3145_),
    .X(_3146_));
 sky130_fd_sc_hd__xor2_1 _6482_ (.A(_1570_),
    .B(_2071_),
    .X(_3147_));
 sky130_fd_sc_hd__xnor2_1 _6483_ (.A(_3146_),
    .B(_3147_),
    .Y(_3148_));
 sky130_fd_sc_hd__xnor2_1 _6484_ (.A(_2213_),
    .B(_2249_),
    .Y(_3149_));
 sky130_fd_sc_hd__xnor2_1 _6485_ (.A(_3148_),
    .B(_3149_),
    .Y(_3150_));
 sky130_fd_sc_hd__xnor2_1 _6486_ (.A(_2416_),
    .B(_2439_),
    .Y(_3151_));
 sky130_fd_sc_hd__xnor2_1 _6487_ (.A(_2475_),
    .B(_2499_),
    .Y(_3152_));
 sky130_fd_sc_hd__xor2_1 _6488_ (.A(_2350_),
    .B(_2378_),
    .X(_3153_));
 sky130_fd_sc_hd__xnor2_1 _6489_ (.A(_3152_),
    .B(_3153_),
    .Y(_3154_));
 sky130_fd_sc_hd__xnor2_1 _6490_ (.A(_3151_),
    .B(_3154_),
    .Y(_3155_));
 sky130_fd_sc_hd__xnor2_1 _6491_ (.A(_3150_),
    .B(_3155_),
    .Y(_3156_));
 sky130_fd_sc_hd__xor2_1 _6492_ (.A(_2534_),
    .B(_2558_),
    .X(_3157_));
 sky130_fd_sc_hd__xnor2_1 _6493_ (.A(_2285_),
    .B(_2320_),
    .Y(_3158_));
 sky130_fd_sc_hd__xnor2_1 _6494_ (.A(_3157_),
    .B(_3158_),
    .Y(_3159_));
 sky130_fd_sc_hd__xnor2_1 _6495_ (.A(_3156_),
    .B(_3159_),
    .Y(_3160_));
 sky130_fd_sc_hd__nand2_1 _6496_ (.A(net204),
    .B(_3119_),
    .Y(_3161_));
 sky130_fd_sc_hd__o211a_1 _6497_ (.A1(_3119_),
    .A2(_3160_),
    .B1(_3161_),
    .C1(_3121_),
    .X(_3162_));
 sky130_fd_sc_hd__nor2_1 _6498_ (.A(_3144_),
    .B(_3162_),
    .Y(_0455_));
 sky130_fd_sc_hd__nand2_4 _6499_ (.A(_1057_),
    .B(_2294_),
    .Y(_3163_));
 sky130_fd_sc_hd__o21ai_4 _6500_ (.A1(_1777_),
    .A2(_3163_),
    .B1(_0668_),
    .Y(_3164_));
 sky130_fd_sc_hd__buf_4 _6501_ (.A(_3164_),
    .X(_3165_));
 sky130_fd_sc_hd__buf_4 _6502_ (.A(_3163_),
    .X(_3166_));
 sky130_fd_sc_hd__buf_4 _6503_ (.A(net37),
    .X(_3167_));
 sky130_fd_sc_hd__mux2_1 _6504_ (.A0(net72),
    .A1(\core_1.execute.mem_stage_pc[0] ),
    .S(_3167_),
    .X(_3168_));
 sky130_fd_sc_hd__buf_4 _6505_ (.A(_3163_),
    .X(_3169_));
 sky130_fd_sc_hd__nor2_1 _6506_ (.A(_0658_),
    .B(_3169_),
    .Y(_3170_));
 sky130_fd_sc_hd__o21a_2 _6507_ (.A1(_1777_),
    .A2(_3163_),
    .B1(_0668_),
    .X(_3171_));
 sky130_fd_sc_hd__buf_4 _6508_ (.A(_3171_),
    .X(_3172_));
 sky130_fd_sc_hd__a211o_1 _6509_ (.A1(_3166_),
    .A2(_3168_),
    .B1(_3170_),
    .C1(_3172_),
    .X(_3173_));
 sky130_fd_sc_hd__o211a_1 _6510_ (.A1(\core_1.execute.sreg_irq_pc.o_d[0] ),
    .A2(_3165_),
    .B1(_3173_),
    .C1(_2813_),
    .X(_0456_));
 sky130_fd_sc_hd__mux2_1 _6511_ (.A0(net79),
    .A1(\core_1.execute.mem_stage_pc[1] ),
    .S(_3167_),
    .X(_3174_));
 sky130_fd_sc_hd__nor2_1 _6512_ (.A(_0650_),
    .B(_3169_),
    .Y(_3175_));
 sky130_fd_sc_hd__a211o_1 _6513_ (.A1(_3166_),
    .A2(_3174_),
    .B1(_3175_),
    .C1(_3172_),
    .X(_3176_));
 sky130_fd_sc_hd__buf_4 _6514_ (.A(_1155_),
    .X(_3177_));
 sky130_fd_sc_hd__o211a_1 _6515_ (.A1(\core_1.execute.sreg_irq_pc.o_d[1] ),
    .A2(_3165_),
    .B1(_3176_),
    .C1(_3177_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_1 _6516_ (.A0(net80),
    .A1(\core_1.execute.mem_stage_pc[2] ),
    .S(_3167_),
    .X(_3178_));
 sky130_fd_sc_hd__nor2_1 _6517_ (.A(_0643_),
    .B(_3169_),
    .Y(_3179_));
 sky130_fd_sc_hd__a211o_1 _6518_ (.A1(_3166_),
    .A2(_3178_),
    .B1(_3179_),
    .C1(_3172_),
    .X(_3180_));
 sky130_fd_sc_hd__o211a_1 _6519_ (.A1(\core_1.execute.sreg_irq_pc.o_d[2] ),
    .A2(_3165_),
    .B1(_3180_),
    .C1(_3177_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_1 _6520_ (.A0(net81),
    .A1(\core_1.execute.mem_stage_pc[3] ),
    .S(_3167_),
    .X(_3181_));
 sky130_fd_sc_hd__nor2_1 _6521_ (.A(_0635_),
    .B(_3169_),
    .Y(_3182_));
 sky130_fd_sc_hd__a211o_1 _6522_ (.A1(_3166_),
    .A2(_3181_),
    .B1(_3182_),
    .C1(_3172_),
    .X(_3183_));
 sky130_fd_sc_hd__o211a_1 _6523_ (.A1(\core_1.execute.sreg_irq_pc.o_d[3] ),
    .A2(_3165_),
    .B1(_3183_),
    .C1(_3177_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_1 _6524_ (.A0(net82),
    .A1(\core_1.execute.mem_stage_pc[4] ),
    .S(_3167_),
    .X(_3184_));
 sky130_fd_sc_hd__buf_4 _6525_ (.A(_3163_),
    .X(_3185_));
 sky130_fd_sc_hd__nor2_1 _6526_ (.A(_0629_),
    .B(_3185_),
    .Y(_3186_));
 sky130_fd_sc_hd__a211o_1 _6527_ (.A1(_3166_),
    .A2(_3184_),
    .B1(_3186_),
    .C1(_3172_),
    .X(_3187_));
 sky130_fd_sc_hd__o211a_1 _6528_ (.A1(\core_1.execute.sreg_irq_pc.o_d[4] ),
    .A2(_3165_),
    .B1(_3187_),
    .C1(_3177_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_1 _6529_ (.A0(net83),
    .A1(\core_1.execute.mem_stage_pc[5] ),
    .S(_3167_),
    .X(_3188_));
 sky130_fd_sc_hd__nor2_1 _6530_ (.A(_0623_),
    .B(_3185_),
    .Y(_3189_));
 sky130_fd_sc_hd__a211o_1 _6531_ (.A1(_3166_),
    .A2(_3188_),
    .B1(_3189_),
    .C1(_3172_),
    .X(_3190_));
 sky130_fd_sc_hd__o211a_1 _6532_ (.A1(\core_1.execute.sreg_irq_pc.o_d[5] ),
    .A2(_3165_),
    .B1(_3190_),
    .C1(_3177_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_1 _6533_ (.A0(net84),
    .A1(\core_1.execute.mem_stage_pc[6] ),
    .S(_3167_),
    .X(_3191_));
 sky130_fd_sc_hd__nor2_1 _6534_ (.A(_0617_),
    .B(_3185_),
    .Y(_3192_));
 sky130_fd_sc_hd__a211o_1 _6535_ (.A1(_3166_),
    .A2(_3191_),
    .B1(_3192_),
    .C1(_3172_),
    .X(_3193_));
 sky130_fd_sc_hd__o211a_1 _6536_ (.A1(\core_1.execute.sreg_irq_pc.o_d[6] ),
    .A2(_3165_),
    .B1(_3193_),
    .C1(_3177_),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_1 _6537_ (.A0(net85),
    .A1(\core_1.execute.mem_stage_pc[7] ),
    .S(_3167_),
    .X(_3194_));
 sky130_fd_sc_hd__nor2_1 _6538_ (.A(_0611_),
    .B(_3185_),
    .Y(_3195_));
 sky130_fd_sc_hd__a211o_1 _6539_ (.A1(_3166_),
    .A2(_3194_),
    .B1(_3195_),
    .C1(_3172_),
    .X(_3196_));
 sky130_fd_sc_hd__o211a_1 _6540_ (.A1(\core_1.execute.sreg_irq_pc.o_d[7] ),
    .A2(_3165_),
    .B1(_3196_),
    .C1(_3177_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_1 _6541_ (.A0(net86),
    .A1(\core_1.execute.mem_stage_pc[8] ),
    .S(_3167_),
    .X(_3197_));
 sky130_fd_sc_hd__nor2_1 _6542_ (.A(_0603_),
    .B(_3185_),
    .Y(_3198_));
 sky130_fd_sc_hd__a211o_1 _6543_ (.A1(_3166_),
    .A2(_3197_),
    .B1(_3198_),
    .C1(_3172_),
    .X(_3199_));
 sky130_fd_sc_hd__o211a_1 _6544_ (.A1(\core_1.execute.sreg_irq_pc.o_d[8] ),
    .A2(_3165_),
    .B1(_3199_),
    .C1(_3177_),
    .X(_0464_));
 sky130_fd_sc_hd__mux2_1 _6545_ (.A0(net87),
    .A1(\core_1.execute.mem_stage_pc[9] ),
    .S(net37),
    .X(_3200_));
 sky130_fd_sc_hd__nor2_1 _6546_ (.A(_0596_),
    .B(_3185_),
    .Y(_3201_));
 sky130_fd_sc_hd__a211o_1 _6547_ (.A1(_3166_),
    .A2(_3200_),
    .B1(_3201_),
    .C1(_3172_),
    .X(_3202_));
 sky130_fd_sc_hd__o211a_1 _6548_ (.A1(\core_1.execute.sreg_irq_pc.o_d[9] ),
    .A2(_3165_),
    .B1(_3202_),
    .C1(_3177_),
    .X(_0465_));
 sky130_fd_sc_hd__mux2_1 _6549_ (.A0(net73),
    .A1(\core_1.execute.mem_stage_pc[10] ),
    .S(net37),
    .X(_3203_));
 sky130_fd_sc_hd__nor2_1 _6550_ (.A(_0588_),
    .B(_3185_),
    .Y(_3204_));
 sky130_fd_sc_hd__a211o_1 _6551_ (.A1(_3169_),
    .A2(_3203_),
    .B1(_3204_),
    .C1(_3171_),
    .X(_3205_));
 sky130_fd_sc_hd__o211a_1 _6552_ (.A1(\core_1.execute.sreg_irq_pc.o_d[10] ),
    .A2(_3164_),
    .B1(_3205_),
    .C1(_3177_),
    .X(_0466_));
 sky130_fd_sc_hd__mux2_1 _6553_ (.A0(net74),
    .A1(\core_1.execute.mem_stage_pc[11] ),
    .S(net37),
    .X(_3206_));
 sky130_fd_sc_hd__nor2_1 _6554_ (.A(_0582_),
    .B(_3185_),
    .Y(_3207_));
 sky130_fd_sc_hd__a211o_1 _6555_ (.A1(_3169_),
    .A2(_3206_),
    .B1(_3207_),
    .C1(_3171_),
    .X(_3208_));
 sky130_fd_sc_hd__clkbuf_8 _6556_ (.A(_1155_),
    .X(_3209_));
 sky130_fd_sc_hd__o211a_1 _6557_ (.A1(\core_1.execute.sreg_irq_pc.o_d[11] ),
    .A2(_3164_),
    .B1(_3208_),
    .C1(_3209_),
    .X(_0467_));
 sky130_fd_sc_hd__mux2_1 _6558_ (.A0(net75),
    .A1(\core_1.execute.mem_stage_pc[12] ),
    .S(net37),
    .X(_3210_));
 sky130_fd_sc_hd__nor2_1 _6559_ (.A(_0575_),
    .B(_3185_),
    .Y(_3211_));
 sky130_fd_sc_hd__a211o_1 _6560_ (.A1(_3169_),
    .A2(_3210_),
    .B1(_3211_),
    .C1(_3171_),
    .X(_3212_));
 sky130_fd_sc_hd__o211a_1 _6561_ (.A1(\core_1.execute.sreg_irq_pc.o_d[12] ),
    .A2(_3164_),
    .B1(_3212_),
    .C1(_3209_),
    .X(_0468_));
 sky130_fd_sc_hd__mux2_1 _6562_ (.A0(net76),
    .A1(\core_1.execute.mem_stage_pc[13] ),
    .S(net37),
    .X(_3213_));
 sky130_fd_sc_hd__nor2_1 _6563_ (.A(_0568_),
    .B(_3185_),
    .Y(_3214_));
 sky130_fd_sc_hd__a211o_1 _6564_ (.A1(_3169_),
    .A2(_3213_),
    .B1(_3214_),
    .C1(_3171_),
    .X(_3215_));
 sky130_fd_sc_hd__o211a_1 _6565_ (.A1(\core_1.execute.sreg_irq_pc.o_d[13] ),
    .A2(_3164_),
    .B1(_3215_),
    .C1(_3209_),
    .X(_0469_));
 sky130_fd_sc_hd__mux2_1 _6566_ (.A0(net77),
    .A1(\core_1.execute.mem_stage_pc[14] ),
    .S(net37),
    .X(_3216_));
 sky130_fd_sc_hd__nor2_1 _6567_ (.A(_0553_),
    .B(_3163_),
    .Y(_3217_));
 sky130_fd_sc_hd__a211o_1 _6568_ (.A1(_3169_),
    .A2(_3216_),
    .B1(_3217_),
    .C1(_3171_),
    .X(_3218_));
 sky130_fd_sc_hd__o211a_1 _6569_ (.A1(\core_1.execute.sreg_irq_pc.o_d[14] ),
    .A2(_3164_),
    .B1(_3218_),
    .C1(_3209_),
    .X(_0470_));
 sky130_fd_sc_hd__mux2_1 _6570_ (.A0(net78),
    .A1(\core_1.execute.mem_stage_pc[15] ),
    .S(net37),
    .X(_3219_));
 sky130_fd_sc_hd__nor2_1 _6571_ (.A(_0545_),
    .B(_3163_),
    .Y(_3220_));
 sky130_fd_sc_hd__a211o_1 _6572_ (.A1(_3169_),
    .A2(_3219_),
    .B1(_3220_),
    .C1(_3171_),
    .X(_3221_));
 sky130_fd_sc_hd__o211a_1 _6573_ (.A1(\core_1.execute.sreg_irq_pc.o_d[15] ),
    .A2(_3164_),
    .B1(_3221_),
    .C1(_3209_),
    .X(_0471_));
 sky130_fd_sc_hd__and4_1 _6574_ (.A(\core_1.execute.sreg_priv_control.o_d[0] ),
    .B(_1057_),
    .C(_0668_),
    .D(_2027_),
    .X(_3222_));
 sky130_fd_sc_hd__a31oi_4 _6575_ (.A1(\core_1.execute.sreg_priv_control.o_d[0] ),
    .A2(_1057_),
    .A3(_2027_),
    .B1(_0667_),
    .Y(_3223_));
 sky130_fd_sc_hd__a22o_1 _6576_ (.A1(net194),
    .A2(_3222_),
    .B1(_3223_),
    .B2(\core_1.execute.sreg_jtr_buff.o_d[0] ),
    .X(_3224_));
 sky130_fd_sc_hd__and2_1 _6577_ (.A(_1178_),
    .B(_3224_),
    .X(_3225_));
 sky130_fd_sc_hd__clkbuf_1 _6578_ (.A(_3225_),
    .X(_0472_));
 sky130_fd_sc_hd__a22o_1 _6579_ (.A1(net201),
    .A2(_3222_),
    .B1(_3223_),
    .B2(\core_1.execute.sreg_jtr_buff.o_d[1] ),
    .X(_3226_));
 sky130_fd_sc_hd__and2_1 _6580_ (.A(_1178_),
    .B(_3226_),
    .X(_3227_));
 sky130_fd_sc_hd__clkbuf_1 _6581_ (.A(_3227_),
    .X(_0473_));
 sky130_fd_sc_hd__a22o_1 _6582_ (.A1(net202),
    .A2(_3222_),
    .B1(_3223_),
    .B2(\core_1.execute.sreg_jtr_buff.o_d[2] ),
    .X(_3228_));
 sky130_fd_sc_hd__and2_1 _6583_ (.A(_1178_),
    .B(_3228_),
    .X(_3229_));
 sky130_fd_sc_hd__clkbuf_1 _6584_ (.A(_3229_),
    .X(_0474_));
 sky130_fd_sc_hd__nand2_1 _6585_ (.A(net106),
    .B(_1048_),
    .Y(_3230_));
 sky130_fd_sc_hd__a21oi_1 _6586_ (.A1(_1046_),
    .A2(_3230_),
    .B1(_1165_),
    .Y(_0475_));
 sky130_fd_sc_hd__a22o_1 _6587_ (.A1(\core_1.execute.sreg_jtr_buff.o_d[1] ),
    .A2(_1047_),
    .B1(_1048_),
    .B2(\core_1.execute.trap_flag ),
    .X(_3231_));
 sky130_fd_sc_hd__and2_1 _6588_ (.A(_1178_),
    .B(_3231_),
    .X(_3232_));
 sky130_fd_sc_hd__clkbuf_1 _6589_ (.A(_3232_),
    .X(_0476_));
 sky130_fd_sc_hd__a22o_1 _6590_ (.A1(\core_1.execute.sreg_jtr_buff.o_d[2] ),
    .A2(_1047_),
    .B1(_1048_),
    .B2(_0670_),
    .X(_3233_));
 sky130_fd_sc_hd__and2_1 _6591_ (.A(_1178_),
    .B(_3233_),
    .X(_3234_));
 sky130_fd_sc_hd__clkbuf_1 _6592_ (.A(_3234_),
    .X(_0477_));
 sky130_fd_sc_hd__and3_1 _6593_ (.A(_1057_),
    .B(_1774_),
    .C(_2293_),
    .X(_3235_));
 sky130_fd_sc_hd__clkbuf_2 _6594_ (.A(_3235_),
    .X(_3236_));
 sky130_fd_sc_hd__clkbuf_4 _6595_ (.A(_3236_),
    .X(_3237_));
 sky130_fd_sc_hd__buf_4 _6596_ (.A(_3236_),
    .X(_3238_));
 sky130_fd_sc_hd__clkbuf_4 _6597_ (.A(_0659_),
    .X(_3239_));
 sky130_fd_sc_hd__a21oi_1 _6598_ (.A1(_0658_),
    .A2(_3238_),
    .B1(_3239_),
    .Y(_3240_));
 sky130_fd_sc_hd__o21a_1 _6599_ (.A1(\core_1.execute.sreg_scratch.o_d[0] ),
    .A2(_3237_),
    .B1(_3240_),
    .X(_0478_));
 sky130_fd_sc_hd__a21oi_1 _6600_ (.A1(_0650_),
    .A2(_3238_),
    .B1(_3239_),
    .Y(_3241_));
 sky130_fd_sc_hd__o21a_1 _6601_ (.A1(\core_1.execute.sreg_scratch.o_d[1] ),
    .A2(_3237_),
    .B1(_3241_),
    .X(_0479_));
 sky130_fd_sc_hd__a21oi_1 _6602_ (.A1(_0643_),
    .A2(_3238_),
    .B1(_3239_),
    .Y(_3242_));
 sky130_fd_sc_hd__o21a_1 _6603_ (.A1(\core_1.execute.sreg_scratch.o_d[2] ),
    .A2(_3237_),
    .B1(_3242_),
    .X(_0480_));
 sky130_fd_sc_hd__a21oi_1 _6604_ (.A1(_0635_),
    .A2(_3238_),
    .B1(_3239_),
    .Y(_3243_));
 sky130_fd_sc_hd__o21a_1 _6605_ (.A1(\core_1.execute.sreg_scratch.o_d[3] ),
    .A2(_3237_),
    .B1(_3243_),
    .X(_0481_));
 sky130_fd_sc_hd__buf_4 _6606_ (.A(_3236_),
    .X(_3244_));
 sky130_fd_sc_hd__a21oi_1 _6607_ (.A1(_0629_),
    .A2(_3244_),
    .B1(_3239_),
    .Y(_3245_));
 sky130_fd_sc_hd__o21a_1 _6608_ (.A1(\core_1.execute.sreg_scratch.o_d[4] ),
    .A2(_3237_),
    .B1(_3245_),
    .X(_0482_));
 sky130_fd_sc_hd__a21oi_1 _6609_ (.A1(_0623_),
    .A2(_3244_),
    .B1(_3239_),
    .Y(_3246_));
 sky130_fd_sc_hd__o21a_1 _6610_ (.A1(\core_1.execute.sreg_scratch.o_d[5] ),
    .A2(_3237_),
    .B1(_3246_),
    .X(_0483_));
 sky130_fd_sc_hd__a21oi_1 _6611_ (.A1(_0617_),
    .A2(_3244_),
    .B1(_3239_),
    .Y(_3247_));
 sky130_fd_sc_hd__o21a_1 _6612_ (.A1(\core_1.execute.sreg_scratch.o_d[6] ),
    .A2(_3237_),
    .B1(_3247_),
    .X(_0484_));
 sky130_fd_sc_hd__a21oi_1 _6613_ (.A1(_0611_),
    .A2(_3244_),
    .B1(_3239_),
    .Y(_3248_));
 sky130_fd_sc_hd__o21a_1 _6614_ (.A1(\core_1.execute.sreg_scratch.o_d[7] ),
    .A2(_3237_),
    .B1(_3248_),
    .X(_0485_));
 sky130_fd_sc_hd__a21oi_1 _6615_ (.A1(_0603_),
    .A2(_3244_),
    .B1(_3239_),
    .Y(_3249_));
 sky130_fd_sc_hd__o21a_1 _6616_ (.A1(\core_1.execute.sreg_scratch.o_d[8] ),
    .A2(_3237_),
    .B1(_3249_),
    .X(_0486_));
 sky130_fd_sc_hd__a21oi_1 _6617_ (.A1(_0596_),
    .A2(_3244_),
    .B1(_1055_),
    .Y(_3250_));
 sky130_fd_sc_hd__o21a_1 _6618_ (.A1(\core_1.execute.sreg_scratch.o_d[9] ),
    .A2(_3237_),
    .B1(_3250_),
    .X(_0487_));
 sky130_fd_sc_hd__a21oi_1 _6619_ (.A1(_0588_),
    .A2(_3244_),
    .B1(_1055_),
    .Y(_3251_));
 sky130_fd_sc_hd__o21a_1 _6620_ (.A1(\core_1.execute.sreg_scratch.o_d[10] ),
    .A2(_3238_),
    .B1(_3251_),
    .X(_0488_));
 sky130_fd_sc_hd__a21oi_1 _6621_ (.A1(_0582_),
    .A2(_3244_),
    .B1(_1055_),
    .Y(_3252_));
 sky130_fd_sc_hd__o21a_1 _6622_ (.A1(\core_1.execute.sreg_scratch.o_d[11] ),
    .A2(_3238_),
    .B1(_3252_),
    .X(_0489_));
 sky130_fd_sc_hd__a21oi_1 _6623_ (.A1(_0575_),
    .A2(_3244_),
    .B1(_1055_),
    .Y(_3253_));
 sky130_fd_sc_hd__o21a_1 _6624_ (.A1(\core_1.execute.sreg_scratch.o_d[12] ),
    .A2(_3238_),
    .B1(_3253_),
    .X(_0490_));
 sky130_fd_sc_hd__a21oi_1 _6625_ (.A1(_0568_),
    .A2(_3244_),
    .B1(_1055_),
    .Y(_3254_));
 sky130_fd_sc_hd__o21a_1 _6626_ (.A1(\core_1.execute.sreg_scratch.o_d[13] ),
    .A2(_3238_),
    .B1(_3254_),
    .X(_0491_));
 sky130_fd_sc_hd__a21oi_1 _6627_ (.A1(_0553_),
    .A2(_3236_),
    .B1(_1055_),
    .Y(_3255_));
 sky130_fd_sc_hd__o21a_1 _6628_ (.A1(\core_1.execute.sreg_scratch.o_d[14] ),
    .A2(_3238_),
    .B1(_3255_),
    .X(_0492_));
 sky130_fd_sc_hd__a21oi_1 _6629_ (.A1(_0545_),
    .A2(_3236_),
    .B1(_1055_),
    .Y(_3256_));
 sky130_fd_sc_hd__o21a_1 _6630_ (.A1(\core_1.execute.sreg_scratch.o_d[15] ),
    .A2(_3238_),
    .B1(_3256_),
    .X(_0493_));
 sky130_fd_sc_hd__clkbuf_4 _6631_ (.A(_1155_),
    .X(_3257_));
 sky130_fd_sc_hd__a32o_1 _6632_ (.A1(\core_1.execute.irq_en ),
    .A2(net18),
    .A3(_3257_),
    .B1(_3029_),
    .B2(\core_1.execute.sreg_irq_flags.o_d[0] ),
    .X(_0494_));
 sky130_fd_sc_hd__inv_2 _6633_ (.A(\core_1.execute.sreg_irq_flags.o_d[1] ),
    .Y(_3258_));
 sky130_fd_sc_hd__nor2_1 _6634_ (.A(_3258_),
    .B(_0666_),
    .Y(_3259_));
 sky130_fd_sc_hd__o21a_1 _6635_ (.A1(\core_1.execute.prev_sys ),
    .A2(_3259_),
    .B1(_1776_),
    .X(_0495_));
 sky130_fd_sc_hd__a22o_1 _6636_ (.A1(\core_1.execute.sreg_irq_flags.i_d[2] ),
    .A2(_3257_),
    .B1(_3029_),
    .B2(\core_1.execute.sreg_irq_flags.o_d[2] ),
    .X(_0496_));
 sky130_fd_sc_hd__a22o_1 _6637_ (.A1(_3167_),
    .A2(_3257_),
    .B1(_3029_),
    .B2(\core_1.execute.sreg_irq_flags.o_d[3] ),
    .X(_0497_));
 sky130_fd_sc_hd__a32o_1 _6638_ (.A1(\core_1.execute.irq_en ),
    .A2(net19),
    .A3(_3257_),
    .B1(_3029_),
    .B2(\core_1.execute.sreg_irq_flags.o_d[4] ),
    .X(_0498_));
 sky130_fd_sc_hd__and2_1 _6639_ (.A(\core_1.dec_sreg_store ),
    .B(_2024_),
    .X(_3260_));
 sky130_fd_sc_hd__clkbuf_4 _6640_ (.A(_3260_),
    .X(_3261_));
 sky130_fd_sc_hd__and2_1 _6641_ (.A(_0670_),
    .B(_1045_),
    .X(_3262_));
 sky130_fd_sc_hd__a31o_1 _6642_ (.A1(_0670_),
    .A2(net77),
    .A3(_3026_),
    .B1(_3262_),
    .X(_3263_));
 sky130_fd_sc_hd__o21a_4 _6643_ (.A1(_3261_),
    .A2(_3263_),
    .B1(_1774_),
    .X(_3264_));
 sky130_fd_sc_hd__clkinv_2 _6644_ (.A(_3264_),
    .Y(_3265_));
 sky130_fd_sc_hd__nand2_1 _6645_ (.A(_0670_),
    .B(_1045_),
    .Y(_3266_));
 sky130_fd_sc_hd__buf_2 _6646_ (.A(_3266_),
    .X(_3267_));
 sky130_fd_sc_hd__nand2_1 _6647_ (.A(\core_1.execute.pc_high_out[0] ),
    .B(_3266_),
    .Y(_3268_));
 sky130_fd_sc_hd__nand2_4 _6648_ (.A(_1057_),
    .B(_2024_),
    .Y(_3269_));
 sky130_fd_sc_hd__o211a_1 _6649_ (.A1(\core_1.execute.pc_high_buff_out[0] ),
    .A2(_3267_),
    .B1(_3268_),
    .C1(_3269_),
    .X(_3270_));
 sky130_fd_sc_hd__a211o_1 _6650_ (.A1(net194),
    .A2(_3261_),
    .B1(_3265_),
    .C1(_3270_),
    .X(_3271_));
 sky130_fd_sc_hd__o211a_1 _6651_ (.A1(\core_1.execute.pc_high_out[0] ),
    .A2(_3264_),
    .B1(_3271_),
    .C1(_3209_),
    .X(_0499_));
 sky130_fd_sc_hd__nand2_1 _6652_ (.A(\core_1.execute.pc_high_out[1] ),
    .B(\core_1.execute.pc_high_out[0] ),
    .Y(_3272_));
 sky130_fd_sc_hd__or2_1 _6653_ (.A(\core_1.execute.pc_high_out[1] ),
    .B(\core_1.execute.pc_high_out[0] ),
    .X(_3273_));
 sky130_fd_sc_hd__and3_1 _6654_ (.A(_3266_),
    .B(_3272_),
    .C(_3273_),
    .X(_3274_));
 sky130_fd_sc_hd__a211o_1 _6655_ (.A1(\core_1.execute.pc_high_buff_out[1] ),
    .A2(_3262_),
    .B1(_3274_),
    .C1(_3261_),
    .X(_3275_));
 sky130_fd_sc_hd__o21ai_1 _6656_ (.A1(net201),
    .A2(_3269_),
    .B1(_3275_),
    .Y(_3276_));
 sky130_fd_sc_hd__nand2_1 _6657_ (.A(_3264_),
    .B(_3276_),
    .Y(_3277_));
 sky130_fd_sc_hd__o211a_1 _6658_ (.A1(\core_1.execute.pc_high_out[1] ),
    .A2(_3264_),
    .B1(_3277_),
    .C1(_3209_),
    .X(_0500_));
 sky130_fd_sc_hd__inv_2 _6659_ (.A(\core_1.execute.pc_high_out[2] ),
    .Y(_3278_));
 sky130_fd_sc_hd__xnor2_1 _6660_ (.A(_3278_),
    .B(_3272_),
    .Y(_3279_));
 sky130_fd_sc_hd__a21o_1 _6661_ (.A1(_3267_),
    .A2(_3279_),
    .B1(_3261_),
    .X(_3280_));
 sky130_fd_sc_hd__nor2_1 _6662_ (.A(\core_1.execute.pc_high_buff_out[2] ),
    .B(_3267_),
    .Y(_3281_));
 sky130_fd_sc_hd__o221a_1 _6663_ (.A1(_0643_),
    .A2(_3269_),
    .B1(_3280_),
    .B2(_3281_),
    .C1(_3264_),
    .X(_3282_));
 sky130_fd_sc_hd__a211oi_1 _6664_ (.A1(_3278_),
    .A2(_3265_),
    .B1(_3282_),
    .C1(_1165_),
    .Y(_0501_));
 sky130_fd_sc_hd__and4_1 _6665_ (.A(\core_1.execute.pc_high_out[3] ),
    .B(\core_1.execute.pc_high_out[2] ),
    .C(\core_1.execute.pc_high_out[1] ),
    .D(\core_1.execute.pc_high_out[0] ),
    .X(_3283_));
 sky130_fd_sc_hd__o21ba_1 _6666_ (.A1(_3278_),
    .A2(_3272_),
    .B1_N(\core_1.execute.pc_high_out[3] ),
    .X(_3284_));
 sky130_fd_sc_hd__o21ai_1 _6667_ (.A1(_3283_),
    .A2(_3284_),
    .B1(_3267_),
    .Y(_3285_));
 sky130_fd_sc_hd__o211a_1 _6668_ (.A1(\core_1.execute.pc_high_buff_out[3] ),
    .A2(_3267_),
    .B1(_3285_),
    .C1(_3269_),
    .X(_3286_));
 sky130_fd_sc_hd__a211o_1 _6669_ (.A1(net203),
    .A2(_3261_),
    .B1(_3265_),
    .C1(_3286_),
    .X(_3287_));
 sky130_fd_sc_hd__o211a_1 _6670_ (.A1(\core_1.execute.pc_high_out[3] ),
    .A2(_3264_),
    .B1(_3287_),
    .C1(_3209_),
    .X(_0502_));
 sky130_fd_sc_hd__inv_2 _6671_ (.A(\core_1.execute.pc_high_out[4] ),
    .Y(_3288_));
 sky130_fd_sc_hd__xnor2_1 _6672_ (.A(\core_1.execute.pc_high_out[4] ),
    .B(_3283_),
    .Y(_3289_));
 sky130_fd_sc_hd__a21o_1 _6673_ (.A1(_3267_),
    .A2(_3289_),
    .B1(_3261_),
    .X(_3290_));
 sky130_fd_sc_hd__nor2_1 _6674_ (.A(\core_1.execute.pc_high_buff_out[4] ),
    .B(_3267_),
    .Y(_3291_));
 sky130_fd_sc_hd__o221a_1 _6675_ (.A1(_0629_),
    .A2(_3269_),
    .B1(_3290_),
    .B2(_3291_),
    .C1(_3264_),
    .X(_3292_));
 sky130_fd_sc_hd__a211oi_1 _6676_ (.A1(_3288_),
    .A2(_3265_),
    .B1(_3292_),
    .C1(_1165_),
    .Y(_0503_));
 sky130_fd_sc_hd__and3_1 _6677_ (.A(\core_1.execute.pc_high_out[5] ),
    .B(\core_1.execute.pc_high_out[4] ),
    .C(_3283_),
    .X(_3293_));
 sky130_fd_sc_hd__a21oi_1 _6678_ (.A1(\core_1.execute.pc_high_out[4] ),
    .A2(_3283_),
    .B1(\core_1.execute.pc_high_out[5] ),
    .Y(_3294_));
 sky130_fd_sc_hd__o21ai_1 _6679_ (.A1(_3293_),
    .A2(_3294_),
    .B1(_3266_),
    .Y(_3295_));
 sky130_fd_sc_hd__o211a_1 _6680_ (.A1(\core_1.execute.pc_high_buff_out[5] ),
    .A2(_3267_),
    .B1(_3295_),
    .C1(_3269_),
    .X(_3296_));
 sky130_fd_sc_hd__a211o_1 _6681_ (.A1(net205),
    .A2(_3261_),
    .B1(_3265_),
    .C1(_3296_),
    .X(_3297_));
 sky130_fd_sc_hd__o211a_1 _6682_ (.A1(\core_1.execute.pc_high_out[5] ),
    .A2(_3264_),
    .B1(_3297_),
    .C1(_3209_),
    .X(_0504_));
 sky130_fd_sc_hd__inv_2 _6683_ (.A(\core_1.execute.pc_high_out[6] ),
    .Y(_3298_));
 sky130_fd_sc_hd__nand2_1 _6684_ (.A(\core_1.execute.pc_high_out[6] ),
    .B(_3293_),
    .Y(_3299_));
 sky130_fd_sc_hd__or2_1 _6685_ (.A(\core_1.execute.pc_high_out[6] ),
    .B(_3293_),
    .X(_3300_));
 sky130_fd_sc_hd__nand2_1 _6686_ (.A(_3299_),
    .B(_3300_),
    .Y(_3301_));
 sky130_fd_sc_hd__a21o_1 _6687_ (.A1(_3267_),
    .A2(_3301_),
    .B1(_3261_),
    .X(_3302_));
 sky130_fd_sc_hd__nor2_1 _6688_ (.A(\core_1.execute.pc_high_buff_out[6] ),
    .B(_3267_),
    .Y(_3303_));
 sky130_fd_sc_hd__o221a_1 _6689_ (.A1(_0617_),
    .A2(_3269_),
    .B1(_3302_),
    .B2(_3303_),
    .C1(_3264_),
    .X(_3304_));
 sky130_fd_sc_hd__a211oi_1 _6690_ (.A1(_3298_),
    .A2(_3265_),
    .B1(_3304_),
    .C1(_3239_),
    .Y(_0505_));
 sky130_fd_sc_hd__xor2_1 _6691_ (.A(\core_1.execute.pc_high_out[7] ),
    .B(_3299_),
    .X(_3305_));
 sky130_fd_sc_hd__nor2_1 _6692_ (.A(_3262_),
    .B(_3305_),
    .Y(_3306_));
 sky130_fd_sc_hd__a211o_1 _6693_ (.A1(\core_1.execute.pc_high_buff_out[7] ),
    .A2(_3262_),
    .B1(_3306_),
    .C1(_3261_),
    .X(_3307_));
 sky130_fd_sc_hd__o211a_1 _6694_ (.A1(net207),
    .A2(_3269_),
    .B1(_3264_),
    .C1(_3307_),
    .X(_3308_));
 sky130_fd_sc_hd__a211o_1 _6695_ (.A1(\core_1.execute.pc_high_out[7] ),
    .A2(_3265_),
    .B1(_3308_),
    .C1(_1165_),
    .X(_0506_));
 sky130_fd_sc_hd__and2_1 _6696_ (.A(\core_1.dec_sreg_store ),
    .B(_2032_),
    .X(_3309_));
 sky130_fd_sc_hd__buf_2 _6697_ (.A(_3309_),
    .X(_3310_));
 sky130_fd_sc_hd__a21oi_1 _6698_ (.A1(_0670_),
    .A2(\core_1.dec_sreg_jal_over ),
    .B1(_3310_),
    .Y(_3311_));
 sky130_fd_sc_hd__nor2_4 _6699_ (.A(_1777_),
    .B(_3311_),
    .Y(_3312_));
 sky130_fd_sc_hd__buf_2 _6700_ (.A(_3310_),
    .X(_3313_));
 sky130_fd_sc_hd__clkinv_2 _6701_ (.A(_3312_),
    .Y(_3314_));
 sky130_fd_sc_hd__nor2_1 _6702_ (.A(_0684_),
    .B(_3313_),
    .Y(_3315_));
 sky130_fd_sc_hd__a211o_1 _6703_ (.A1(net194),
    .A2(_3313_),
    .B1(_3314_),
    .C1(_3315_),
    .X(_3316_));
 sky130_fd_sc_hd__o211a_1 _6704_ (.A1(\core_1.execute.pc_high_buff_out[0] ),
    .A2(_3312_),
    .B1(_3316_),
    .C1(_3209_),
    .X(_0507_));
 sky130_fd_sc_hd__nor2_1 _6705_ (.A(_0674_),
    .B(_3313_),
    .Y(_3317_));
 sky130_fd_sc_hd__a211o_1 _6706_ (.A1(net201),
    .A2(_3313_),
    .B1(_3314_),
    .C1(_3317_),
    .X(_3318_));
 sky130_fd_sc_hd__o211a_1 _6707_ (.A1(\core_1.execute.pc_high_buff_out[1] ),
    .A2(_3312_),
    .B1(_3318_),
    .C1(_3257_),
    .X(_0508_));
 sky130_fd_sc_hd__nor2_1 _6708_ (.A(_0672_),
    .B(_3310_),
    .Y(_3319_));
 sky130_fd_sc_hd__a211o_1 _6709_ (.A1(net202),
    .A2(_3313_),
    .B1(_3314_),
    .C1(_3319_),
    .X(_3320_));
 sky130_fd_sc_hd__o211a_1 _6710_ (.A1(\core_1.execute.pc_high_buff_out[2] ),
    .A2(_3312_),
    .B1(_3320_),
    .C1(_3257_),
    .X(_0509_));
 sky130_fd_sc_hd__nor2_1 _6711_ (.A(_0669_),
    .B(_3310_),
    .Y(_3321_));
 sky130_fd_sc_hd__a211o_1 _6712_ (.A1(net203),
    .A2(_3313_),
    .B1(_3314_),
    .C1(_3321_),
    .X(_3322_));
 sky130_fd_sc_hd__o211a_1 _6713_ (.A1(\core_1.execute.pc_high_buff_out[3] ),
    .A2(_3312_),
    .B1(_3322_),
    .C1(_3257_),
    .X(_0510_));
 sky130_fd_sc_hd__nor2_1 _6714_ (.A(_0680_),
    .B(_3310_),
    .Y(_3323_));
 sky130_fd_sc_hd__a211o_1 _6715_ (.A1(net204),
    .A2(_3313_),
    .B1(_3314_),
    .C1(_3323_),
    .X(_3324_));
 sky130_fd_sc_hd__o211a_1 _6716_ (.A1(\core_1.execute.pc_high_buff_out[4] ),
    .A2(_3312_),
    .B1(_3324_),
    .C1(_3257_),
    .X(_0511_));
 sky130_fd_sc_hd__nor2_1 _6717_ (.A(_0677_),
    .B(_3310_),
    .Y(_3325_));
 sky130_fd_sc_hd__a211o_1 _6718_ (.A1(net205),
    .A2(_3313_),
    .B1(_3314_),
    .C1(_3325_),
    .X(_3326_));
 sky130_fd_sc_hd__o211a_1 _6719_ (.A1(\core_1.execute.pc_high_buff_out[5] ),
    .A2(_3312_),
    .B1(_3326_),
    .C1(_3257_),
    .X(_0512_));
 sky130_fd_sc_hd__nor2_1 _6720_ (.A(_0671_),
    .B(_3310_),
    .Y(_3327_));
 sky130_fd_sc_hd__a211o_1 _6721_ (.A1(net206),
    .A2(_3313_),
    .B1(_3314_),
    .C1(_3327_),
    .X(_3328_));
 sky130_fd_sc_hd__o211a_1 _6722_ (.A1(\core_1.execute.pc_high_buff_out[6] ),
    .A2(_3312_),
    .B1(_3328_),
    .C1(_3257_),
    .X(_0513_));
 sky130_fd_sc_hd__nand2_1 _6723_ (.A(_0611_),
    .B(_3310_),
    .Y(_3329_));
 sky130_fd_sc_hd__o211a_1 _6724_ (.A1(net115),
    .A2(_3313_),
    .B1(_3312_),
    .C1(_3329_),
    .X(_3330_));
 sky130_fd_sc_hd__a211o_1 _6725_ (.A1(\core_1.execute.pc_high_buff_out[7] ),
    .A2(_3314_),
    .B1(_3330_),
    .C1(_1165_),
    .X(_0514_));
 sky130_fd_sc_hd__dfxtp_4 _6726_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0015_),
    .Q(\core_1.decode.o_submit ));
 sky130_fd_sc_hd__dfxtp_2 _6727_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0016_),
    .Q(net178));
 sky130_fd_sc_hd__dfxtp_4 _6728_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0017_),
    .Q(net185));
 sky130_fd_sc_hd__dfxtp_4 _6729_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0018_),
    .Q(net186));
 sky130_fd_sc_hd__dfxtp_4 _6730_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0019_),
    .Q(net187));
 sky130_fd_sc_hd__dfxtp_4 _6731_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0020_),
    .Q(net188));
 sky130_fd_sc_hd__dfxtp_4 _6732_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0021_),
    .Q(net189));
 sky130_fd_sc_hd__dfxtp_4 _6733_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0022_),
    .Q(net190));
 sky130_fd_sc_hd__dfxtp_4 _6734_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0023_),
    .Q(net191));
 sky130_fd_sc_hd__dfxtp_4 _6735_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0024_),
    .Q(net192));
 sky130_fd_sc_hd__dfxtp_4 _6736_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0025_),
    .Q(net193));
 sky130_fd_sc_hd__dfxtp_4 _6737_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0026_),
    .Q(net179));
 sky130_fd_sc_hd__dfxtp_4 _6738_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0027_),
    .Q(net180));
 sky130_fd_sc_hd__dfxtp_4 _6739_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0028_),
    .Q(net181));
 sky130_fd_sc_hd__dfxtp_4 _6740_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0029_),
    .Q(net182));
 sky130_fd_sc_hd__dfxtp_4 _6741_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0030_),
    .Q(net183));
 sky130_fd_sc_hd__dfxtp_4 _6742_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0031_),
    .Q(net184));
 sky130_fd_sc_hd__dfxtp_1 _6743_ (.CLK(clknet_leaf_34_i_clk),
    .D(_0032_),
    .Q(\core_1.dec_pc_inc ));
 sky130_fd_sc_hd__dfxtp_2 _6744_ (.CLK(clknet_leaf_1_i_clk),
    .D(_0033_),
    .Q(\core_1.dec_r_bus_imm ));
 sky130_fd_sc_hd__dfxtp_1 _6745_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0034_),
    .Q(\core_1.dec_alu_flags_ie ));
 sky130_fd_sc_hd__dfxtp_1 _6746_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0035_),
    .Q(\core_1.dec_alu_carry_en ));
 sky130_fd_sc_hd__dfxtp_4 _6747_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0036_),
    .Q(\core_1.dec_l_reg_sel[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6748_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0037_),
    .Q(\core_1.dec_l_reg_sel[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6749_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0038_),
    .Q(\core_1.dec_l_reg_sel[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6750_ (.CLK(clknet_leaf_1_i_clk),
    .D(_0039_),
    .Q(\core_1.dec_rf_ie[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6751_ (.CLK(clknet_leaf_1_i_clk),
    .D(_0040_),
    .Q(\core_1.dec_rf_ie[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6752_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0041_),
    .Q(\core_1.dec_rf_ie[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6753_ (.CLK(clknet_leaf_1_i_clk),
    .D(_0042_),
    .Q(\core_1.dec_rf_ie[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6754_ (.CLK(clknet_leaf_1_i_clk),
    .D(_0043_),
    .Q(\core_1.dec_rf_ie[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6755_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0044_),
    .Q(\core_1.dec_rf_ie[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6756_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0045_),
    .Q(\core_1.dec_rf_ie[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6757_ (.CLK(clknet_leaf_1_i_clk),
    .D(_0046_),
    .Q(\core_1.dec_rf_ie[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6758_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0047_),
    .Q(\core_1.dec_r_reg_sel[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6759_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0048_),
    .Q(\core_1.dec_r_reg_sel[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6760_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0049_),
    .Q(\core_1.dec_r_reg_sel[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6761_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0050_),
    .Q(\core_1.dec_jump_cond_code[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6762_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0051_),
    .Q(\core_1.dec_jump_cond_code[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6763_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0052_),
    .Q(\core_1.dec_jump_cond_code[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6764_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0053_),
    .Q(\core_1.dec_jump_cond_code[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6765_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0054_),
    .Q(\core_1.dec_jump_cond_code[4] ));
 sky130_fd_sc_hd__dfxtp_2 _6766_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0055_),
    .Q(\core_1.de_jmp_pred ));
 sky130_fd_sc_hd__dfxtp_2 _6767_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0056_),
    .Q(\core_1.dec_mem_access ));
 sky130_fd_sc_hd__dfxtp_2 _6768_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0057_),
    .Q(\core_1.dec_mem_we ));
 sky130_fd_sc_hd__dfxtp_1 _6769_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0058_),
    .Q(\core_1.dec_used_operands[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6770_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0059_),
    .Q(\core_1.dec_used_operands[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6771_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0060_),
    .Q(\core_1.dec_sreg_load ));
 sky130_fd_sc_hd__dfxtp_4 _6772_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0061_),
    .Q(\core_1.dec_sreg_store ));
 sky130_fd_sc_hd__dfxtp_4 _6773_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0062_),
    .Q(\core_1.dec_sreg_jal_over ));
 sky130_fd_sc_hd__dfxtp_1 _6774_ (.CLK(clknet_leaf_34_i_clk),
    .D(_0063_),
    .Q(\core_1.dec_sreg_irt ));
 sky130_fd_sc_hd__dfxtp_1 _6775_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0064_),
    .Q(\core_1.dec_sys ));
 sky130_fd_sc_hd__dfxtp_1 _6776_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0065_),
    .Q(\core_1.dec_mem_width ));
 sky130_fd_sc_hd__dfxtp_1 _6777_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0066_),
    .Q(\core_1.decode.input_valid ));
 sky130_fd_sc_hd__dfxtp_2 _6778_ (.CLK(clknet_leaf_34_i_clk),
    .D(_0067_),
    .Q(\core_1.execute.sreg_priv_control.o_d[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6779_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0068_),
    .Q(\core_1.execute.sreg_data_page ));
 sky130_fd_sc_hd__dfxtp_1 _6780_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0069_),
    .Q(\core_1.execute.sreg_long_ptr_en ));
 sky130_fd_sc_hd__dfxtp_1 _6781_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0070_),
    .Q(\core_1.execute.sreg_priv_control.o_d[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6782_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0071_),
    .Q(\core_1.execute.sreg_priv_control.o_d[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6783_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0072_),
    .Q(\core_1.execute.sreg_priv_control.o_d[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6784_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0073_),
    .Q(\core_1.execute.sreg_priv_control.o_d[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6785_ (.CLK(clknet_leaf_34_i_clk),
    .D(_0074_),
    .Q(\core_1.execute.sreg_priv_control.o_d[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6786_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0075_),
    .Q(\core_1.execute.sreg_priv_control.o_d[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6787_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0076_),
    .Q(\core_1.execute.sreg_priv_control.o_d[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6788_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0077_),
    .Q(\core_1.execute.sreg_priv_control.o_d[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6789_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0078_),
    .Q(\core_1.execute.sreg_priv_control.o_d[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6790_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0079_),
    .Q(\core_1.execute.sreg_priv_control.o_d[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6791_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0080_),
    .Q(\core_1.execute.sreg_priv_control.o_d[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6792_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0081_),
    .Q(\core_1.execute.sreg_priv_control.o_d[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6793_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0082_),
    .Q(\core_1.execute.alu_mul_div.comp ));
 sky130_fd_sc_hd__dfxtp_1 _6794_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0083_),
    .Q(\core_1.fetch.out_buffer_data_instr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6795_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0084_),
    .Q(\core_1.fetch.out_buffer_data_instr[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6796_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0085_),
    .Q(\core_1.fetch.out_buffer_data_instr[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6797_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0086_),
    .Q(\core_1.fetch.out_buffer_data_instr[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6798_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0087_),
    .Q(\core_1.fetch.out_buffer_data_instr[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6799_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0088_),
    .Q(\core_1.fetch.out_buffer_data_instr[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6800_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0089_),
    .Q(\core_1.fetch.out_buffer_data_instr[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6801_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0090_),
    .Q(\core_1.fetch.out_buffer_data_instr[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6802_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0091_),
    .Q(\core_1.fetch.out_buffer_data_instr[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6803_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0092_),
    .Q(\core_1.fetch.out_buffer_data_instr[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6804_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0093_),
    .Q(\core_1.fetch.out_buffer_data_instr[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6805_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0094_),
    .Q(\core_1.fetch.out_buffer_data_instr[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6806_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0095_),
    .Q(\core_1.fetch.out_buffer_data_instr[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6807_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0096_),
    .Q(\core_1.fetch.out_buffer_data_instr[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6808_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0097_),
    .Q(\core_1.fetch.out_buffer_data_instr[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6809_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0098_),
    .Q(\core_1.fetch.out_buffer_data_instr[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6810_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0099_),
    .Q(\core_1.fetch.out_buffer_data_instr[16] ));
 sky130_fd_sc_hd__dfxtp_1 _6811_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0100_),
    .Q(\core_1.fetch.out_buffer_data_instr[17] ));
 sky130_fd_sc_hd__dfxtp_1 _6812_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0101_),
    .Q(\core_1.fetch.out_buffer_data_instr[18] ));
 sky130_fd_sc_hd__dfxtp_1 _6813_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0102_),
    .Q(\core_1.fetch.out_buffer_data_instr[19] ));
 sky130_fd_sc_hd__dfxtp_1 _6814_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0103_),
    .Q(\core_1.fetch.out_buffer_data_instr[20] ));
 sky130_fd_sc_hd__dfxtp_1 _6815_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0104_),
    .Q(\core_1.fetch.out_buffer_data_instr[21] ));
 sky130_fd_sc_hd__dfxtp_1 _6816_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0105_),
    .Q(\core_1.fetch.out_buffer_data_instr[22] ));
 sky130_fd_sc_hd__dfxtp_1 _6817_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0106_),
    .Q(\core_1.fetch.out_buffer_data_instr[23] ));
 sky130_fd_sc_hd__dfxtp_1 _6818_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0107_),
    .Q(\core_1.fetch.out_buffer_data_instr[24] ));
 sky130_fd_sc_hd__dfxtp_1 _6819_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0108_),
    .Q(\core_1.fetch.out_buffer_data_instr[25] ));
 sky130_fd_sc_hd__dfxtp_1 _6820_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0109_),
    .Q(\core_1.fetch.out_buffer_data_instr[26] ));
 sky130_fd_sc_hd__dfxtp_1 _6821_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0110_),
    .Q(\core_1.fetch.out_buffer_data_instr[27] ));
 sky130_fd_sc_hd__dfxtp_1 _6822_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0111_),
    .Q(\core_1.fetch.out_buffer_data_instr[28] ));
 sky130_fd_sc_hd__dfxtp_1 _6823_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0112_),
    .Q(\core_1.fetch.out_buffer_data_instr[29] ));
 sky130_fd_sc_hd__dfxtp_1 _6824_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0113_),
    .Q(\core_1.fetch.out_buffer_data_instr[30] ));
 sky130_fd_sc_hd__dfxtp_1 _6825_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0114_),
    .Q(\core_1.fetch.out_buffer_data_instr[31] ));
 sky130_fd_sc_hd__dfxtp_2 _6826_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0115_),
    .Q(\core_1.fetch.out_buffer_valid ));
 sky130_fd_sc_hd__dfxtp_1 _6827_ (.CLK(clknet_leaf_18_i_clk),
    .D(\core_1.fetch.current_req_branch_pred ),
    .Q(\core_1.fetch.prev_req_branch_pred ));
 sky130_fd_sc_hd__dfxtp_1 _6828_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0116_),
    .Q(\core_1.fetch.out_buffer_data_pred ));
 sky130_fd_sc_hd__dfxtp_1 _6829_ (.CLK(clknet_leaf_21_i_clk),
    .D(\core_1.fetch.submitable ),
    .Q(\core_1.decode.i_submit ));
 sky130_fd_sc_hd__dfxtp_2 _6830_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0117_),
    .Q(\core_1.fetch.prev_request_pc[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6831_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0118_),
    .Q(\core_1.fetch.prev_request_pc[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6832_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0119_),
    .Q(\core_1.fetch.prev_request_pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6833_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0120_),
    .Q(\core_1.fetch.prev_request_pc[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6834_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0121_),
    .Q(\core_1.fetch.prev_request_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6835_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0122_),
    .Q(\core_1.fetch.prev_request_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6836_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0123_),
    .Q(\core_1.fetch.prev_request_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6837_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0124_),
    .Q(\core_1.fetch.prev_request_pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6838_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0125_),
    .Q(\core_1.fetch.prev_request_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6839_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0126_),
    .Q(\core_1.fetch.prev_request_pc[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6840_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0127_),
    .Q(\core_1.fetch.prev_request_pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6841_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0128_),
    .Q(\core_1.fetch.prev_request_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6842_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0129_),
    .Q(\core_1.fetch.prev_request_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6843_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0130_),
    .Q(\core_1.fetch.prev_request_pc[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6844_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0131_),
    .Q(\core_1.fetch.prev_request_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6845_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0132_),
    .Q(\core_1.fetch.prev_request_pc[15] ));
 sky130_fd_sc_hd__dfxtp_4 _6846_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0133_),
    .Q(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6847_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0134_),
    .Q(\core_1.decode.i_instr_l[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6848_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0135_),
    .Q(\core_1.decode.i_instr_l[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6849_ (.CLK(clknet_leaf_1_i_clk),
    .D(_0136_),
    .Q(\core_1.decode.i_instr_l[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6850_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0137_),
    .Q(\core_1.decode.i_instr_l[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6851_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0138_),
    .Q(\core_1.decode.i_instr_l[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6852_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0139_),
    .Q(\core_1.decode.i_instr_l[6] ));
 sky130_fd_sc_hd__dfxtp_2 _6853_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0140_),
    .Q(\core_1.decode.i_instr_l[7] ));
 sky130_fd_sc_hd__dfxtp_2 _6854_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0141_),
    .Q(\core_1.decode.i_instr_l[8] ));
 sky130_fd_sc_hd__dfxtp_2 _6855_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0142_),
    .Q(\core_1.decode.i_instr_l[9] ));
 sky130_fd_sc_hd__dfxtp_2 _6856_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0143_),
    .Q(\core_1.decode.i_instr_l[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6857_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0144_),
    .Q(\core_1.decode.i_instr_l[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6858_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0145_),
    .Q(\core_1.decode.i_instr_l[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6859_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0146_),
    .Q(\core_1.decode.i_instr_l[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6860_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0147_),
    .Q(\core_1.decode.i_instr_l[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6861_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0148_),
    .Q(\core_1.decode.i_instr_l[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6862_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0149_),
    .Q(\core_1.decode.i_imm_pass[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6863_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0150_),
    .Q(\core_1.decode.i_imm_pass[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6864_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0151_),
    .Q(\core_1.decode.i_imm_pass[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6865_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0152_),
    .Q(\core_1.decode.i_imm_pass[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6866_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0153_),
    .Q(\core_1.decode.i_imm_pass[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6867_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0154_),
    .Q(\core_1.decode.i_imm_pass[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6868_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0155_),
    .Q(\core_1.decode.i_imm_pass[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6869_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0156_),
    .Q(\core_1.decode.i_imm_pass[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6870_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0157_),
    .Q(\core_1.decode.i_imm_pass[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6871_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0158_),
    .Q(\core_1.decode.i_imm_pass[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6872_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0159_),
    .Q(\core_1.decode.i_imm_pass[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6873_ (.CLK(clknet_leaf_15_i_clk),
    .D(_0160_),
    .Q(\core_1.decode.i_imm_pass[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6874_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0161_),
    .Q(\core_1.decode.i_imm_pass[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6875_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0162_),
    .Q(\core_1.decode.i_imm_pass[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6876_ (.CLK(clknet_leaf_14_i_clk),
    .D(_0163_),
    .Q(\core_1.decode.i_imm_pass[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6877_ (.CLK(clknet_leaf_16_i_clk),
    .D(_0164_),
    .Q(\core_1.decode.i_imm_pass[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6878_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0165_),
    .Q(\core_1.fetch.dbg_out ));
 sky130_fd_sc_hd__dfxtp_1 _6879_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0166_),
    .Q(\core_1.fetch.flush_event_invalidate ));
 sky130_fd_sc_hd__dfxtp_1 _6880_ (.CLK(clknet_leaf_18_i_clk),
    .D(_0167_),
    .Q(\core_1.fetch.pc_flush_override ));
 sky130_fd_sc_hd__dfxtp_1 _6881_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0168_),
    .Q(\core_1.fetch.pc_reset_override ));
 sky130_fd_sc_hd__dfxtp_4 _6882_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0169_),
    .Q(net156));
 sky130_fd_sc_hd__dfxtp_1 _6883_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0170_),
    .Q(\core_1.decode.i_jmp_pred_pass ));
 sky130_fd_sc_hd__dfxtp_4 _6884_ (.CLK(clknet_leaf_34_i_clk),
    .D(_0171_),
    .Q(net79));
 sky130_fd_sc_hd__dfxtp_1 _6885_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0004_),
    .Q(\core_1.decode.oc_alu_mode[1] ));
 sky130_fd_sc_hd__dfxtp_4 _6886_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0005_),
    .Q(\core_1.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6887_ (.CLK(clknet_leaf_1_i_clk),
    .D(_0006_),
    .Q(\core_1.decode.oc_alu_mode[3] ));
 sky130_fd_sc_hd__dfxtp_4 _6888_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0007_),
    .Q(\core_1.decode.oc_alu_mode[4] ));
 sky130_fd_sc_hd__dfxtp_4 _6889_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0008_),
    .Q(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__dfxtp_4 _6890_ (.CLK(clknet_leaf_1_i_clk),
    .D(_0009_),
    .Q(\core_1.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__dfxtp_4 _6891_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0010_),
    .Q(\core_1.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__dfxtp_2 _6892_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0011_),
    .Q(\core_1.execute.alu_mul_div.i_mul ));
 sky130_fd_sc_hd__dfxtp_4 _6893_ (.CLK(clknet_leaf_1_i_clk),
    .D(_0012_),
    .Q(\core_1.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__dfxtp_4 _6894_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0000_),
    .Q(\core_1.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__dfxtp_1 _6895_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0001_),
    .Q(\core_1.decode.oc_alu_mode[11] ));
 sky130_fd_sc_hd__dfxtp_4 _6896_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0002_),
    .Q(\core_1.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__dfxtp_2 _6897_ (.CLK(clknet_leaf_36_i_clk),
    .D(_0003_),
    .Q(\core_1.decode.oc_alu_mode[13] ));
 sky130_fd_sc_hd__dfxtp_2 _6898_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0172_),
    .Q(\core_1.execute.alu_mul_div.div_cur[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6899_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0173_),
    .Q(\core_1.execute.alu_mul_div.div_cur[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6900_ (.CLK(clknet_leaf_38_i_clk),
    .D(_0174_),
    .Q(\core_1.execute.alu_mul_div.div_cur[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6901_ (.CLK(clknet_leaf_38_i_clk),
    .D(_0175_),
    .Q(\core_1.execute.alu_mul_div.div_cur[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6902_ (.CLK(clknet_leaf_37_i_clk),
    .D(_0176_),
    .Q(\core_1.execute.alu_mul_div.div_cur[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6903_ (.CLK(clknet_leaf_38_i_clk),
    .D(_0177_),
    .Q(\core_1.execute.alu_mul_div.div_cur[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6904_ (.CLK(clknet_leaf_38_i_clk),
    .D(_0178_),
    .Q(\core_1.execute.alu_mul_div.div_cur[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6905_ (.CLK(clknet_leaf_38_i_clk),
    .D(_0179_),
    .Q(\core_1.execute.alu_mul_div.div_cur[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6906_ (.CLK(clknet_leaf_38_i_clk),
    .D(_0180_),
    .Q(\core_1.execute.alu_mul_div.div_cur[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6907_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0181_),
    .Q(\core_1.execute.alu_mul_div.div_cur[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6908_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0182_),
    .Q(\core_1.execute.alu_mul_div.div_cur[11] ));
 sky130_fd_sc_hd__dfxtp_2 _6909_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0183_),
    .Q(\core_1.execute.alu_mul_div.div_cur[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6910_ (.CLK(clknet_leaf_38_i_clk),
    .D(_0184_),
    .Q(\core_1.execute.alu_mul_div.div_cur[13] ));
 sky130_fd_sc_hd__dfxtp_2 _6911_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0185_),
    .Q(\core_1.execute.alu_mul_div.div_cur[14] ));
 sky130_fd_sc_hd__dfxtp_2 _6912_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0186_),
    .Q(\core_1.execute.alu_mul_div.div_cur[15] ));
 sky130_fd_sc_hd__dfxtp_2 _6913_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0187_),
    .Q(\core_1.execute.alu_mul_div.div_cur[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6914_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0188_),
    .Q(\core_1.execute.alu_mul_div.cbit[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6915_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0189_),
    .Q(\core_1.execute.alu_mul_div.cbit[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6916_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0190_),
    .Q(\core_1.execute.alu_mul_div.cbit[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6917_ (.CLK(clknet_leaf_35_i_clk),
    .D(_0191_),
    .Q(\core_1.dec_mem_long ));
 sky130_fd_sc_hd__dfxtp_1 _6918_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0192_),
    .Q(net104));
 sky130_fd_sc_hd__dfxtp_1 _6919_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0014_),
    .Q(net107));
 sky130_fd_sc_hd__dfxtp_1 _6920_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0193_),
    .Q(\core_1.execute.mem_stage_pc[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6921_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0194_),
    .Q(\core_1.execute.mem_stage_pc[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6922_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0195_),
    .Q(\core_1.execute.mem_stage_pc[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6923_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0196_),
    .Q(\core_1.execute.mem_stage_pc[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6924_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0197_),
    .Q(\core_1.execute.mem_stage_pc[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6925_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0198_),
    .Q(\core_1.execute.mem_stage_pc[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6926_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0199_),
    .Q(\core_1.execute.mem_stage_pc[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6927_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0200_),
    .Q(\core_1.execute.mem_stage_pc[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6928_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0201_),
    .Q(\core_1.execute.mem_stage_pc[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6929_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0202_),
    .Q(\core_1.execute.mem_stage_pc[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6930_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0203_),
    .Q(\core_1.execute.mem_stage_pc[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6931_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0204_),
    .Q(\core_1.execute.mem_stage_pc[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6932_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0205_),
    .Q(\core_1.execute.mem_stage_pc[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6933_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0206_),
    .Q(\core_1.execute.mem_stage_pc[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6934_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0207_),
    .Q(\core_1.execute.mem_stage_pc[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6935_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0208_),
    .Q(\core_1.execute.mem_stage_pc[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6936_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0209_),
    .Q(\core_1.execute.prev_pc_high[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6937_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0210_),
    .Q(\core_1.execute.prev_pc_high[1] ));
 sky130_fd_sc_hd__dfxtp_1 _6938_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0211_),
    .Q(\core_1.execute.prev_pc_high[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6939_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0212_),
    .Q(\core_1.execute.prev_pc_high[3] ));
 sky130_fd_sc_hd__dfxtp_1 _6940_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0213_),
    .Q(\core_1.execute.prev_pc_high[4] ));
 sky130_fd_sc_hd__dfxtp_1 _6941_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0214_),
    .Q(\core_1.execute.prev_pc_high[5] ));
 sky130_fd_sc_hd__dfxtp_1 _6942_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0215_),
    .Q(\core_1.execute.prev_pc_high[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6943_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0216_),
    .Q(\core_1.execute.prev_pc_high[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6944_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0217_),
    .Q(\core_1.execute.sreg_irq_flags.i_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _6945_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0218_),
    .Q(\core_1.execute.prev_sys ));
 sky130_fd_sc_hd__dfxtp_1 _6946_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0219_),
    .Q(net159));
 sky130_fd_sc_hd__dfxtp_1 _6947_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0220_),
    .Q(\core_1.ew_addr_high[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6948_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0221_),
    .Q(net132));
 sky130_fd_sc_hd__dfxtp_1 _6949_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0222_),
    .Q(net133));
 sky130_fd_sc_hd__dfxtp_1 _6950_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0223_),
    .Q(net134));
 sky130_fd_sc_hd__dfxtp_2 _6951_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0224_),
    .Q(net135));
 sky130_fd_sc_hd__dfxtp_2 _6952_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0225_),
    .Q(net136));
 sky130_fd_sc_hd__dfxtp_2 _6953_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0226_),
    .Q(net137));
 sky130_fd_sc_hd__dfxtp_2 _6954_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0227_),
    .Q(net138));
 sky130_fd_sc_hd__dfxtp_1 _6955_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0228_),
    .Q(\core_1.ew_submit ));
 sky130_fd_sc_hd__dfxtp_2 _6956_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0229_),
    .Q(\core_1.ew_data[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6957_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0230_),
    .Q(\core_1.ew_data[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6958_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0231_),
    .Q(\core_1.ew_data[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6959_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0232_),
    .Q(\core_1.ew_data[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6960_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0233_),
    .Q(\core_1.ew_data[4] ));
 sky130_fd_sc_hd__dfxtp_2 _6961_ (.CLK(clknet_leaf_25_i_clk),
    .D(_0234_),
    .Q(\core_1.ew_data[5] ));
 sky130_fd_sc_hd__dfxtp_2 _6962_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0235_),
    .Q(\core_1.ew_data[6] ));
 sky130_fd_sc_hd__dfxtp_1 _6963_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0236_),
    .Q(\core_1.ew_data[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6964_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0237_),
    .Q(\core_1.ew_data[8] ));
 sky130_fd_sc_hd__dfxtp_1 _6965_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0238_),
    .Q(\core_1.ew_data[9] ));
 sky130_fd_sc_hd__dfxtp_1 _6966_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0239_),
    .Q(\core_1.ew_data[10] ));
 sky130_fd_sc_hd__dfxtp_1 _6967_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0240_),
    .Q(\core_1.ew_data[11] ));
 sky130_fd_sc_hd__dfxtp_1 _6968_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0241_),
    .Q(\core_1.ew_data[12] ));
 sky130_fd_sc_hd__dfxtp_1 _6969_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0242_),
    .Q(\core_1.ew_data[13] ));
 sky130_fd_sc_hd__dfxtp_1 _6970_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0243_),
    .Q(\core_1.ew_data[14] ));
 sky130_fd_sc_hd__dfxtp_1 _6971_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0244_),
    .Q(\core_1.ew_data[15] ));
 sky130_fd_sc_hd__dfxtp_1 _6972_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0245_),
    .Q(\core_1.ew_addr[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6973_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0246_),
    .Q(net116));
 sky130_fd_sc_hd__dfxtp_1 _6974_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0247_),
    .Q(net123));
 sky130_fd_sc_hd__dfxtp_1 _6975_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0248_),
    .Q(net124));
 sky130_fd_sc_hd__dfxtp_1 _6976_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0249_),
    .Q(net125));
 sky130_fd_sc_hd__dfxtp_1 _6977_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0250_),
    .Q(net126));
 sky130_fd_sc_hd__dfxtp_1 _6978_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0251_),
    .Q(net127));
 sky130_fd_sc_hd__dfxtp_1 _6979_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0252_),
    .Q(net128));
 sky130_fd_sc_hd__dfxtp_1 _6980_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0253_),
    .Q(net129));
 sky130_fd_sc_hd__dfxtp_1 _6981_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0254_),
    .Q(net130));
 sky130_fd_sc_hd__dfxtp_1 _6982_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0255_),
    .Q(net131));
 sky130_fd_sc_hd__dfxtp_1 _6983_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0256_),
    .Q(net117));
 sky130_fd_sc_hd__dfxtp_1 _6984_ (.CLK(clknet_leaf_17_i_clk),
    .D(_0257_),
    .Q(net118));
 sky130_fd_sc_hd__dfxtp_1 _6985_ (.CLK(clknet_leaf_19_i_clk),
    .D(_0258_),
    .Q(net119));
 sky130_fd_sc_hd__dfxtp_1 _6986_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0259_),
    .Q(net120));
 sky130_fd_sc_hd__dfxtp_1 _6987_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0260_),
    .Q(net121));
 sky130_fd_sc_hd__dfxtp_2 _6988_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0261_),
    .Q(\core_1.ew_reg_ie[0] ));
 sky130_fd_sc_hd__dfxtp_1 _6989_ (.CLK(clknet_leaf_1_i_clk),
    .D(_0262_),
    .Q(\core_1.ew_reg_ie[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6990_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0263_),
    .Q(\core_1.ew_reg_ie[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6991_ (.CLK(clknet_leaf_1_i_clk),
    .D(_0264_),
    .Q(\core_1.ew_reg_ie[3] ));
 sky130_fd_sc_hd__dfxtp_4 _6992_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0265_),
    .Q(\core_1.ew_reg_ie[4] ));
 sky130_fd_sc_hd__dfxtp_2 _6993_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0266_),
    .Q(\core_1.ew_reg_ie[5] ));
 sky130_fd_sc_hd__dfxtp_2 _6994_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0267_),
    .Q(\core_1.ew_reg_ie[6] ));
 sky130_fd_sc_hd__dfxtp_2 _6995_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0268_),
    .Q(\core_1.ew_reg_ie[7] ));
 sky130_fd_sc_hd__dfxtp_1 _6996_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0269_),
    .Q(\core_1.ew_mem_access ));
 sky130_fd_sc_hd__dfxtp_2 _6997_ (.CLK(clknet_leaf_9_i_clk),
    .D(_0270_),
    .Q(\core_1.ew_mem_width ));
 sky130_fd_sc_hd__dfxtp_4 _6998_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0013_),
    .Q(\core_1.decode.i_flush ));
 sky130_fd_sc_hd__dfxtp_4 _6999_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0271_),
    .Q(net155));
 sky130_fd_sc_hd__dfxtp_1 _7000_ (.CLK(clknet_leaf_34_i_clk),
    .D(_0272_),
    .Q(\core_1.execute.hold_valid ));
 sky130_fd_sc_hd__dfxtp_1 _7001_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0273_),
    .Q(\core_1.execute.rf.reg_outputs[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7002_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0274_),
    .Q(\core_1.execute.rf.reg_outputs[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7003_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0275_),
    .Q(\core_1.execute.rf.reg_outputs[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7004_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0276_),
    .Q(\core_1.execute.rf.reg_outputs[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7005_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0277_),
    .Q(\core_1.execute.rf.reg_outputs[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7006_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0278_),
    .Q(\core_1.execute.rf.reg_outputs[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7007_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0279_),
    .Q(\core_1.execute.rf.reg_outputs[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7008_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0280_),
    .Q(\core_1.execute.rf.reg_outputs[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7009_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0281_),
    .Q(\core_1.execute.rf.reg_outputs[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7010_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0282_),
    .Q(\core_1.execute.rf.reg_outputs[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7011_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0283_),
    .Q(\core_1.execute.rf.reg_outputs[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7012_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0284_),
    .Q(\core_1.execute.rf.reg_outputs[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7013_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0285_),
    .Q(\core_1.execute.rf.reg_outputs[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7014_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0286_),
    .Q(\core_1.execute.rf.reg_outputs[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7015_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0287_),
    .Q(\core_1.execute.rf.reg_outputs[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7016_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0288_),
    .Q(\core_1.execute.rf.reg_outputs[7][15] ));
 sky130_fd_sc_hd__dfxtp_2 _7017_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0289_),
    .Q(\core_1.execute.rf.reg_outputs[6][0] ));
 sky130_fd_sc_hd__dfxtp_2 _7018_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0290_),
    .Q(\core_1.execute.rf.reg_outputs[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7019_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0291_),
    .Q(\core_1.execute.rf.reg_outputs[6][2] ));
 sky130_fd_sc_hd__dfxtp_2 _7020_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0292_),
    .Q(\core_1.execute.rf.reg_outputs[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7021_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0293_),
    .Q(\core_1.execute.rf.reg_outputs[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7022_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0294_),
    .Q(\core_1.execute.rf.reg_outputs[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7023_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0295_),
    .Q(\core_1.execute.rf.reg_outputs[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7024_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0296_),
    .Q(\core_1.execute.rf.reg_outputs[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7025_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0297_),
    .Q(\core_1.execute.rf.reg_outputs[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7026_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0298_),
    .Q(\core_1.execute.rf.reg_outputs[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7027_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0299_),
    .Q(\core_1.execute.rf.reg_outputs[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7028_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0300_),
    .Q(\core_1.execute.rf.reg_outputs[6][11] ));
 sky130_fd_sc_hd__dfxtp_2 _7029_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0301_),
    .Q(\core_1.execute.rf.reg_outputs[6][12] ));
 sky130_fd_sc_hd__dfxtp_2 _7030_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0302_),
    .Q(\core_1.execute.rf.reg_outputs[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7031_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0303_),
    .Q(\core_1.execute.rf.reg_outputs[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7032_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0304_),
    .Q(\core_1.execute.rf.reg_outputs[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7033_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0305_),
    .Q(\core_1.execute.rf.reg_outputs[5][0] ));
 sky130_fd_sc_hd__dfxtp_2 _7034_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0306_),
    .Q(\core_1.execute.rf.reg_outputs[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7035_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0307_),
    .Q(\core_1.execute.rf.reg_outputs[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7036_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0308_),
    .Q(\core_1.execute.rf.reg_outputs[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7037_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0309_),
    .Q(\core_1.execute.rf.reg_outputs[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7038_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0310_),
    .Q(\core_1.execute.rf.reg_outputs[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7039_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0311_),
    .Q(\core_1.execute.rf.reg_outputs[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7040_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0312_),
    .Q(\core_1.execute.rf.reg_outputs[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7041_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0313_),
    .Q(\core_1.execute.rf.reg_outputs[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7042_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0314_),
    .Q(\core_1.execute.rf.reg_outputs[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7043_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0315_),
    .Q(\core_1.execute.rf.reg_outputs[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7044_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0316_),
    .Q(\core_1.execute.rf.reg_outputs[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7045_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0317_),
    .Q(\core_1.execute.rf.reg_outputs[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7046_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0318_),
    .Q(\core_1.execute.rf.reg_outputs[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7047_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0319_),
    .Q(\core_1.execute.rf.reg_outputs[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7048_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0320_),
    .Q(\core_1.execute.rf.reg_outputs[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7049_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0321_),
    .Q(\core_1.execute.rf.reg_outputs[4][0] ));
 sky130_fd_sc_hd__dfxtp_2 _7050_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0322_),
    .Q(\core_1.execute.rf.reg_outputs[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7051_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0323_),
    .Q(\core_1.execute.rf.reg_outputs[4][2] ));
 sky130_fd_sc_hd__dfxtp_2 _7052_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0324_),
    .Q(\core_1.execute.rf.reg_outputs[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7053_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0325_),
    .Q(\core_1.execute.rf.reg_outputs[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7054_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0326_),
    .Q(\core_1.execute.rf.reg_outputs[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7055_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0327_),
    .Q(\core_1.execute.rf.reg_outputs[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7056_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0328_),
    .Q(\core_1.execute.rf.reg_outputs[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7057_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0329_),
    .Q(\core_1.execute.rf.reg_outputs[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7058_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0330_),
    .Q(\core_1.execute.rf.reg_outputs[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7059_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0331_),
    .Q(\core_1.execute.rf.reg_outputs[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7060_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0332_),
    .Q(\core_1.execute.rf.reg_outputs[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7061_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0333_),
    .Q(\core_1.execute.rf.reg_outputs[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7062_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0334_),
    .Q(\core_1.execute.rf.reg_outputs[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7063_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0335_),
    .Q(\core_1.execute.rf.reg_outputs[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7064_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0336_),
    .Q(\core_1.execute.rf.reg_outputs[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7065_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0337_),
    .Q(\core_1.execute.rf.reg_outputs[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7066_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0338_),
    .Q(\core_1.execute.rf.reg_outputs[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7067_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0339_),
    .Q(\core_1.execute.rf.reg_outputs[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7068_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0340_),
    .Q(\core_1.execute.rf.reg_outputs[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7069_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0341_),
    .Q(\core_1.execute.rf.reg_outputs[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7070_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0342_),
    .Q(\core_1.execute.rf.reg_outputs[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7071_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0343_),
    .Q(\core_1.execute.rf.reg_outputs[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7072_ (.CLK(clknet_leaf_3_i_clk),
    .D(_0344_),
    .Q(\core_1.execute.rf.reg_outputs[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7073_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0345_),
    .Q(\core_1.execute.rf.reg_outputs[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7074_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0346_),
    .Q(\core_1.execute.rf.reg_outputs[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7075_ (.CLK(clknet_leaf_12_i_clk),
    .D(_0347_),
    .Q(\core_1.execute.rf.reg_outputs[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7076_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0348_),
    .Q(\core_1.execute.rf.reg_outputs[3][11] ));
 sky130_fd_sc_hd__dfxtp_2 _7077_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0349_),
    .Q(\core_1.execute.rf.reg_outputs[3][12] ));
 sky130_fd_sc_hd__dfxtp_2 _7078_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0350_),
    .Q(\core_1.execute.rf.reg_outputs[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7079_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0351_),
    .Q(\core_1.execute.rf.reg_outputs[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7080_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0352_),
    .Q(\core_1.execute.rf.reg_outputs[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7081_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0353_),
    .Q(\core_1.execute.rf.reg_outputs[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7082_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0354_),
    .Q(\core_1.execute.rf.reg_outputs[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7083_ (.CLK(clknet_leaf_5_i_clk),
    .D(_0355_),
    .Q(\core_1.execute.rf.reg_outputs[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _7084_ (.CLK(clknet_leaf_7_i_clk),
    .D(_0356_),
    .Q(\core_1.execute.rf.reg_outputs[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7085_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0357_),
    .Q(\core_1.execute.rf.reg_outputs[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7086_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0358_),
    .Q(\core_1.execute.rf.reg_outputs[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7087_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0359_),
    .Q(\core_1.execute.rf.reg_outputs[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7088_ (.CLK(clknet_leaf_4_i_clk),
    .D(_0360_),
    .Q(\core_1.execute.rf.reg_outputs[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7089_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0361_),
    .Q(\core_1.execute.rf.reg_outputs[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7090_ (.CLK(clknet_leaf_7_i_clk),
    .D(_0362_),
    .Q(\core_1.execute.rf.reg_outputs[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7091_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0363_),
    .Q(\core_1.execute.rf.reg_outputs[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7092_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0364_),
    .Q(\core_1.execute.rf.reg_outputs[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7093_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0365_),
    .Q(\core_1.execute.rf.reg_outputs[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7094_ (.CLK(clknet_leaf_7_i_clk),
    .D(_0366_),
    .Q(\core_1.execute.rf.reg_outputs[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7095_ (.CLK(clknet_leaf_6_i_clk),
    .D(_0367_),
    .Q(\core_1.execute.rf.reg_outputs[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7096_ (.CLK(clknet_leaf_7_i_clk),
    .D(_0368_),
    .Q(\core_1.execute.rf.reg_outputs[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _7097_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0369_),
    .Q(\core_1.execute.rf.reg_outputs[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _7098_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0370_),
    .Q(\core_1.execute.rf.reg_outputs[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _7099_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0371_),
    .Q(\core_1.execute.rf.reg_outputs[1][2] ));
 sky130_fd_sc_hd__dfxtp_2 _7100_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0372_),
    .Q(\core_1.execute.rf.reg_outputs[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _7101_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0373_),
    .Q(\core_1.execute.rf.reg_outputs[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _7102_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0374_),
    .Q(\core_1.execute.rf.reg_outputs[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _7103_ (.CLK(clknet_leaf_2_i_clk),
    .D(_0375_),
    .Q(\core_1.execute.rf.reg_outputs[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _7104_ (.CLK(clknet_leaf_8_i_clk),
    .D(_0376_),
    .Q(\core_1.execute.rf.reg_outputs[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _7105_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0377_),
    .Q(\core_1.execute.rf.reg_outputs[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _7106_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0378_),
    .Q(\core_1.execute.rf.reg_outputs[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _7107_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0379_),
    .Q(\core_1.execute.rf.reg_outputs[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _7108_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0380_),
    .Q(\core_1.execute.rf.reg_outputs[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _7109_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0381_),
    .Q(\core_1.execute.rf.reg_outputs[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _7110_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0382_),
    .Q(\core_1.execute.rf.reg_outputs[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _7111_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0383_),
    .Q(\core_1.execute.rf.reg_outputs[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _7112_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0384_),
    .Q(\core_1.execute.rf.reg_outputs[1][15] ));
 sky130_fd_sc_hd__dfxtp_4 _7113_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0385_),
    .Q(net88));
 sky130_fd_sc_hd__dfxtp_4 _7114_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0386_),
    .Q(net95));
 sky130_fd_sc_hd__dfxtp_4 _7115_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0387_),
    .Q(net96));
 sky130_fd_sc_hd__dfxtp_4 _7116_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0388_),
    .Q(net97));
 sky130_fd_sc_hd__dfxtp_4 _7117_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0389_),
    .Q(net98));
 sky130_fd_sc_hd__dfxtp_4 _7118_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0390_),
    .Q(net99));
 sky130_fd_sc_hd__dfxtp_4 _7119_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0391_),
    .Q(net100));
 sky130_fd_sc_hd__dfxtp_4 _7120_ (.CLK(clknet_leaf_10_i_clk),
    .D(_0392_),
    .Q(net101));
 sky130_fd_sc_hd__dfxtp_4 _7121_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0393_),
    .Q(net102));
 sky130_fd_sc_hd__dfxtp_4 _7122_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0394_),
    .Q(net103));
 sky130_fd_sc_hd__dfxtp_4 _7123_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0395_),
    .Q(net89));
 sky130_fd_sc_hd__dfxtp_4 _7124_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0396_),
    .Q(net90));
 sky130_fd_sc_hd__dfxtp_2 _7125_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0397_),
    .Q(net91));
 sky130_fd_sc_hd__dfxtp_2 _7126_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0398_),
    .Q(net92));
 sky130_fd_sc_hd__dfxtp_4 _7127_ (.CLK(clknet_leaf_13_i_clk),
    .D(_0399_),
    .Q(net93));
 sky130_fd_sc_hd__dfxtp_4 _7128_ (.CLK(clknet_leaf_11_i_clk),
    .D(_0400_),
    .Q(net94));
 sky130_fd_sc_hd__dfxtp_2 _7129_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0401_),
    .Q(\core_1.execute.irq_en ));
 sky130_fd_sc_hd__dfxtp_2 _7130_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0402_),
    .Q(\core_1.execute.alu_mul_div.cbit[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7131_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0403_),
    .Q(\core_1.execute.alu_mul_div.mul_res[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7132_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0404_),
    .Q(\core_1.execute.alu_mul_div.mul_res[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7133_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0405_),
    .Q(\core_1.execute.alu_mul_div.mul_res[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7134_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0406_),
    .Q(\core_1.execute.alu_mul_div.mul_res[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7135_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0407_),
    .Q(\core_1.execute.alu_mul_div.mul_res[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7136_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0408_),
    .Q(\core_1.execute.alu_mul_div.mul_res[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7137_ (.CLK(clknet_leaf_0_i_clk),
    .D(_0409_),
    .Q(\core_1.execute.alu_mul_div.mul_res[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7138_ (.CLK(clknet_leaf_0_i_clk),
    .D(_0410_),
    .Q(\core_1.execute.alu_mul_div.mul_res[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7139_ (.CLK(clknet_leaf_0_i_clk),
    .D(_0411_),
    .Q(\core_1.execute.alu_mul_div.mul_res[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7140_ (.CLK(clknet_leaf_0_i_clk),
    .D(_0412_),
    .Q(\core_1.execute.alu_mul_div.mul_res[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7141_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0413_),
    .Q(\core_1.execute.alu_mul_div.mul_res[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7142_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0414_),
    .Q(\core_1.execute.alu_mul_div.mul_res[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7143_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0415_),
    .Q(\core_1.execute.alu_mul_div.mul_res[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7144_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0416_),
    .Q(\core_1.execute.alu_mul_div.mul_res[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7145_ (.CLK(clknet_leaf_43_i_clk),
    .D(_0417_),
    .Q(\core_1.execute.alu_mul_div.mul_res[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7146_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0418_),
    .Q(\core_1.execute.alu_mul_div.mul_res[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7147_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0419_),
    .Q(\core_1.execute.next_ready_delayed ));
 sky130_fd_sc_hd__dfxtp_1 _7148_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0420_),
    .Q(\core_1.execute.alu_mul_div.div_res[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7149_ (.CLK(clknet_leaf_42_i_clk),
    .D(_0421_),
    .Q(\core_1.execute.alu_mul_div.div_res[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7150_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0422_),
    .Q(\core_1.execute.alu_mul_div.div_res[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7151_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0423_),
    .Q(\core_1.execute.alu_mul_div.div_res[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7152_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0424_),
    .Q(\core_1.execute.alu_mul_div.div_res[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7153_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0425_),
    .Q(\core_1.execute.alu_mul_div.div_res[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7154_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0426_),
    .Q(\core_1.execute.alu_mul_div.div_res[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7155_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0427_),
    .Q(\core_1.execute.alu_mul_div.div_res[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7156_ (.CLK(clknet_leaf_41_i_clk),
    .D(_0428_),
    .Q(\core_1.execute.alu_mul_div.div_res[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7157_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0429_),
    .Q(\core_1.execute.alu_mul_div.div_res[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7158_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0430_),
    .Q(\core_1.execute.alu_mul_div.div_res[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7159_ (.CLK(clknet_leaf_40_i_clk),
    .D(_0431_),
    .Q(\core_1.execute.alu_mul_div.div_res[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7160_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0432_),
    .Q(\core_1.execute.alu_mul_div.div_res[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7161_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0433_),
    .Q(\core_1.execute.alu_mul_div.div_res[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7162_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0434_),
    .Q(\core_1.execute.alu_mul_div.div_res[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7163_ (.CLK(clknet_leaf_39_i_clk),
    .D(_0435_),
    .Q(\core_1.execute.alu_mul_div.div_res[15] ));
 sky130_fd_sc_hd__dfxtp_4 _7164_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0436_),
    .Q(net72));
 sky130_fd_sc_hd__dfxtp_4 _7165_ (.CLK(clknet_leaf_34_i_clk),
    .D(_0437_),
    .Q(net80));
 sky130_fd_sc_hd__dfxtp_2 _7166_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0438_),
    .Q(net81));
 sky130_fd_sc_hd__dfxtp_4 _7167_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0439_),
    .Q(net82));
 sky130_fd_sc_hd__dfxtp_4 _7168_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0440_),
    .Q(net83));
 sky130_fd_sc_hd__dfxtp_4 _7169_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0441_),
    .Q(net84));
 sky130_fd_sc_hd__dfxtp_4 _7170_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0442_),
    .Q(net85));
 sky130_fd_sc_hd__dfxtp_4 _7171_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0443_),
    .Q(net86));
 sky130_fd_sc_hd__dfxtp_4 _7172_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0444_),
    .Q(net87));
 sky130_fd_sc_hd__dfxtp_4 _7173_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0445_),
    .Q(net73));
 sky130_fd_sc_hd__dfxtp_4 _7174_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0446_),
    .Q(net74));
 sky130_fd_sc_hd__dfxtp_4 _7175_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0447_),
    .Q(net75));
 sky130_fd_sc_hd__dfxtp_4 _7176_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0448_),
    .Q(net76));
 sky130_fd_sc_hd__dfxtp_4 _7177_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0449_),
    .Q(net77));
 sky130_fd_sc_hd__dfxtp_4 _7178_ (.CLK(clknet_leaf_24_i_clk),
    .D(_0450_),
    .Q(net78));
 sky130_fd_sc_hd__dfxtp_2 _7179_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0451_),
    .Q(\core_1.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7180_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0452_),
    .Q(\core_1.execute.alu_flag_reg.o_d[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7181_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0453_),
    .Q(\core_1.execute.alu_flag_reg.o_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7182_ (.CLK(clknet_leaf_34_i_clk),
    .D(_0454_),
    .Q(\core_1.execute.alu_flag_reg.o_d[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7183_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0455_),
    .Q(\core_1.execute.alu_flag_reg.o_d[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7184_ (.CLK(clknet_leaf_34_i_clk),
    .D(_0456_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7185_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0457_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7186_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0458_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7187_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0459_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7188_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0460_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7189_ (.CLK(clknet_leaf_26_i_clk),
    .D(_0461_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7190_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0462_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7191_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0463_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7192_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0464_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7193_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0465_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7194_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0466_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7195_ (.CLK(clknet_leaf_20_i_clk),
    .D(_0467_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7196_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0468_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7197_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0469_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7198_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0470_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7199_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0471_),
    .Q(\core_1.execute.sreg_irq_pc.o_d[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7200_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0472_),
    .Q(\core_1.execute.sreg_jtr_buff.o_d[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7201_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0473_),
    .Q(\core_1.execute.sreg_jtr_buff.o_d[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7202_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0474_),
    .Q(\core_1.execute.sreg_jtr_buff.o_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7203_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0475_),
    .Q(net106));
 sky130_fd_sc_hd__dfxtp_1 _7204_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0476_),
    .Q(\core_1.execute.trap_flag ));
 sky130_fd_sc_hd__dfxtp_2 _7205_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0477_),
    .Q(net105));
 sky130_fd_sc_hd__dfxtp_1 _7206_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0478_),
    .Q(\core_1.execute.sreg_scratch.o_d[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7207_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0479_),
    .Q(\core_1.execute.sreg_scratch.o_d[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7208_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0480_),
    .Q(\core_1.execute.sreg_scratch.o_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7209_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0481_),
    .Q(\core_1.execute.sreg_scratch.o_d[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7210_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0482_),
    .Q(\core_1.execute.sreg_scratch.o_d[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7211_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0483_),
    .Q(\core_1.execute.sreg_scratch.o_d[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7212_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0484_),
    .Q(\core_1.execute.sreg_scratch.o_d[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7213_ (.CLK(clknet_leaf_33_i_clk),
    .D(_0485_),
    .Q(\core_1.execute.sreg_scratch.o_d[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7214_ (.CLK(clknet_leaf_34_i_clk),
    .D(_0486_),
    .Q(\core_1.execute.sreg_scratch.o_d[8] ));
 sky130_fd_sc_hd__dfxtp_1 _7215_ (.CLK(clknet_leaf_23_i_clk),
    .D(_0487_),
    .Q(\core_1.execute.sreg_scratch.o_d[9] ));
 sky130_fd_sc_hd__dfxtp_1 _7216_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0488_),
    .Q(\core_1.execute.sreg_scratch.o_d[10] ));
 sky130_fd_sc_hd__dfxtp_1 _7217_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0489_),
    .Q(\core_1.execute.sreg_scratch.o_d[11] ));
 sky130_fd_sc_hd__dfxtp_1 _7218_ (.CLK(clknet_leaf_21_i_clk),
    .D(_0490_),
    .Q(\core_1.execute.sreg_scratch.o_d[12] ));
 sky130_fd_sc_hd__dfxtp_1 _7219_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0491_),
    .Q(\core_1.execute.sreg_scratch.o_d[13] ));
 sky130_fd_sc_hd__dfxtp_1 _7220_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0492_),
    .Q(\core_1.execute.sreg_scratch.o_d[14] ));
 sky130_fd_sc_hd__dfxtp_1 _7221_ (.CLK(clknet_leaf_22_i_clk),
    .D(_0493_),
    .Q(\core_1.execute.sreg_scratch.o_d[15] ));
 sky130_fd_sc_hd__dfxtp_1 _7222_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0494_),
    .Q(\core_1.execute.sreg_irq_flags.o_d[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7223_ (.CLK(clknet_leaf_32_i_clk),
    .D(_0495_),
    .Q(\core_1.execute.sreg_irq_flags.o_d[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7224_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0496_),
    .Q(\core_1.execute.sreg_irq_flags.o_d[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7225_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0497_),
    .Q(\core_1.execute.sreg_irq_flags.o_d[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7226_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0498_),
    .Q(\core_1.execute.sreg_irq_flags.o_d[4] ));
 sky130_fd_sc_hd__dfxtp_2 _7227_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0499_),
    .Q(\core_1.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__dfxtp_2 _7228_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0500_),
    .Q(\core_1.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__dfxtp_2 _7229_ (.CLK(clknet_leaf_31_i_clk),
    .D(_0501_),
    .Q(\core_1.execute.pc_high_out[2] ));
 sky130_fd_sc_hd__dfxtp_2 _7230_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0502_),
    .Q(\core_1.execute.pc_high_out[3] ));
 sky130_fd_sc_hd__dfxtp_2 _7231_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0503_),
    .Q(\core_1.execute.pc_high_out[4] ));
 sky130_fd_sc_hd__dfxtp_2 _7232_ (.CLK(clknet_leaf_29_i_clk),
    .D(_0504_),
    .Q(\core_1.execute.pc_high_out[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7233_ (.CLK(clknet_leaf_30_i_clk),
    .D(_0505_),
    .Q(\core_1.execute.pc_high_out[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7234_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0506_),
    .Q(\core_1.execute.pc_high_out[7] ));
 sky130_fd_sc_hd__dfxtp_1 _7235_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0507_),
    .Q(\core_1.execute.pc_high_buff_out[0] ));
 sky130_fd_sc_hd__dfxtp_1 _7236_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0508_),
    .Q(\core_1.execute.pc_high_buff_out[1] ));
 sky130_fd_sc_hd__dfxtp_1 _7237_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0509_),
    .Q(\core_1.execute.pc_high_buff_out[2] ));
 sky130_fd_sc_hd__dfxtp_1 _7238_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0510_),
    .Q(\core_1.execute.pc_high_buff_out[3] ));
 sky130_fd_sc_hd__dfxtp_1 _7239_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0511_),
    .Q(\core_1.execute.pc_high_buff_out[4] ));
 sky130_fd_sc_hd__dfxtp_1 _7240_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0512_),
    .Q(\core_1.execute.pc_high_buff_out[5] ));
 sky130_fd_sc_hd__dfxtp_1 _7241_ (.CLK(clknet_leaf_28_i_clk),
    .D(_0513_),
    .Q(\core_1.execute.pc_high_buff_out[6] ));
 sky130_fd_sc_hd__dfxtp_1 _7242_ (.CLK(clknet_leaf_27_i_clk),
    .D(_0514_),
    .Q(\core_1.execute.pc_high_buff_out[7] ));
 sky130_fd_sc_hd__conb_1 core1_213 (.LO(net213));
 sky130_fd_sc_hd__conb_1 core1_214 (.LO(net214));
 sky130_fd_sc_hd__conb_1 core1_215 (.LO(net215));
 sky130_fd_sc_hd__conb_1 core1_216 (.LO(net216));
 sky130_fd_sc_hd__conb_1 core1_217 (.LO(net217));
 sky130_fd_sc_hd__conb_1 core1_218 (.LO(net218));
 sky130_fd_sc_hd__conb_1 core1_219 (.LO(net219));
 sky130_fd_sc_hd__conb_1 core1_220 (.LO(net220));
 sky130_fd_sc_hd__conb_1 core1_221 (.LO(net221));
 sky130_fd_sc_hd__conb_1 core1_222 (.LO(net222));
 sky130_fd_sc_hd__conb_1 core1_223 (.LO(net223));
 sky130_fd_sc_hd__conb_1 core1_224 (.LO(net224));
 sky130_fd_sc_hd__conb_1 core1_225 (.LO(net225));
 sky130_fd_sc_hd__conb_1 core1_226 (.LO(net226));
 sky130_fd_sc_hd__conb_1 core1_227 (.LO(net227));
 sky130_fd_sc_hd__conb_1 core1_228 (.LO(net228));
 sky130_fd_sc_hd__conb_1 core1_229 (.LO(net229));
 sky130_fd_sc_hd__conb_1 core1_230 (.LO(net230));
 sky130_fd_sc_hd__conb_1 core1_231 (.LO(net231));
 sky130_fd_sc_hd__conb_1 core1_232 (.LO(net232));
 sky130_fd_sc_hd__conb_1 core1_233 (.LO(net233));
 sky130_fd_sc_hd__conb_1 core1_234 (.LO(net234));
 sky130_fd_sc_hd__conb_1 core1_235 (.LO(net235));
 sky130_fd_sc_hd__conb_1 core1_236 (.LO(net236));
 sky130_fd_sc_hd__conb_1 core1_237 (.LO(net237));
 sky130_fd_sc_hd__conb_1 core1_238 (.LO(net238));
 sky130_fd_sc_hd__conb_1 core1_239 (.LO(net239));
 sky130_fd_sc_hd__conb_1 core1_240 (.LO(net240));
 sky130_fd_sc_hd__conb_1 core1_241 (.LO(net241));
 sky130_fd_sc_hd__conb_1 core1_242 (.LO(net242));
 sky130_fd_sc_hd__conb_1 core1_243 (.LO(net243));
 sky130_fd_sc_hd__conb_1 core1_244 (.LO(net244));
 sky130_fd_sc_hd__conb_1 core1_245 (.LO(net245));
 sky130_fd_sc_hd__conb_1 core1_246 (.LO(net246));
 sky130_fd_sc_hd__conb_1 core1_247 (.LO(net247));
 sky130_fd_sc_hd__conb_1 core1_248 (.LO(net248));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(i_core_int_sreg[0]),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(i_core_int_sreg[10]),
    .X(net2));
 sky130_fd_sc_hd__dlymetal6s2s_1 input3 (.A(i_core_int_sreg[11]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(i_core_int_sreg[12]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(i_core_int_sreg[13]),
    .X(net5));
 sky130_fd_sc_hd__buf_2 input6 (.A(i_core_int_sreg[14]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 input7 (.A(i_core_int_sreg[15]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(i_core_int_sreg[1]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(i_core_int_sreg[2]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(i_core_int_sreg[3]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(i_core_int_sreg[4]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(i_core_int_sreg[5]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(i_core_int_sreg[6]),
    .X(net13));
 sky130_fd_sc_hd__buf_2 input14 (.A(i_core_int_sreg[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(i_core_int_sreg[8]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(i_core_int_sreg[9]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(i_disable),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(i_irq),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(i_mc_core_int),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_4 input20 (.A(i_mem_ack),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(i_mem_data[0]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(i_mem_data[10]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(i_mem_data[11]),
    .X(net23));
 sky130_fd_sc_hd__dlymetal6s2s_1 input24 (.A(i_mem_data[12]),
    .X(net24));
 sky130_fd_sc_hd__dlymetal6s2s_1 input25 (.A(i_mem_data[13]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(i_mem_data[14]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 input27 (.A(i_mem_data[15]),
    .X(net27));
 sky130_fd_sc_hd__buf_2 input28 (.A(i_mem_data[1]),
    .X(net28));
 sky130_fd_sc_hd__buf_2 input29 (.A(i_mem_data[2]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input30 (.A(i_mem_data[3]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(i_mem_data[4]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(i_mem_data[5]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(i_mem_data[6]),
    .X(net33));
 sky130_fd_sc_hd__dlymetal6s2s_1 input34 (.A(i_mem_data[7]),
    .X(net34));
 sky130_fd_sc_hd__dlymetal6s2s_1 input35 (.A(i_mem_data[8]),
    .X(net35));
 sky130_fd_sc_hd__dlymetal6s2s_1 input36 (.A(i_mem_data[9]),
    .X(net36));
 sky130_fd_sc_hd__buf_6 input37 (.A(i_mem_exception),
    .X(net37));
 sky130_fd_sc_hd__dlymetal6s2s_1 input38 (.A(i_req_data[0]),
    .X(net38));
 sky130_fd_sc_hd__dlymetal6s2s_1 input39 (.A(i_req_data[10]),
    .X(net39));
 sky130_fd_sc_hd__dlymetal6s2s_1 input40 (.A(i_req_data[11]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(i_req_data[12]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_1 input42 (.A(i_req_data[13]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(i_req_data[14]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(i_req_data[15]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(i_req_data[16]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(i_req_data[17]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(i_req_data[18]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input48 (.A(i_req_data[19]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(i_req_data[1]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(i_req_data[20]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(i_req_data[21]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 input52 (.A(i_req_data[22]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 input53 (.A(i_req_data[23]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(i_req_data[24]),
    .X(net54));
 sky130_fd_sc_hd__dlymetal6s2s_1 input55 (.A(i_req_data[25]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 input56 (.A(i_req_data[26]),
    .X(net56));
 sky130_fd_sc_hd__dlymetal6s2s_1 input57 (.A(i_req_data[27]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(i_req_data[28]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(i_req_data[29]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(i_req_data[2]),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 input61 (.A(i_req_data[30]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 input62 (.A(i_req_data[31]),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 input63 (.A(i_req_data[3]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(i_req_data[4]),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 input65 (.A(i_req_data[5]),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 input66 (.A(i_req_data[6]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(i_req_data[7]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(i_req_data[8]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(i_req_data[9]),
    .X(net69));
 sky130_fd_sc_hd__buf_4 input70 (.A(i_req_data_valid),
    .X(net70));
 sky130_fd_sc_hd__buf_4 input71 (.A(i_rst),
    .X(net71));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(dbg_pc[0]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(dbg_pc[10]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(dbg_pc[11]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(dbg_pc[12]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(dbg_pc[13]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(dbg_pc[14]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(dbg_pc[15]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(dbg_pc[1]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(dbg_pc[2]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(dbg_pc[3]));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(dbg_pc[4]));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(dbg_pc[5]));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(dbg_pc[6]));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(dbg_pc[7]));
 sky130_fd_sc_hd__buf_2 output86 (.A(net86),
    .X(dbg_pc[8]));
 sky130_fd_sc_hd__buf_2 output87 (.A(net87),
    .X(dbg_pc[9]));
 sky130_fd_sc_hd__buf_2 output88 (.A(net88),
    .X(dbg_r0[0]));
 sky130_fd_sc_hd__buf_2 output89 (.A(net89),
    .X(dbg_r0[10]));
 sky130_fd_sc_hd__buf_2 output90 (.A(net90),
    .X(dbg_r0[11]));
 sky130_fd_sc_hd__buf_2 output91 (.A(net91),
    .X(dbg_r0[12]));
 sky130_fd_sc_hd__buf_2 output92 (.A(net92),
    .X(dbg_r0[13]));
 sky130_fd_sc_hd__buf_2 output93 (.A(net93),
    .X(dbg_r0[14]));
 sky130_fd_sc_hd__buf_2 output94 (.A(net94),
    .X(dbg_r0[15]));
 sky130_fd_sc_hd__buf_2 output95 (.A(net95),
    .X(dbg_r0[1]));
 sky130_fd_sc_hd__buf_2 output96 (.A(net96),
    .X(dbg_r0[2]));
 sky130_fd_sc_hd__buf_2 output97 (.A(net97),
    .X(dbg_r0[3]));
 sky130_fd_sc_hd__buf_2 output98 (.A(net98),
    .X(dbg_r0[4]));
 sky130_fd_sc_hd__buf_2 output99 (.A(net99),
    .X(dbg_r0[5]));
 sky130_fd_sc_hd__buf_2 output100 (.A(net100),
    .X(dbg_r0[6]));
 sky130_fd_sc_hd__buf_2 output101 (.A(net101),
    .X(dbg_r0[7]));
 sky130_fd_sc_hd__buf_2 output102 (.A(net102),
    .X(dbg_r0[8]));
 sky130_fd_sc_hd__buf_2 output103 (.A(net103),
    .X(dbg_r0[9]));
 sky130_fd_sc_hd__buf_2 output104 (.A(net104),
    .X(o_c_data_page));
 sky130_fd_sc_hd__buf_2 output105 (.A(net105),
    .X(o_c_instr_long));
 sky130_fd_sc_hd__buf_2 output106 (.A(net106),
    .X(o_c_instr_page));
 sky130_fd_sc_hd__buf_2 output107 (.A(net107),
    .X(o_icache_flush));
 sky130_fd_sc_hd__buf_2 output108 (.A(net108),
    .X(o_instr_long_addr[0]));
 sky130_fd_sc_hd__buf_2 output109 (.A(net109),
    .X(o_instr_long_addr[1]));
 sky130_fd_sc_hd__buf_2 output110 (.A(net110),
    .X(o_instr_long_addr[2]));
 sky130_fd_sc_hd__buf_2 output111 (.A(net111),
    .X(o_instr_long_addr[3]));
 sky130_fd_sc_hd__buf_2 output112 (.A(net112),
    .X(o_instr_long_addr[4]));
 sky130_fd_sc_hd__buf_2 output113 (.A(net113),
    .X(o_instr_long_addr[5]));
 sky130_fd_sc_hd__buf_2 output114 (.A(net114),
    .X(o_instr_long_addr[6]));
 sky130_fd_sc_hd__buf_2 output115 (.A(net115),
    .X(o_instr_long_addr[7]));
 sky130_fd_sc_hd__buf_2 output116 (.A(net116),
    .X(o_mem_addr[0]));
 sky130_fd_sc_hd__buf_2 output117 (.A(net117),
    .X(o_mem_addr[10]));
 sky130_fd_sc_hd__buf_2 output118 (.A(net118),
    .X(o_mem_addr[11]));
 sky130_fd_sc_hd__buf_2 output119 (.A(net119),
    .X(o_mem_addr[12]));
 sky130_fd_sc_hd__buf_2 output120 (.A(net120),
    .X(o_mem_addr[13]));
 sky130_fd_sc_hd__buf_2 output121 (.A(net121),
    .X(o_mem_addr[14]));
 sky130_fd_sc_hd__buf_2 output122 (.A(net122),
    .X(o_mem_addr[15]));
 sky130_fd_sc_hd__buf_2 output123 (.A(net123),
    .X(o_mem_addr[1]));
 sky130_fd_sc_hd__buf_2 output124 (.A(net124),
    .X(o_mem_addr[2]));
 sky130_fd_sc_hd__buf_2 output125 (.A(net125),
    .X(o_mem_addr[3]));
 sky130_fd_sc_hd__buf_2 output126 (.A(net126),
    .X(o_mem_addr[4]));
 sky130_fd_sc_hd__buf_2 output127 (.A(net127),
    .X(o_mem_addr[5]));
 sky130_fd_sc_hd__buf_2 output128 (.A(net128),
    .X(o_mem_addr[6]));
 sky130_fd_sc_hd__buf_2 output129 (.A(net129),
    .X(o_mem_addr[7]));
 sky130_fd_sc_hd__buf_2 output130 (.A(net130),
    .X(o_mem_addr[8]));
 sky130_fd_sc_hd__buf_2 output131 (.A(net131),
    .X(o_mem_addr[9]));
 sky130_fd_sc_hd__buf_2 output132 (.A(net132),
    .X(o_mem_addr_high[0]));
 sky130_fd_sc_hd__buf_2 output133 (.A(net133),
    .X(o_mem_addr_high[1]));
 sky130_fd_sc_hd__buf_2 output134 (.A(net134),
    .X(o_mem_addr_high[2]));
 sky130_fd_sc_hd__buf_2 output135 (.A(net135),
    .X(o_mem_addr_high[3]));
 sky130_fd_sc_hd__buf_2 output136 (.A(net136),
    .X(o_mem_addr_high[4]));
 sky130_fd_sc_hd__buf_2 output137 (.A(net137),
    .X(o_mem_addr_high[5]));
 sky130_fd_sc_hd__buf_2 output138 (.A(net138),
    .X(o_mem_addr_high[6]));
 sky130_fd_sc_hd__buf_2 output139 (.A(net139),
    .X(o_mem_data[0]));
 sky130_fd_sc_hd__buf_2 output140 (.A(net140),
    .X(o_mem_data[10]));
 sky130_fd_sc_hd__buf_2 output141 (.A(net141),
    .X(o_mem_data[11]));
 sky130_fd_sc_hd__buf_2 output142 (.A(net142),
    .X(o_mem_data[12]));
 sky130_fd_sc_hd__buf_2 output143 (.A(net143),
    .X(o_mem_data[13]));
 sky130_fd_sc_hd__buf_2 output144 (.A(net144),
    .X(o_mem_data[14]));
 sky130_fd_sc_hd__buf_2 output145 (.A(net145),
    .X(o_mem_data[15]));
 sky130_fd_sc_hd__buf_2 output146 (.A(net146),
    .X(o_mem_data[1]));
 sky130_fd_sc_hd__buf_2 output147 (.A(net147),
    .X(o_mem_data[2]));
 sky130_fd_sc_hd__buf_2 output148 (.A(net148),
    .X(o_mem_data[3]));
 sky130_fd_sc_hd__buf_2 output149 (.A(net149),
    .X(o_mem_data[4]));
 sky130_fd_sc_hd__buf_2 output150 (.A(net150),
    .X(o_mem_data[5]));
 sky130_fd_sc_hd__buf_2 output151 (.A(net151),
    .X(o_mem_data[6]));
 sky130_fd_sc_hd__buf_2 output152 (.A(net152),
    .X(o_mem_data[7]));
 sky130_fd_sc_hd__buf_2 output153 (.A(net153),
    .X(o_mem_data[8]));
 sky130_fd_sc_hd__buf_2 output154 (.A(net154),
    .X(o_mem_data[9]));
 sky130_fd_sc_hd__buf_2 output155 (.A(net155),
    .X(o_mem_long));
 sky130_fd_sc_hd__buf_2 output156 (.A(net156),
    .X(o_mem_req));
 sky130_fd_sc_hd__buf_2 output157 (.A(net157),
    .X(o_mem_sel[0]));
 sky130_fd_sc_hd__buf_2 output158 (.A(net158),
    .X(o_mem_sel[1]));
 sky130_fd_sc_hd__buf_2 output159 (.A(net159),
    .X(o_mem_we));
 sky130_fd_sc_hd__buf_2 output160 (.A(net160),
    .X(o_req_active));
 sky130_fd_sc_hd__buf_2 output161 (.A(net161),
    .X(o_req_addr[0]));
 sky130_fd_sc_hd__buf_2 output162 (.A(net162),
    .X(o_req_addr[10]));
 sky130_fd_sc_hd__buf_2 output163 (.A(net163),
    .X(o_req_addr[11]));
 sky130_fd_sc_hd__buf_2 output164 (.A(net164),
    .X(o_req_addr[12]));
 sky130_fd_sc_hd__buf_2 output165 (.A(net165),
    .X(o_req_addr[13]));
 sky130_fd_sc_hd__buf_2 output166 (.A(net166),
    .X(o_req_addr[14]));
 sky130_fd_sc_hd__buf_2 output167 (.A(net167),
    .X(o_req_addr[15]));
 sky130_fd_sc_hd__buf_2 output168 (.A(net168),
    .X(o_req_addr[1]));
 sky130_fd_sc_hd__buf_2 output169 (.A(net169),
    .X(o_req_addr[2]));
 sky130_fd_sc_hd__buf_2 output170 (.A(net170),
    .X(o_req_addr[3]));
 sky130_fd_sc_hd__buf_2 output171 (.A(net171),
    .X(o_req_addr[4]));
 sky130_fd_sc_hd__buf_2 output172 (.A(net172),
    .X(o_req_addr[5]));
 sky130_fd_sc_hd__buf_2 output173 (.A(net173),
    .X(o_req_addr[6]));
 sky130_fd_sc_hd__buf_2 output174 (.A(net174),
    .X(o_req_addr[7]));
 sky130_fd_sc_hd__buf_2 output175 (.A(net175),
    .X(o_req_addr[8]));
 sky130_fd_sc_hd__buf_2 output176 (.A(net176),
    .X(o_req_addr[9]));
 sky130_fd_sc_hd__buf_2 output177 (.A(net177),
    .X(o_req_ppl_submit));
 sky130_fd_sc_hd__buf_2 output178 (.A(net211),
    .X(sr_bus_addr[0]));
 sky130_fd_sc_hd__buf_2 output179 (.A(net179),
    .X(sr_bus_addr[10]));
 sky130_fd_sc_hd__buf_2 output180 (.A(net180),
    .X(sr_bus_addr[11]));
 sky130_fd_sc_hd__buf_2 output181 (.A(net181),
    .X(sr_bus_addr[12]));
 sky130_fd_sc_hd__buf_2 output182 (.A(net182),
    .X(sr_bus_addr[13]));
 sky130_fd_sc_hd__buf_2 output183 (.A(net183),
    .X(sr_bus_addr[14]));
 sky130_fd_sc_hd__buf_2 output184 (.A(net184),
    .X(sr_bus_addr[15]));
 sky130_fd_sc_hd__buf_2 output185 (.A(net185),
    .X(sr_bus_addr[1]));
 sky130_fd_sc_hd__buf_2 output186 (.A(net186),
    .X(sr_bus_addr[2]));
 sky130_fd_sc_hd__buf_2 output187 (.A(net187),
    .X(sr_bus_addr[3]));
 sky130_fd_sc_hd__buf_2 output188 (.A(net188),
    .X(sr_bus_addr[4]));
 sky130_fd_sc_hd__buf_2 output189 (.A(net189),
    .X(sr_bus_addr[5]));
 sky130_fd_sc_hd__buf_2 output190 (.A(net190),
    .X(sr_bus_addr[6]));
 sky130_fd_sc_hd__buf_2 output191 (.A(net191),
    .X(sr_bus_addr[7]));
 sky130_fd_sc_hd__buf_2 output192 (.A(net192),
    .X(sr_bus_addr[8]));
 sky130_fd_sc_hd__buf_2 output193 (.A(net193),
    .X(sr_bus_addr[9]));
 sky130_fd_sc_hd__buf_2 output194 (.A(net194),
    .X(sr_bus_data_o[0]));
 sky130_fd_sc_hd__buf_2 output195 (.A(net195),
    .X(sr_bus_data_o[10]));
 sky130_fd_sc_hd__buf_2 output196 (.A(net196),
    .X(sr_bus_data_o[11]));
 sky130_fd_sc_hd__buf_2 output197 (.A(net197),
    .X(sr_bus_data_o[12]));
 sky130_fd_sc_hd__buf_2 output198 (.A(net198),
    .X(sr_bus_data_o[13]));
 sky130_fd_sc_hd__buf_2 output199 (.A(net199),
    .X(sr_bus_data_o[14]));
 sky130_fd_sc_hd__buf_2 output200 (.A(net200),
    .X(sr_bus_data_o[15]));
 sky130_fd_sc_hd__buf_2 output201 (.A(net201),
    .X(sr_bus_data_o[1]));
 sky130_fd_sc_hd__buf_2 output202 (.A(net202),
    .X(sr_bus_data_o[2]));
 sky130_fd_sc_hd__buf_2 output203 (.A(net203),
    .X(sr_bus_data_o[3]));
 sky130_fd_sc_hd__buf_2 output204 (.A(net204),
    .X(sr_bus_data_o[4]));
 sky130_fd_sc_hd__buf_2 output205 (.A(net205),
    .X(sr_bus_data_o[5]));
 sky130_fd_sc_hd__buf_2 output206 (.A(net206),
    .X(sr_bus_data_o[6]));
 sky130_fd_sc_hd__buf_2 output207 (.A(net207),
    .X(sr_bus_data_o[7]));
 sky130_fd_sc_hd__buf_2 output208 (.A(net208),
    .X(sr_bus_data_o[8]));
 sky130_fd_sc_hd__buf_2 output209 (.A(net209),
    .X(sr_bus_data_o[9]));
 sky130_fd_sc_hd__buf_2 output210 (.A(net210),
    .X(sr_bus_we));
 sky130_fd_sc_hd__buf_4 fanout211 (.A(net178),
    .X(net211));
 sky130_fd_sc_hd__conb_1 core1_212 (.LO(net212));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_i_clk (.A(i_clk),
    .X(clknet_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_1_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_1_i_clk (.A(clknet_1_0_0_i_clk),
    .X(clknet_1_0_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_1_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_1_i_clk (.A(clknet_1_1_0_i_clk),
    .X(clknet_1_1_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_i_clk (.A(clknet_1_0_1_i_clk),
    .X(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_i_clk (.A(clknet_1_0_1_i_clk),
    .X(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_i_clk (.A(clknet_1_1_1_i_clk),
    .X(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_i_clk (.A(clknet_1_1_1_i_clk),
    .X(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6726__D (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4089__A2 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4074__A2 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4072__A2 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__A2 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4056__A2 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__A2 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__A2 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4025__A2 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__A2 (.DIODE(_0015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6826__D (.DIODE(_0115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__D (.DIODE(_0228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__B (.DIODE(_0228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__B (.DIODE(_0228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__B (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__B (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__B (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__A2_N (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3425__B (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3418__A2 (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3409__B1 (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3401__B (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3333__A (.DIODE(_0516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4378__A2 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__A2 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__A2 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__B1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__B1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3456__B1 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3393__B (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__A2 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3369__B (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3361__A2 (.DIODE(_0517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__A2 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__A2 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3452__A2 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__A2 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__B1 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3421__A2 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3397__A2 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3389__A2 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__A2 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3345__A2 (.DIODE(_0519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3465__B (.DIODE(_0525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__B1 (.DIODE(_0525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3344__A2 (.DIODE(_0525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__A2 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__A2 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__A2 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__A2 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__A2 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__A2 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3396__A2 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__A2 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3364__A2 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3344__B1 (.DIODE(_0527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__B1 (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__B1 (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__B1 (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__B1 (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3452__B1 (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__B1 (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__B1 (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3389__B1 (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3368__B1 (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3360__A2 (.DIODE(_0532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4058__A1 (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3555__A1 (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3461__B (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3460__A_N (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__B (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3390__A_N (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3382__B (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__A_N (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3378__D (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3351__A (.DIODE(_0534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3554__A (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3355__A2 (.DIODE(_0535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__A2 (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3462__A2 (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__A2 (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__B1 (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__A2 (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3417__A2 (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__A2 (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__A2 (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3368__A2 (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__A2 (.DIODE(_0541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__A2 (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__A2 (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__B1 (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__B1 (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3367__A2 (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__B1 (.DIODE(_0542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__A1 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6571__A (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__A1 (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4147__B (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3362__A (.DIODE(_0545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__A1 (.DIODE(_0553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6567__A (.DIODE(_0553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6437__A1 (.DIODE(_0553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4143__A1_N (.DIODE(_0553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3371__A (.DIODE(_0553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__B1 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__B1 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__B1 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__A2 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3420__B1 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3414__A2 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3404__B1 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3396__B1 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__B1 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__A2 (.DIODE(_0554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4056__A1 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__S1 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__S1 (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3461__D (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__D (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3390__C (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3382__D (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3378__B (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3377__A_N (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3375__B_N (.DIODE(_0555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4054__A1 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__S0 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__S0 (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3461__C (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__C (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3390__B (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3382__C (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__B (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3378__A_N (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3377__B (.DIODE(_0558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3478__D1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3462__D1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3455__D1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__C1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__C1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3434__D1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3424__D1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3417__D1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__D1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__D1 (.DIODE(_0566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6625__A1 (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6563__A (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__B (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3387__A (.DIODE(_0568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__A1 (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__A1 (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4424__A2 (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4137__A1_N (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3395__A (.DIODE(_0575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__A1 (.DIODE(_0582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6554__A (.DIODE(_0582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__A1 (.DIODE(_0582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__A1 (.DIODE(_0582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__A1_N (.DIODE(_0582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3403__A (.DIODE(_0582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__A1 (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6550__A (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6405__A1 (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__A1_N (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3410__A (.DIODE(_0588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__A1 (.DIODE(_0596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__A (.DIODE(_0596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6399__A1 (.DIODE(_0596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__A2 (.DIODE(_0596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__A1_N (.DIODE(_0596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3419__A (.DIODE(_0596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6615__A1 (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6542__A (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A1 (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__A1_N (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3427__A (.DIODE(_0603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6723__A (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6613__A1 (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6538__A (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6385__A1 (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__A1_N (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3436__A (.DIODE(_0611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__A1 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__A1 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6534__A (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6378__A1 (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__A1_N (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3443__A (.DIODE(_0617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__A1 (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6530__A (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__A1 (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4519__A2 (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4413__A2 (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4115__B (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3450__A (.DIODE(_0623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__A1 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__A1 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6526__A (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__A1 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__A2 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__A2 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__A2 (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4111__A1_N (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3457__A (.DIODE(_0629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__A1 (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6521__A (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6476__A1 (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6355__A1 (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4462__A2 (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4417__A2 (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__A1_N (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3464__A (.DIODE(_0635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__A1 (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6602__A1 (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6517__A (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6470__A1 (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6351__A (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__B (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__A1 (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3473__A (.DIODE(_0643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__A1 (.DIODE(_0644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3480__A1 (.DIODE(_0644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__A3 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3480__A3 (.DIODE(_0648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6600__A1 (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__A (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6467__A1 (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__A1 (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__A1_N (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3481__A (.DIODE(_0650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4378__B1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__B1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__B1 (.DIODE(_0652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4378__B2 (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__B2 (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__B2 (.DIODE(_0657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6598__A1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6506__A (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6465__A1 (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__A (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3490__A (.DIODE(_0658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6597__A (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__A (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__A (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__B (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4163__A (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__B (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4116__A (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__A (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3948__A (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3611__A (.DIODE(_0659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3599__S (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3597__A1 (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3595__A1 (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3592__A1 (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3591__B_N (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3588__S (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3583__S (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3572__S (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__S (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3495__A (.DIODE(_0662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__S (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3767__S (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3766__S (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__A1 (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3606__S (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3605__S (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3604__S (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3575__S (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3574__S (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3496__A (.DIODE(_0663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4353__S (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4304__S (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4301__S (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4298__S (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4295__S (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__S (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4232__B1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3892__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3769__S (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__A1 (.DIODE(_0664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6575__B1 (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6100__B (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4098__B (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__A (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3500__A (.DIODE(_0667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6574__C (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6507__B1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6500__B1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__C1 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__A (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3941__A2 (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__A (.DIODE(_0668_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__A1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6645__A (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__A1 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__A (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6590__B2 (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__B (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3512__B (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__B (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__B (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3503__B (.DIODE(_0670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__C1 (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3520__B (.DIODE(_0687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__B (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__A2 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__B (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__A2 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4433__A (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4430__A (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3545__C1 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3541__A1 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3537__A (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3536__C1 (.DIODE(_0693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__A (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__B (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4569__A (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__A (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__B (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__B (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4450__B1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4386__B1 (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3533__A (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__A (.DIODE(_0694_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__C (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__C (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__C (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4025__A1 (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__C_N (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__C_N (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__B (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__S1 (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__B1 (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3528__B (.DIODE(_0695_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__C (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__C (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__B (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__A_N (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__C (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__B (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__B (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4384__A_N (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3532__B (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3531__A_N (.DIODE(_0698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__B2 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__B2 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__B1 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__B2 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__B2 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4514__B2 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__B1 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__B2 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4395__B (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3535__A2 (.DIODE(_0700_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4610__B1 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4603__A1 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__B2 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__B (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4023__A1 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__A (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__A (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3542__A (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__S0 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__A1 (.DIODE(_0701_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__A1 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3540__B1 (.DIODE(_0707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4595__B (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4578__B (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4563__B (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4449__A_N (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__B (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__B (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4388__C_N (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4387__A (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4385__A_N (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3549__A (.DIODE(_0716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4607__B (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__B (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4585__B_N (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4532__B_N (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__B_N (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__B_N (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4434__A (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4429__A (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4027__A1 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__C1 (.DIODE(_0717_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3556__B2 (.DIODE(_0723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__A (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3897__A (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3565__B (.DIODE(_0724_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6295__B (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__S (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__B (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__B (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__A (.DIODE(_0726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6264__B (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__A1 (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6150__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6125__A (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3562__B (.DIODE(_0729_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__D_N (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__D_N (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3935__C (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3564__B (.DIODE(_0731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__B (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3651__B1 (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3568__A (.DIODE(_0735_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__A0 (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3582__D_N (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3573__A (.DIODE(_0739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__A0 (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__D_N (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3582__A (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3573__B_N (.DIODE(_0740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4273__A0 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__B1 (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__A (.DIODE(_0742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__A0 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3603__C1 (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3576__B (.DIODE(_0743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__A0 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__A1 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__A2 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__A2 (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__A (.DIODE(_0746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__A0 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__A1 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__B1 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__A2 (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__B (.DIODE(_0747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4328__A0 (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__A1 (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3751__A2 (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__B1 (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3582__B (.DIODE(_0748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__A0 (.DIODE(_0749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A1 (.DIODE(_0749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3756__A2 (.DIODE(_0749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__A1_N (.DIODE(_0749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3582__C (.DIODE(_0749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__A0 (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__A1 (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__A2 (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3728__A2_N (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__A (.DIODE(_0751_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__A0 (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__A1 (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__A2 (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3742__B1 (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__B (.DIODE(_0752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__A0 (.DIODE(_0753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__A1 (.DIODE(_0753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3741__B1 (.DIODE(_0753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3740__A2 (.DIODE(_0753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__C (.DIODE(_0753_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4322__A0 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__B1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__B1 (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3587__D (.DIODE(_0754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__A0 (.DIODE(_0756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__A1 (.DIODE(_0756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3761__A2 (.DIODE(_0756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3760__A2 (.DIODE(_0756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__A (.DIODE(_0756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4307__A0 (.DIODE(_0757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__A1 (.DIODE(_0757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3739__B1 (.DIODE(_0757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__B (.DIODE(_0757_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4318__A0 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__A1 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__B1 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3743__B1 (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3593__C (.DIODE(_0758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__A0 (.DIODE(_0763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__A1 (.DIODE(_0763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__A (.DIODE(_0763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__A0 (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__A1 (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__B (.DIODE(_0765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__A0 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__A1 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3745__A2 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3744__A2 (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__C (.DIODE(_0766_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__A0 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__A1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3763__B1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3761__B1 (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3600__D (.DIODE(_0767_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3602__D (.DIODE(_0769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4277__A0 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3772__A (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3608__B1 (.DIODE(_0772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4281__A0 (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__B (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3607__A (.DIODE(_0773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__A0 (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3771__C (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3607__B (.DIODE(_0774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__C1 (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__C1 (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__C1 (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__C1 (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__C1 (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__C1 (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3779__A (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3610__C1 (.DIODE(_0777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4266__S (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4264__S (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4262__S (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4260__S (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4258__S (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4256__S (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4254__S (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4252__S (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3612__A (.DIODE(_0779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6454__A1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5657__A1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5620__A1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__A1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5545__B1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__A1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5436__A1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__A1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5066__C1 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__A0 (.DIODE(_0780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4033__A1 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4006__B1 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3999__A (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__B2 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3704__A (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3692__A2 (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3683__A (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3669__B (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3647__A (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__A (.DIODE(_0799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4086__A (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__A1 (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3699__A (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3642__B (.DIODE(_0800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__A (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__A (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4030__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4001__B1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3995__B1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__B1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3715__B1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3702__A (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3700__A (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__A1 (.DIODE(_0803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__A1 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__A2 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__A2 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4018__A2 (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3648__B1_N (.DIODE(_0806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__A1 (.DIODE(_0808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4081__B (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__A (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__A (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4059__B (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3990__C1 (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3989__A (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3674__A (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3662__A (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3657__A (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3652__A (.DIODE(_0810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4842__S (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__S (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4075__S (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4069__S (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__S (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4034__B1 (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3976__A (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3955__A (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3653__A (.DIODE(_0811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__A2 (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__A2 (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3991__A2 (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3954__A (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3722__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3693__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3654__S (.DIODE(_0812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__B2 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__B2 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__A1 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__B2 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__A1 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__B1 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__B1 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__A1 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__A1 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__A1 (.DIODE(_0814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__C1 (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__C1 (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__C1 (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__C1 (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__B1 (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__C1 (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__C1 (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__C1 (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3669__A (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3658__A (.DIODE(_0815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4064__A2 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4046__B1 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__B1 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4038__A2 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__A2 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__A2 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__A2 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__A2 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__A2 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__A2 (.DIODE(_0816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__B2 (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__B1 (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__B1 (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__B1 (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__A2 (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3664__B1 (.DIODE(_0820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__A1 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__A1 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__A1 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__A1 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__A1 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__A1 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4471__A (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__A1 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__A1 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3670__A1 (.DIODE(_0822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__A2 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__A2 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__A2 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__A2 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__A2 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__B1 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__B1 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__A2 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__B1 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__B1 (.DIODE(_0830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__C1 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__C1 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__C1 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__C1 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5469__C1 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5402__C1 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__C1 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5291__C1 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__C1 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__B2 (.DIODE(_0831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__A1 (.DIODE(_0832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__B2 (.DIODE(_0832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__A1 (.DIODE(_0832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__B2 (.DIODE(_0832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5461__A1 (.DIODE(_0832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5433__B2 (.DIODE(_0832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5354__A1 (.DIODE(_0832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__B2 (.DIODE(_0832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5159__A1 (.DIODE(_0832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3680__A1 (.DIODE(_0832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__A2 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5624__A2 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__A2 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__A2 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__A2 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__A2 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__A2 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__A2 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__A2 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__A0 (.DIODE(_0835_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__C1 (.DIODE(_0837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3684__A1 (.DIODE(_0837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5679__A1 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5648__A1 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5553__B2 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5524__A1 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5434__A1 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__A1 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__A1 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5318__A1 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__A1 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3691__A1 (.DIODE(_0839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__A1 (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__A1 (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A1 (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__A1 (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__A1 (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__A1 (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__A1 (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__B1 (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__A1 (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3707__A0 (.DIODE(_0846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__A1 (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__A (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__A1 (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__A (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__A1 (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__A (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__A1 (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__A1 (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__A1 (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3710__A (.DIODE(_0859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__C1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__B (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__A1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__A1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__A1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5498__A1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__A (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5328__A1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5241__A1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__A1 (.DIODE(_0860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4048__C1 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3712__B2 (.DIODE(_0861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5677__A1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5652__A1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5454__A (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5398__B1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__A1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__B2 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__A1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5034__B1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__B1 (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3714__A (.DIODE(_0862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__A1 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6474__A1 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5621__A1 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A1 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5558__A (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5529__A1 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__A1 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5353__A (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__C1 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3716__A0 (.DIODE(_0863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__A2 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__A2 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__B (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__A2 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__B1 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__B1 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__A2 (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__B (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3725__A (.DIODE(_0870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__A2 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__A2 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__A2 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__A2 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__A2 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__A2 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__A2 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__A2 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A2 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__A2 (.DIODE(_0871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3759__A1 (.DIODE(_0891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3750__B (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3749__A2_N (.DIODE(_0893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3757__A2 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3755__A2_N (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3754__B2 (.DIODE(_0899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4287__A0 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__A1 (.DIODE(_0912_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__A0 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__A2 (.DIODE(_0913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__A0 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__A3 (.DIODE(_0914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__A0 (.DIODE(_0915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3770__A4 (.DIODE(_0915_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3773__A2 (.DIODE(_0916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3773__B1 (.DIODE(_0918_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3844__B1_N (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3822__A1 (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3817__A1 (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3774__A (.DIODE(_0919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__A1 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__A2 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__A2 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3835__S (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__A2 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3826__A (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3789__A (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3783__S (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3777__A (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__A2 (.DIODE(_0920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3849__B1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3845__C1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__B1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3827__B1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3781__A (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3776__B1 (.DIODE(_0921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__B1 (.DIODE(_0922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3848__A (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3840__A (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3831__A (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3812__A (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3808__A (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3803__A (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3798__A (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3794__A (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3788__A (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3778__B (.DIODE(_0923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__C1 (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__C1 (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__C1 (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__C1 (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__C1 (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__C1 (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__C1 (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__C1 (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__C1 (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__C1 (.DIODE(_0925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__C (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3837__A1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__B1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__B1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__B1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__B1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__B1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__B1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__B1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3785__A1 (.DIODE(_0926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3841__A2 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3832__A2 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3823__A2 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3818__A2 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3813__A2 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3809__A2 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3804__A2 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3799__A2 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3795__A2 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3790__A2 (.DIODE(_0933_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__S (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__S (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__S (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__S (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__S (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__S (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__S (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__S (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__S (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3855__A (.DIODE(_0983_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3889__A (.DIODE(_1000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4338__S (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4336__S (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4315__A (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4289__A (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4268__A (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3893__A (.DIODE(_1002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3895__A (.DIODE(_1003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6101__A1 (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__C (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4899__B (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4883__B (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4881__B (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4879__B (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4877__B (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4875__B (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4873__B (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3899__A (.DIODE(_1006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4869__B (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4867__B (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4865__B (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4863__B (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4861__B (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4859__B (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4857__B (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4855__B (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4853__B (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3947__A1 (.DIODE(_1007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__B (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__B (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__B (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__A1 (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__A (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__A (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__A_N (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5122__A (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__A (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3909__A (.DIODE(_1009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5124__C (.DIODE(_1010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__A0 (.DIODE(_1010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__B (.DIODE(_1010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__C (.DIODE(_1011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__B (.DIODE(_1011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__C (.DIODE(_1011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__B (.DIODE(_1011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__C (.DIODE(_1011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__B (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__C (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__C (.DIODE(_1013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__C (.DIODE(_1014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3943__C (.DIODE(_1014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__D (.DIODE(_1014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__B (.DIODE(_1015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5132__B (.DIODE(_1015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3908__A (.DIODE(_1015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__B (.DIODE(_1017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__A2 (.DIODE(_1017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__A2 (.DIODE(_1017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__A2 (.DIODE(_1017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5448__B (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5415__B (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5377__B (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__B (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5303__B (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5266__A1 (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5265__B (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5253__A1 (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__A1 (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3911__A (.DIODE(_1018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5643__A1 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5642__B (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5579__B (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5568__B1 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5563__B (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5514__B (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5500__B (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5449__A1 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4093__A (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__B1 (.DIODE(_1019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6421__A1 (.DIODE(_1043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6367__A1 (.DIODE(_1043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__B (.DIODE(_1043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4847__A (.DIODE(_1043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3937__A (.DIODE(_1043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6645__B (.DIODE(_1045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6641__B (.DIODE(_1045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3938__B (.DIODE(_1045_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6590__A2 (.DIODE(_1047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__A2 (.DIODE(_1047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3940__B (.DIODE(_1047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__A2 (.DIODE(_1051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__B (.DIODE(_1053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3946__C_N (.DIODE(_1053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__B1 (.DIODE(_1055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__B1 (.DIODE(_1055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6625__B1 (.DIODE(_1055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__B1 (.DIODE(_1055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__B1 (.DIODE(_1055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__B1 (.DIODE(_1055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__B1 (.DIODE(_1055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4345__A (.DIODE(_1055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4340__A (.DIODE(_1055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3949__A (.DIODE(_1055_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6295__A (.DIODE(_1056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4891__A (.DIODE(_1056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4890__A (.DIODE(_1056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4889__A (.DIODE(_1056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4888__A (.DIODE(_1056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4887__A (.DIODE(_1056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4886__A (.DIODE(_1056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4885__A (.DIODE(_1056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4634__A (.DIODE(_1056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3950__A (.DIODE(_1056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6648__A (.DIODE(_1057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__A (.DIODE(_1057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6575__A2 (.DIODE(_1057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6574__B (.DIODE(_1057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6499__A (.DIODE(_1057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6453__A (.DIODE(_1057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__B (.DIODE(_1057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__B (.DIODE(_1057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4077__A0 (.DIODE(_1057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__B (.DIODE(_1057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3953__A (.DIODE(_1058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__S (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__S (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__S (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__S (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__S (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__S (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__S (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__S (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__S (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__S (.DIODE(_1059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__S (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4014__S (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4011__S (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4003__S (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__S (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__S (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__S (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__S (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__S (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__S (.DIODE(_1070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__B (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__A2 (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__A2 (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__A2 (.DIODE(_1104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4071__C (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4050__B (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__B1 (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__B1 (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__B1 (.DIODE(_1105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__B (.DIODE(_1115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__B (.DIODE(_1115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__B (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__A2 (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__A2 (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__A2 (.DIODE(_1122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4073__C (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__B1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__B1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__B1 (.DIODE(_1125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__B2 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__B2 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__B2 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5567__A (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__B2 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__B2 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__B2 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__B2 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5207__A1 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4082__A1 (.DIODE(_1138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__A (.DIODE(_1141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6099__A (.DIODE(_1141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5691__S (.DIODE(_1141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5630__S (.DIODE(_1141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5580__A1 (.DIODE(_1141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5515__A1 (.DIODE(_1141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5504__A (.DIODE(_1141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4359__A (.DIODE(_1141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4095__A (.DIODE(_1141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4085__A1 (.DIODE(_1141_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__A2 (.DIODE(_1144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__A2 (.DIODE(_1144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5299__A2 (.DIODE(_1144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A2 (.DIODE(_1144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A2 (.DIODE(_1144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__A2 (.DIODE(_1144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__A2 (.DIODE(_1144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4092__A (.DIODE(_1144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__A2 (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__A2 (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__A2 (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__A2 (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__A2 (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__A2 (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__A2 (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__A2 (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__A2 (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__A3 (.DIODE(_1145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6446__A2 (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__A2 (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6340__A (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5251__A1 (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5146__A1 (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4362__A (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4147__A (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__A (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4115__A (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__B1 (.DIODE(_1146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4143__A2_N (.DIODE(_1148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4137__A2_N (.DIODE(_1148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4133__A2_N (.DIODE(_1148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4130__A2_N (.DIODE(_1148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4127__A2_N (.DIODE(_1148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4099__A (.DIODE(_1148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4096__B (.DIODE(_1148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4146__B (.DIODE(_1150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4140__B (.DIODE(_1150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__B1 (.DIODE(_1150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__B1 (.DIODE(_1150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__B1 (.DIODE(_1150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4114__B (.DIODE(_1150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4111__B1 (.DIODE(_1150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__B1 (.DIODE(_1150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__B1 (.DIODE(_1150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4101__A2 (.DIODE(_1150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4147__C (.DIODE(_1152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4141__C (.DIODE(_1152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4124__A2_N (.DIODE(_1152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4121__A2_N (.DIODE(_1152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4118__A2_N (.DIODE(_1152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4115__C (.DIODE(_1152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4111__A2_N (.DIODE(_1152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__A2_N (.DIODE(_1152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4105__A2_N (.DIODE(_1152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4100__B (.DIODE(_1152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6631__A (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6556__A (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6514__A (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6089__A (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6067__A (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6042__A (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6018__A (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4870__A (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4849__A (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4104__A (.DIODE(_1155_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__B1 (.DIODE(_1156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4134__A (.DIODE(_1156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4131__A (.DIODE(_1156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4128__A (.DIODE(_1156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4125__A (.DIODE(_1156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4122__A (.DIODE(_1156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4119__A (.DIODE(_1156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4112__A (.DIODE(_1156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4109__A (.DIODE(_1156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4106__A (.DIODE(_1156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6725__C1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__C1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6676__C1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6664__C1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6586__B1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5754__A (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4892__A (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4148__B1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4142__B1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4117__B1 (.DIODE(_1165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6591__A (.DIODE(_1178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6588__A (.DIODE(_1178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6583__A (.DIODE(_1178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6580__A (.DIODE(_1178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6577__A (.DIODE(_1178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4845__A (.DIODE(_1178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4351__A (.DIODE(_1178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4343__A (.DIODE(_1178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4144__A (.DIODE(_1178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4138__A (.DIODE(_1178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6220__C1 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__A1 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6199__A1 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6198__B (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6186__A (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6179__A (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6158__A1 (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6157__B (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6154__B (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4150__A (.DIODE(_1187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6319__A (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6245__A (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6232__A (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__C1 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6122__A (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__A1 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4823__B2 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__C1 (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4708__A (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4158__A (.DIODE(_1188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6244__S (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6231__A1 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6230__A (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__A1 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6197__S (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6178__S (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__B2 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6153__A (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6146__A2 (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4153__A (.DIODE(_1190_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__A (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6334__A (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6315__A (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6313__A (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6268__S1 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6256__S (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__C1 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__C1 (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4807__A (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4157__A (.DIODE(_1191_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__S0 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6217__S (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__S0 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__S (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6109__A (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6106__A1 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__S0 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__S0 (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__S (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__A (.DIODE(_1192_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__A1 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6243__A1 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__S1 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__B (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__A (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__S1 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__S1 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__A1 (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__B (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4156__B (.DIODE(_1193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__B (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__A1 (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6117__B2 (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__A1 (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__A1 (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4157__B (.DIODE(_1194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4796__A (.DIODE(_1196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4766__A (.DIODE(_1196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4755__A (.DIODE(_1196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4728__A (.DIODE(_1196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__A (.DIODE(_1196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4691__A1 (.DIODE(_1196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4159__A (.DIODE(_1196_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6297__A (.DIODE(_1197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__A1 (.DIODE(_1197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4795__A (.DIODE(_1197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4785__A1 (.DIODE(_1197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4736__A1 (.DIODE(_1197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4722__A1 (.DIODE(_1197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__A1 (.DIODE(_1197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__A (.DIODE(_1197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4694__A1 (.DIODE(_1197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__A2 (.DIODE(_1197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4836__B (.DIODE(_1198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4161__B1_N (.DIODE(_1198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4234__S (.DIODE(_1201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4230__S (.DIODE(_1201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4228__S (.DIODE(_1201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4207__A (.DIODE(_1201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4186__A (.DIODE(_1201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4165__A (.DIODE(_1201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4184__S (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4182__S (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4180__S (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4178__S (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4176__S (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4174__S (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4172__S (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4170__S (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4168__S (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__S (.DIODE(_1202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4205__S (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4203__S (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4201__S (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4199__S (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4197__S (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4195__S (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4193__S (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4191__S (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4189__S (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__S (.DIODE(_1213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4226__S (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4224__S (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4222__S (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4220__S (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4218__S (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4216__S (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4214__S (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4212__S (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4210__S (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4208__S (.DIODE(_1224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4287__S (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__S (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__S (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4281__S (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4279__S (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4277__S (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4275__S (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4273__S (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__S (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__S (.DIODE(_1255_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4313__S (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4311__S (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4309__S (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4307__S (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__S (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__S (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__S (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__S (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__S (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__S (.DIODE(_1266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4334__S (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4332__S (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4330__S (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4328__S (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4326__S (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4324__S (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4322__S (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4320__S (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4318__S (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4316__S (.DIODE(_1282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__B (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__S (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__S (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__S (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__S (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__S (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__S (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__S (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__S (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4349__A (.DIODE(_1299_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__B2 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__B2 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__B2 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__B2 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__B2 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__B2 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__B2 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__B2 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__A0 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4350__A1 (.DIODE(_1300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6421__A2 (.DIODE(_1305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6367__A2 (.DIODE(_1305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4357__B (.DIODE(_1305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6446__C1 (.DIODE(_1306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__C1 (.DIODE(_1306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6375__C1 (.DIODE(_1306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6356__A (.DIODE(_1306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4631__A (.DIODE(_1306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4358__A (.DIODE(_1306_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6432__B1 (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6409__B1 (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6402__A (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6389__B1 (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6382__B1 (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6373__B1 (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6361__B1 (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__A1 (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6344__B1 (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4633__A1 (.DIODE(_1307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6437__A2 (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6419__A2 (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6374__A2 (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4360__A (.DIODE(_1308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__A2 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6405__A2 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6399__A2 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6392__A2 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6385__A2 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6378__A2 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6364__A2 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6355__A2 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6341__A2 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4626__A2 (.DIODE(_1309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6438__A1 (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__A1 (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6375__A1 (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6354__A (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__A (.DIODE(_1311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__B (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__A1 (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__A (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__A (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__A (.DIODE(_1317_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__C (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__A2 (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4477__B (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__B (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4370__B (.DIODE(_1318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5274__S (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__A1 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__A1 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__A (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__A (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__B2 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4521__A (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__A2 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__B2 (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__A (.DIODE(_1319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__B (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__S (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4405__S (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__S (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4403__S (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4401__A (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__S (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__S (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4378__C1 (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4373__B (.DIODE(_1321_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__A1 (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__B1 (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4375__A (.DIODE(_1322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__A2 (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__C1 (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4375__B (.DIODE(_1323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4518__S (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4457__A (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4376__B (.DIODE(_1324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__B (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__A1 (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__A1 (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__A1 (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__C (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__A (.DIODE(_1326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__C (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__A2 (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__A2 (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__A2 (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4415__D (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4379__B (.DIODE(_1327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__S (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__S (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__A1 (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__A (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__S (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4539__A (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4380__B (.DIODE(_1328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__B1 (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__B1 (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__B1 (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__B1 (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__B1 (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__B1 (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__B1 (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__B1 (.DIODE(_1337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4394__B (.DIODE(_1338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__A2 (.DIODE(_1340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__A2 (.DIODE(_1340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__B1 (.DIODE(_1340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4514__A2 (.DIODE(_1340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__B1 (.DIODE(_1340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4435__A (.DIODE(_1340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4393__B1 (.DIODE(_1340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__A2 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__A2 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__C1 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__C1 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__A2 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__A2 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__C1 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__A2 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__C1 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4393__C1 (.DIODE(_1341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__B (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__A (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__B1 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__A1 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__A3 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__B1 (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__A (.DIODE(_1343_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__C (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5150__B (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4491__C1 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4490__A2 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4481__A4 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4479__B2 (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4397__B (.DIODE(_1345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__A3 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6167__A1 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6135__B2 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6133__A3 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__B2 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4445__A2 (.DIODE(_1346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__A2 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__A2 (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__A (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__A (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__A (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4648__A (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__A (.DIODE(_1347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__A (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4651__A (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4400__B (.DIODE(_1348_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__S (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4641__S (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4616__A1 (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__S (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4461__A1 (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__S (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4420__A1 (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4418__S (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4409__S (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__S (.DIODE(_1350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__B2 (.DIODE(_1351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__A2 (.DIODE(_1351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__A (.DIODE(_1351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__A (.DIODE(_1351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__A (.DIODE(_1351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__A1 (.DIODE(_1351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__A_N (.DIODE(_1351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__A (.DIODE(_1351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__B (.DIODE(_1351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__B (.DIODE(_1351_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6112__A1 (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__A2 (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__A (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__A (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4643__A (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__A (.DIODE(_1352_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__A2 (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__A (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__A1 (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__B (.DIODE(_1353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__B2 (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__A2 (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5013__A1 (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5012__A1 (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__A (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__A (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4676__A_N (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4647__B_N (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__C (.DIODE(_1354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__A2 (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__A2 (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__A (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__A (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__A (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__A1 (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4673__B (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4672__A_N (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4407__D (.DIODE(_1355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__A (.DIODE(_1358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__A (.DIODE(_1358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__A (.DIODE(_1358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__A (.DIODE(_1358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__B (.DIODE(_1358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__B (.DIODE(_1358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4410__D_N (.DIODE(_1358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__A_N (.DIODE(_1359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__B (.DIODE(_1359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4442__A_N (.DIODE(_1359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__B2 (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5148__B1 (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__A (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__A1 (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4908__A1 (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4907__A1 (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4668__B (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4655__B (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4468__B1 (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4426__A2 (.DIODE(_1363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__A (.DIODE(_1366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__A (.DIODE(_1366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__A1 (.DIODE(_1366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4665__B (.DIODE(_1366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4659__B (.DIODE(_1366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4555__A (.DIODE(_1366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__A2 (.DIODE(_1366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__A (.DIODE(_1367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__B (.DIODE(_1367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4469__A (.DIODE(_1367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4421__A3 (.DIODE(_1367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6114__A1 (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__A2 (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5029__A1 (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__A (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__A (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4637__A (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__A (.DIODE(_1371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__B (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__A2 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__A (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__A (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A1 (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4681__B (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4639__A (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4425__B (.DIODE(_1373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__A2 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__A2 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__A2 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4594__B1 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__A1 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__B1 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__A2 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__B1 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__A2 (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4428__A (.DIODE(_1376_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__A2 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__A2 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__A2 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__A2 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__A2 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__A2 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__A2 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__B1 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__A2 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__A2 (.DIODE(_1377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4550__A2 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__B1 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4526__A2 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__A2 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4439__A2 (.DIODE(_1378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__A2 (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__A2 (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__A2 (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__A2 (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__A2 (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__A2 (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__A2 (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__A2 (.DIODE(_1379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__B1 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4584__B1 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__A2 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4546__B1 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__B1 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4531__B1 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__B1 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4512__B1 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__B1 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4432__B1 (.DIODE(_1380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__A2 (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__A2 (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__A2 (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__A2 (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__A2 (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__A2 (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__A2 (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__A2 (.DIODE(_1382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4587__B1 (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__B1 (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__A2 (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__B1 (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__B1 (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__B1 (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__B1 (.DIODE(_1383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__A2 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__A2 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__B1 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__B1 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__A2 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__B1 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__A2 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__B1 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__B1 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__A2 (.DIODE(_1384_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__B1 (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__B1 (.DIODE(_1388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__A2 (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__A (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__A0 (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5065__B (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4951__B (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__A2 (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__B (.DIODE(_1389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4453__A (.DIODE(_1395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__A2 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__A2 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__A2 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4583__C (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__A2 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__A2 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__A2 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4530__C (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4510__A (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__A2 (.DIODE(_1400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__A1 (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4983__A1 (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__A0 (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4615__A2 (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__B (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__B (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4485__A1 (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4484__B1 (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4455__A (.DIODE(_1403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6166__A0 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__A1 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__B1 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4456__A2 (.DIODE(_1404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5611__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5546__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5485__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__S (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4458__A (.DIODE(_1406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6127__B (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5216__S (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__B (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__S (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4942__S (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4939__S (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4923__S (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4911__S (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__B (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4459__S (.DIODE(_1407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6120__A2 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A2 (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__A (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__A (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__A (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4467__A (.DIODE(_1410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__A (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__B (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4464__A (.DIODE(_1412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A1 (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5279__A (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__A (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__A2 (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__A (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__A (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4556__A (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4554__S (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4475__A (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4465__B (.DIODE(_1413_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__A1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__A1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__A1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4906__A2 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__A1 (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__C (.DIODE(_1414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__C (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__B (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__B (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5311__B (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5273__B (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__C1 (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__C1 (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__A (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4924__A (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4470__B (.DIODE(_1418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4606__A (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4537__A (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4487__A (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4486__A (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4483__B1 (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4482__A (.DIODE(_1427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__A2 (.DIODE(_1445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__A1 (.DIODE(_1445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__B1 (.DIODE(_1445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__B1 (.DIODE(_1445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__B1 (.DIODE(_1445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__A1 (.DIODE(_1445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__B1 (.DIODE(_1445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__A1 (.DIODE(_1445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__B (.DIODE(_1445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__B (.DIODE(_1445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__B1 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__B1 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__B1 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__B1 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__B2 (.DIODE(_1446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6117__B1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__A (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__B1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__B1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5320__A (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A2 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5281__A1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__C1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5179__A1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4620__A1 (.DIODE(_1451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5008__B (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4508__A (.DIODE(_1456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__A0 (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__A0 (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__B2 (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__A2 (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__B (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__A2 (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5009__B (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4938__A2 (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__A0 (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4509__A (.DIODE(_1457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A2 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__A2 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5103__A2 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5097__A2 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A2 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5092__A2 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__A2 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__B (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4904__A2 (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4511__C (.DIODE(_1459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__A3 (.DIODE(_1464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__A1 (.DIODE(_1465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6228__B2 (.DIODE(_1465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6217__A0 (.DIODE(_1465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__B2 (.DIODE(_1465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4995__B (.DIODE(_1465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4994__B (.DIODE(_1465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4937__A2 (.DIODE(_1465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__A1 (.DIODE(_1465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4517__A (.DIODE(_1465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6120__B2 (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__A (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__A (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4520__A (.DIODE(_1468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__B1 (.DIODE(_1472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4609__B (.DIODE(_1472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__B1 (.DIODE(_1472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__B1 (.DIODE(_1472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4579__B1 (.DIODE(_1472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__B1 (.DIODE(_1472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__B1 (.DIODE(_1472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__C (.DIODE(_1472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6267__A0 (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__B1 (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__A2 (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__B2 (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4964__B (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4941__A2 (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__A0 (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4529__A (.DIODE(_1477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__A0 (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5027__B (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__B (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4962__A2 (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__A0 (.DIODE(_1478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__B1 (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__B1 (.DIODE(_1480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__B2 (.DIODE(_1483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__B2 (.DIODE(_1483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5162__A1 (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__B (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5024__A (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__B (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4966__A2 (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4536__A1 (.DIODE(_1484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5424__S (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5345__S (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5309__S (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5269__S (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5164__S (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4928__A (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4920__S (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4915__S (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__B (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4553__A1 (.DIODE(_1488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__B2 (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6267__A1 (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__B2 (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5028__A (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4960__B (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4959__B (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4957__A2 (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4933__A2 (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__B2 (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4545__A (.DIODE(_1493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__B1 (.DIODE(_1499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__B1 (.DIODE(_1499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__B1 (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5165__A1 (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5033__B (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4953__A2 (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4552__A1 (.DIODE(_1500_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5465__A1 (.DIODE(_1504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__B2 (.DIODE(_1504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5384__A (.DIODE(_1504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5322__A1 (.DIODE(_1504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__C1 (.DIODE(_1504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5228__A1 (.DIODE(_1504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5178__A1 (.DIODE(_1504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4946__A (.DIODE(_1504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4718__B (.DIODE(_1504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4619__A1 (.DIODE(_1504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6118__A1 (.DIODE(_1505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5551__A1 (.DIODE(_1505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5387__A1 (.DIODE(_1505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5358__A1 (.DIODE(_1505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5357__A (.DIODE(_1505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5319__A (.DIODE(_1505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5226__A1 (.DIODE(_1505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5221__A1 (.DIODE(_1505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5167__S (.DIODE(_1505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__A (.DIODE(_1505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5280__A2 (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5278__A (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5275__B (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5272__B (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5224__B1 (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5223__A (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__A2 (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5219__B (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5218__B (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4558__B (.DIODE(_1506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5109__B1 (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4565__B (.DIODE(_1513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5391__B2 (.DIODE(_1515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4976__B (.DIODE(_1515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__A2 (.DIODE(_1515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__B (.DIODE(_1515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__A0 (.DIODE(_1515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__A0 (.DIODE(_1515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__A1 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__B2 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5355__A2 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5053__B (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5051__B (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4978__B (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4977__A2 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4967__B (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4914__A2 (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4574__A (.DIODE(_1522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__A0 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__A0 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A2 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__A0 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__A1 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4575__A1 (.DIODE(_1523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4581__A2 (.DIODE(_1526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__B1 (.DIODE(_1528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__B1 (.DIODE(_1528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5046__B (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5037__B (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__B (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4972__B (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4582__A (.DIODE(_1530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__A3 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__B2 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__A1 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__B (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5432__B2 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__A1 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__A2 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4909__A2 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__A3 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4590__A2 (.DIODE(_1531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__B1 (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__B1 (.DIODE(_1533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__B2 (.DIODE(_1536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__B2 (.DIODE(_1536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5161__A1 (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4998__B (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4997__A2 (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4589__B (.DIODE(_1537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__B1 (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__B1 (.DIODE(_1543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__B1 (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4597__B (.DIODE(_1545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6193__A1 (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__A1 (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5168__A1 (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__B (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4969__B (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4968__B (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__A2 (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__A0 (.DIODE(_1547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__B1 (.DIODE(_1552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__A2 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__A3 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__A2 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4990__B (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4986__B (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4985__B (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4918__A (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4816__A3 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4605__A1 (.DIODE(_1553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__A (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A1 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5277__S (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5276__S (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5222__S (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5220__A1 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A1 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__A1 (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5173__A (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__A (.DIODE(_1555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__B2 (.DIODE(_1561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__A3 (.DIODE(_1562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__A2 (.DIODE(_1562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5231__B (.DIODE(_1562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5043__B (.DIODE(_1562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5042__B (.DIODE(_1562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4984__B (.DIODE(_1562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4982__B (.DIODE(_1562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4921__A (.DIODE(_1562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__A1 (.DIODE(_1562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4614__C (.DIODE(_1562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5039__A (.DIODE(_1565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4657__B (.DIODE(_1565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4656__B (.DIODE(_1565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4617__B1 (.DIODE(_1565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5457__B (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5392__A1 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5359__B1 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5321__C1 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5288__A1 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5227__A (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5177__B1 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4618__B1 (.DIODE(_1566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4621__C1 (.DIODE(_1569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6482__A (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6458__A (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4623__A2 (.DIODE(_1570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__A1 (.DIODE(_1573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__A (.DIODE(_1573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4625__B (.DIODE(_1573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__B1 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6441__B1 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6416__B1 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6396__B1 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6352__D1 (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6349__A (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4632__C (.DIODE(_1580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5035__A (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4957__A1 (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4781__B (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4684__B (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4638__B (.DIODE(_1585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4963__A (.DIODE(_1587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4683__A2 (.DIODE(_1587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__B (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5060__A (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5025__A1 (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5015__A (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4679__B (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4642__B (.DIODE(_1589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5018__A (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5017__A1 (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4645__B (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4644__B (.DIODE(_1591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5004__A (.DIODE(_1596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5003__A1 (.DIODE(_1596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4650__B (.DIODE(_1596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4649__B (.DIODE(_1596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6119__A (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__A (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5390__A2 (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5389__A2 (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__A (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__A (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4974__A1 (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4973__A (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4653__B (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4652__A_N (.DIODE(_1599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__A2 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__A2 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__A2 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__A2 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__A2 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__A2 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__A2 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__A2 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__A2 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__A2 (.DIODE(_1640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__A2 (.DIODE(_1641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4797__B1 (.DIODE(_1641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__A2 (.DIODE(_1641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__A2 (.DIODE(_1641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__A2 (.DIODE(_1641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__A2 (.DIODE(_1641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__A2 (.DIODE(_1641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__A2 (.DIODE(_1641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__A2 (.DIODE(_1641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__A2 (.DIODE(_1641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4793__A (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4779__A (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4774__A (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4763__A (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4751__A (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4695__A (.DIODE(_1642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__B1 (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4786__B1 (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4768__B1 (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4757__B1 (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4743__A (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4737__B1 (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4730__B1 (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__B1 (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__B1 (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__B1 (.DIODE(_1643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4714__A2 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4703__A2 (.DIODE(_1646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__A2 (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4701__B (.DIODE(_1648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6330__A (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6327__A (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6324__A (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6321__A (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6307__A (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6304__A (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6301__A (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__S (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4744__A (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4706__A (.DIODE(_1653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6337__B1 (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6335__B1 (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6316__B1 (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6314__B1 (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6298__B1 (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4738__C1 (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4731__C1 (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4724__C1 (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__C1 (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__C1 (.DIODE(_1654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4721__B (.DIODE(_1659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4713__B (.DIODE(_1659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__C1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__C1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4787__C1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4780__C1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4775__C1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4769__C1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4764__C1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4758__C1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4752__C1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4745__C1 (.DIODE(_1687_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6475__B2 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6473__A (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6293__B2 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5682__A1 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5032__B (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__B (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4931__C (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4826__A0 (.DIODE(_1733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6255__A3 (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6253__B2 (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__A1 (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__B2 (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5014__B (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4940__A2 (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4802__A1 (.DIODE(_1734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__C1 (.DIODE(_1736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4804__A (.DIODE(_1736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6267__S (.DIODE(_1737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6241__S (.DIODE(_1737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__S (.DIODE(_1737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6166__S1 (.DIODE(_1737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__S0 (.DIODE(_1737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6108__A (.DIODE(_1737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__A1 (.DIODE(_1737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4834__A (.DIODE(_1737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4817__S (.DIODE(_1737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4805__A (.DIODE(_1737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6336__B (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__A2 (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6315__B (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__A2 (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6116__B (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4806__B1 (.DIODE(_1738_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6288__A1 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6287__B1 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__A2 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6220__A1 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6219__A (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6121__C1 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__C1 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4832__A (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__B2 (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__A (.DIODE(_1741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6286__A1 (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6165__B (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6120__A1 (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6117__A1 (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6113__A (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6111__A1 (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4831__A2 (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4811__B (.DIODE(_1743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6338__A1 (.DIODE(_1744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6317__A1 (.DIODE(_1744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6208__A2 (.DIODE(_1744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6133__A2 (.DIODE(_1744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__A1 (.DIODE(_1744_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__A1 (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5656__A2 (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4955__B (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4954__B (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4932__A2 (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4815__A2 (.DIODE(_1745_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6217__A1 (.DIODE(_1746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__B2 (.DIODE(_1746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__A2 (.DIODE(_1746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__A2 (.DIODE(_1746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5001__B (.DIODE(_1746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5000__B (.DIODE(_1746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4910__A2 (.DIODE(_1746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4814__A2 (.DIODE(_1746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6334__B (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__A2 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6313__B (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6300__A2 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4820__B1 (.DIODE(_1752_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6279__B (.DIODE(_1756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6278__B (.DIODE(_1756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4824__B1 (.DIODE(_1756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6106__S (.DIODE(_1760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4841__A2 (.DIODE(_1760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__A2 (.DIODE(_1760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4830__B (.DIODE(_1760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4829__B (.DIODE(_1760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6329__A1 (.DIODE(_1763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6326__A1 (.DIODE(_1763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6323__A1 (.DIODE(_1763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6320__A1 (.DIODE(_1763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6310__A (.DIODE(_1763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6306__A1 (.DIODE(_1763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6303__A1 (.DIODE(_1763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6300__A1 (.DIODE(_1763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4837__A1 (.DIODE(_1763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__A (.DIODE(_1763_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6320__A2 (.DIODE(_1765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6110__A (.DIODE(_1765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4835__B (.DIODE(_1765_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6299__A (.DIODE(_1769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6289__S (.DIODE(_1769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6269__S (.DIODE(_1769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6257__S (.DIODE(_1769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6246__A1 (.DIODE(_1769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6221__A1 (.DIODE(_1769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6207__C1 (.DIODE(_1769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6133__A1 (.DIODE(_1769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6123__A1 (.DIODE(_1769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4840__A (.DIODE(_1769_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6643__B1 (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__B (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6342__A (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__A2 (.DIODE(_1774_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6635__B1 (.DIODE(_1776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__C1 (.DIODE(_1776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__C1 (.DIODE(_1776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__C1 (.DIODE(_1776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__C1 (.DIODE(_1776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__C1 (.DIODE(_1776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__C1 (.DIODE(_1776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__C1 (.DIODE(_1776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__C1 (.DIODE(_1776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4850__C1 (.DIODE(_1776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6699__A (.DIODE(_1777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6507__A1 (.DIODE(_1777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6500__A1 (.DIODE(_1777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4893__B (.DIODE(_1777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__A2 (.DIODE(_1777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__A2 (.DIODE(_1777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__A2 (.DIODE(_1777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__A2 (.DIODE(_1777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__A2 (.DIODE(_1777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4852__A (.DIODE(_1777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__A2 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__A2 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__A2 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__A2 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__A2 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__A2 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__A2 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__A2 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__A2 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__A2 (.DIODE(_1778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5996__A (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5972__A (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5947__A (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5925__A (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5901__A (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5879__A (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5854__A (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5826__A (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5779__A (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4871__A (.DIODE(_1788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__C1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5769__C1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__C1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__C1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__C1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__C1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__C1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__C1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__C1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__C1 (.DIODE(_1789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__B1 (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A2 (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5100__B1 (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4894__A (.DIODE(_1796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5510__A2 (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__S (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__S (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__S (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__S (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__S (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__S (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__S (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5070__S (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__S (.DIODE(_1801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__A2 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__B1 (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__C (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5069__A (.DIODE(_1803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6115__A2 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__A2 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__A1 (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__A (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4950__A (.DIODE(_1804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6205__A0 (.DIODE(_1811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6194__A0 (.DIODE(_1811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__B2 (.DIODE(_1811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5420__B (.DIODE(_1811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5169__A0 (.DIODE(_1811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5055__B (.DIODE(_1811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5050__B (.DIODE(_1811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4913__A2 (.DIODE(_1811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__A1 (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6166__A3 (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__B2 (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5040__B (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4917__A2 (.DIODE(_1815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6166__A1 (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__A3 (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__A0 (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4970__A2 (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4919__A2 (.DIODE(_1817_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6166__A2 (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__A1 (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__B2 (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5172__A1 (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4922__A2 (.DIODE(_1820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__A2 (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6117__A2 (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5667__A1 (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5666__A (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5381__A2 (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5217__A2 (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__A (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__A2 (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4936__A1 (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4934__S (.DIODE(_1827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__B1 (.DIODE(_1870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4981__A1 (.DIODE(_1870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__A1 (.DIODE(_1887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5325__A2 (.DIODE(_1887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5324__A (.DIODE(_1887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__A (.DIODE(_1887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5396__A2 (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4993__B (.DIODE(_1891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5649__A3 (.DIODE(_1925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5608__C1 (.DIODE(_1925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5607__A2 (.DIODE(_1925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5596__A2 (.DIODE(_1925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5030__A3 (.DIODE(_1925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6468__A1 (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5090__A (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5083__A1 (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5082__B (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5078__B1_N (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5068__B (.DIODE(_1966_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5076__A2 (.DIODE(_1971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5074__B (.DIODE(_1971_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5080__A1 (.DIODE(_1977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5086__A1 (.DIODE(_1982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5094__A1 (.DIODE(_1989_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6453__B (.DIODE(_2013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__B (.DIODE(_2013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__A2 (.DIODE(_2013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__B1 (.DIODE(_2013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A2 (.DIODE(_2013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__A2 (.DIODE(_2013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5199__C (.DIODE(_2016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__B (.DIODE(_2016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5136__C (.DIODE(_2016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5130__B (.DIODE(_2016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__C (.DIODE(_2016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5409__A (.DIODE(_2021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5374__B1 (.DIODE(_2021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__B1 (.DIODE(_2021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__B1 (.DIODE(_2021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__A2 (.DIODE(_2021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5248__B1 (.DIODE(_2021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__A2 (.DIODE(_2021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__C1 (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5640__A (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5628__A (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5297__C1 (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__B1 (.DIODE(_2030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5681__A1 (.DIODE(_2039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5594__C1 (.DIODE(_2039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__A1 (.DIODE(_2039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__B2 (.DIODE(_2039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5344__A (.DIODE(_2039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5160__A1 (.DIODE(_2039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6155__A0 (.DIODE(_2041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6132__D (.DIODE(_2041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5174__B (.DIODE(_2041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__A (.DIODE(_2041_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5356__A1 (.DIODE(_2042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5289__A1 (.DIODE(_2042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5152__B (.DIODE(_2042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5527__A (.DIODE(_2046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5362__A1 (.DIODE(_2046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5314__B1 (.DIODE(_2046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__B2 (.DIODE(_2046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5234__A1_N (.DIODE(_2046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__B1 (.DIODE(_2046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5479__B1 (.DIODE(_2047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5284__A1 (.DIODE(_2047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5157__B2 (.DIODE(_2047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5225__A2 (.DIODE(_2063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5176__A2 (.DIODE(_2063_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5180__B (.DIODE(_2070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6482__B (.DIODE(_2071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6458__B (.DIODE(_2071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__B (.DIODE(_2071_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6341__B1 (.DIODE(_2076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__A1 (.DIODE(_2076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__A1 (.DIODE(_2076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__B1 (.DIODE(_2077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5307__B1 (.DIODE(_2077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5254__A (.DIODE(_2077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5194__A (.DIODE(_2077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5187__A (.DIODE(_2077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__B1 (.DIODE(_2078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__S (.DIODE(_2078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__S (.DIODE(_2078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__S (.DIODE(_2078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__S (.DIODE(_2078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__S (.DIODE(_2078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__S (.DIODE(_2078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__S (.DIODE(_2078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__S (.DIODE(_2078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5188__S (.DIODE(_2078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5540__S (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5472__S (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__S (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__S (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__S (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__S (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__S (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__S (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__S (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__S (.DIODE(_2081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__A1 (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__A1 (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5632__A (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__A1 (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__A1 (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__B1 (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__B1 (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A1 (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5209__A1 (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5208__B (.DIODE(_2084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5574__S (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5541__S (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5473__S (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__S (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__S (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__S (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__S (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__S (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__S (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__S (.DIODE(_2101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__B1 (.DIODE(_2103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5239__B1 (.DIODE(_2117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__A (.DIODE(_2128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6457__A (.DIODE(_2128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5240__B (.DIODE(_2128_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6352__A2 (.DIODE(_2131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__A1 (.DIODE(_2131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5255__A2 (.DIODE(_2131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5292__B1 (.DIODE(_2156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6480__B (.DIODE(_2177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6457__B (.DIODE(_2177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5290__B (.DIODE(_2177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__A2 (.DIODE(_2180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__A1 (.DIODE(_2180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5293__A1 (.DIODE(_2180_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5329__B1 (.DIODE(_2195_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__A (.DIODE(_2213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6460__A (.DIODE(_2213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5327__B (.DIODE(_2213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6365__A2 (.DIODE(_2216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__A1 (.DIODE(_2216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5330__B2 (.DIODE(_2216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__A (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__A (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5342__B (.DIODE(_2227_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5366__B1 (.DIODE(_2229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6484__B (.DIODE(_2249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6459__A (.DIODE(_2249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5365__A2 (.DIODE(_2249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6375__A2 (.DIODE(_2252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__A1 (.DIODE(_2252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5367__A1 (.DIODE(_2252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__A2 (.DIODE(_2256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__A2_N (.DIODE(_2256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__A2 (.DIODE(_2256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__A2 (.DIODE(_2256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5564__B (.DIODE(_2256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__A2 (.DIODE(_2256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__A2 (.DIODE(_2256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__A2 (.DIODE(_2256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A2 (.DIODE(_2256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__A2 (.DIODE(_2256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__A2 (.DIODE(_2257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__B1 (.DIODE(_2257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__B1 (.DIODE(_2257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__A2 (.DIODE(_2257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__A2 (.DIODE(_2257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__A2 (.DIODE(_2257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__A2 (.DIODE(_2257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__A2 (.DIODE(_2257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__A2 (.DIODE(_2257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A2 (.DIODE(_2257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5408__B_N (.DIODE(_2263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5379__B (.DIODE(_2263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__B1 (.DIODE(_2265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__B1 (.DIODE(_2277_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5395__B (.DIODE(_2278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5394__A1 (.DIODE(_2278_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5400__C1 (.DIODE(_2284_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6493__A (.DIODE(_2285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6456__A (.DIODE(_2285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5401__B (.DIODE(_2285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6379__A2 (.DIODE(_2288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5711__A1 (.DIODE(_2288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5404__A1 (.DIODE(_2288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6593__C (.DIODE(_2293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__B1 (.DIODE(_2293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__B1 (.DIODE(_2293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__B1 (.DIODE(_2293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__B1 (.DIODE(_2293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__B1 (.DIODE(_2293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__B1 (.DIODE(_2293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__B1 (.DIODE(_2293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__B1 (.DIODE(_2293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5412__B1 (.DIODE(_2293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6499__B (.DIODE(_2294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5689__B1 (.DIODE(_2294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5639__A2 (.DIODE(_2294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5627__A2 (.DIODE(_2294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5577__B1 (.DIODE(_2294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5566__B1 (.DIODE(_2294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5512__B1 (.DIODE(_2294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5502__B1 (.DIODE(_2294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5446__B1 (.DIODE(_2294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__A2 (.DIODE(_2294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5444__B_N (.DIODE(_2300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5417__B (.DIODE(_2300_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__B1 (.DIODE(_2302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5435__B1 (.DIODE(_2311_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__B1 (.DIODE(_2312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5431__B1 (.DIODE(_2312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6493__B (.DIODE(_2320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6461__B (.DIODE(_2320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5438__A2 (.DIODE(_2320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6386__A2 (.DIODE(_2323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__A1 (.DIODE(_2323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5440__A1 (.DIODE(_2323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5505__B_N (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5450__B (.DIODE(_2332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__B1 (.DIODE(_2334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5467__A (.DIODE(_2338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5680__B2 (.DIODE(_2340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5651__B (.DIODE(_2340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5618__A2 (.DIODE(_2340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5591__A2 (.DIODE(_2340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5554__B2 (.DIODE(_2340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5528__A2 (.DIODE(_2340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__B1 (.DIODE(_2340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5464__A2 (.DIODE(_2340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5678__C1 (.DIODE(_2341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5647__C1 (.DIODE(_2341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__C1 (.DIODE(_2341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__C1 (.DIODE(_2341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5552__C1 (.DIODE(_2341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5523__C1 (.DIODE(_2341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__C1 (.DIODE(_2341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__C1 (.DIODE(_2341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6488__A (.DIODE(_2350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__A (.DIODE(_2350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5468__B (.DIODE(_2350_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__A2 (.DIODE(_2353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__A1 (.DIODE(_2353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5471__A1 (.DIODE(_2353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5499__B1 (.DIODE(_2358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5495__B1 (.DIODE(_2371_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6488__B (.DIODE(_2378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6463__B (.DIODE(_2378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5497__B (.DIODE(_2378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__A2 (.DIODE(_2381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__A1 (.DIODE(_2381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__A2 (.DIODE(_2381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6399__B1 (.DIODE(_2382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5507__A2 (.DIODE(_2382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5506__A1 (.DIODE(_2382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5569__B_N (.DIODE(_2396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5516__B (.DIODE(_2396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5535__B1 (.DIODE(_2410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6486__A (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6462__A_N (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5537__A2 (.DIODE(_2416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6406__A2 (.DIODE(_2419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__A1 (.DIODE(_2419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5539__A1 (.DIODE(_2419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5562__B1 (.DIODE(_2423_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5555__A2 (.DIODE(_2430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6486__B (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6462__B (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5560__B (.DIODE(_2439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__A2 (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__A1 (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5572__A2 (.DIODE(_2442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6412__B1 (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5571__A2 (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5570__A1 (.DIODE(_2443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5625__B_N (.DIODE(_2459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5581__B (.DIODE(_2459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5595__C1 (.DIODE(_2473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__A (.DIODE(_2475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6455__A (.DIODE(_2475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5597__B (.DIODE(_2475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__A2 (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__A1 (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5600__A1 (.DIODE(_2478_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5708__S (.DIODE(_2481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5706__S (.DIODE(_2481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5704__S (.DIODE(_2481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5702__S (.DIODE(_2481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5700__S (.DIODE(_2481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5698__S (.DIODE(_2481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5696__S (.DIODE(_2481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5664__S (.DIODE(_2481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5635__S (.DIODE(_2481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5603__S (.DIODE(_2481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6487__B (.DIODE(_2499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6455__B (.DIODE(_2499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5622__B (.DIODE(_2499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__A2 (.DIODE(_2502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__A1 (.DIODE(_2502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5633__A2 (.DIODE(_2502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__B (.DIODE(_2508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5637__B (.DIODE(_2508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5631__B (.DIODE(_2508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5687__C (.DIODE(_2520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5644__B (.DIODE(_2520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__A (.DIODE(_2534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5658__B (.DIODE(_2534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6438__A2 (.DIODE(_2538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__A1 (.DIODE(_2538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5662__A1 (.DIODE(_2538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6492__B (.DIODE(_2558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6473__B (.DIODE(_2558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6471__A1 (.DIODE(_2558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6454__C1 (.DIODE(_2558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5684__A2 (.DIODE(_2558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__B2 (.DIODE(_2561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__A2 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__A1 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5694__A2 (.DIODE(_2562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5693__A2 (.DIODE(_2567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5692__B (.DIODE(_2567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__S (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__S (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5725__S (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5723__S (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5721__S (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5719__S (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5717__S (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5715__S (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5713__S (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5711__S (.DIODE(_2579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__S (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__S (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__S (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__S (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__S (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__S (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__S (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__S (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5734__S (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__S (.DIODE(_2590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6062__B (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6025__B (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__B (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__B (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__B (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__B (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5756__A (.DIODE(_2602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__B (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6024__B (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__B (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5949__B (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__B (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__B (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5873__B (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__B (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__B (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__B (.DIODE(_2603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__A1 (.DIODE(_2604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A1 (.DIODE(_2604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A1 (.DIODE(_2604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__A1 (.DIODE(_2604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A1 (.DIODE(_2604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__A1 (.DIODE(_2604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5769__A1 (.DIODE(_2604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__A1 (.DIODE(_2604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__A1 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__A1 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__A1 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A1 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__A1 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5877__A1 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__A1 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5764__A2 (.DIODE(_2607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5801__A (.DIODE(_2608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5799__B (.DIODE(_2608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5794__B (.DIODE(_2608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5789__B (.DIODE(_2608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5784__B (.DIODE(_2608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5762__A (.DIODE(_2608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__A (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__A (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__A (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__A (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__A (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__A (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__B (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5773__B (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__B (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5763__B (.DIODE(_2609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__A1 (.DIODE(_2613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__A1 (.DIODE(_2613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5992__A1 (.DIODE(_2613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__A1 (.DIODE(_2613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__A1 (.DIODE(_2613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__A1 (.DIODE(_2613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__A1 (.DIODE(_2613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5769__A2 (.DIODE(_2613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6070__A1 (.DIODE(_2617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__A1 (.DIODE(_2617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5994__A1 (.DIODE(_2617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__A1 (.DIODE(_2617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__A1 (.DIODE(_2617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__A1 (.DIODE(_2617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__A1 (.DIODE(_2617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5774__A2 (.DIODE(_2617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__A1 (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__A1 (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__A1 (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5959__A1 (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__A1 (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__A1 (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5846__A1 (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__A2 (.DIODE(_2621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__C1 (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5818__C1 (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5814__C1 (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__C1 (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5807__C1 (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__C1 (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__C1 (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__C1 (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__C1 (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5780__C1 (.DIODE(_2623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__A1 (.DIODE(_2626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__A1 (.DIODE(_2626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__A1 (.DIODE(_2626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__A1 (.DIODE(_2626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__A1 (.DIODE(_2626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__A1 (.DIODE(_2626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__A1 (.DIODE(_2626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5785__A2 (.DIODE(_2626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6076__A1 (.DIODE(_2630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__A1 (.DIODE(_2630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6001__A1 (.DIODE(_2630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5963__A1 (.DIODE(_2630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__A1 (.DIODE(_2630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__A1 (.DIODE(_2630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5850__A1 (.DIODE(_2630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5790__A2 (.DIODE(_2630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5965__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__A1 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5795__A2 (.DIODE(_2634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__A1 (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__A1 (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6005__A1 (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A1 (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__A1 (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5892__A1 (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__A1 (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5800__A2 (.DIODE(_2638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A2_N (.DIODE(_2642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__A2_N (.DIODE(_2642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5824__A2_N (.DIODE(_2642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5820__A2_N (.DIODE(_2642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5816__A2_N (.DIODE(_2642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5812__A2_N (.DIODE(_2642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__A2_N (.DIODE(_2642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__A2_N (.DIODE(_2642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6082__A (.DIODE(_2644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__A (.DIODE(_2644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6007__A (.DIODE(_2644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__A (.DIODE(_2644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__A (.DIODE(_2644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5894__A (.DIODE(_2644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5857__A (.DIODE(_2644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5806__B (.DIODE(_2644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6084__A (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__A (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6009__A (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__A (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__A (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5896__A (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5859__A (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5809__B (.DIODE(_2646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__A (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__A (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6011__A (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__A (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__A (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__A (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5861__A (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5813__B (.DIODE(_2649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__A (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6051__A (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__A (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__A (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__A (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__A (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5863__A (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5817__B (.DIODE(_2652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6091__A (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__A (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__A (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__A (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__A (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__A (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5865__A (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5821__B (.DIODE(_2655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__A (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__A (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6017__A (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5980__A (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__A (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__A (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5867__A (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5825__B (.DIODE(_2658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5852__C1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5850__C1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5848__C1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5846__C1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5844__C1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5842__C1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5840__C1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5835__C1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5831__C1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5827__C1 (.DIODE(_2660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6095__A (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__A (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__A (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5982__A (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__A (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__A (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5869__A (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5830__B (.DIODE(_2662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__A (.DIODE(_2665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__A (.DIODE(_2665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__A (.DIODE(_2665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__A (.DIODE(_2665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__A (.DIODE(_2665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__A (.DIODE(_2665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5871__A (.DIODE(_2665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5834__B (.DIODE(_2665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5877__C1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__C1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__C1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__C1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__C1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__C1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__C1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__C1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__C1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5855__C1 (.DIODE(_2678_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5909__B (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5907__B (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5905__B (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5903__B (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5900__B (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5898__B (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5883__B (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5881__B (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__B (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__B (.DIODE(_2690_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__C1 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5897__C1 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5895__C1 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5892__C1 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5890__C1 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5888__C1 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5886__C1 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5884__C1 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5882__C1 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5880__C1 (.DIODE(_2693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5923__C1 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5921__C1 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5919__C1 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5917__C1 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5915__C1 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5910__C1 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5908__C1 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__C1 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5904__C1 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5902__C1 (.DIODE(_2705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5946__B (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5944__B (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5942__B (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5940__B (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5938__B (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5936__B (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__B (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__B (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__B (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__B (.DIODE(_2712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5943__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5930__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5928__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5926__C1 (.DIODE(_2719_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__A2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__A2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5943__A2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__A2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5939__A2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__A2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5934__B (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5933__A2 (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5932__B (.DIODE(_2722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__C1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__C1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5965__C1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5963__C1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__C1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5959__C1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__C1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__C1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__C1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__C1 (.DIODE(_2731_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5967__A2 (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5965__A2 (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5963__A2 (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5961__A2 (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5959__A2 (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5957__A2 (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5955__A2 (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5953__A2 (.DIODE(_2732_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5968__A (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5966__B (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5964__B (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5962__B (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5960__B (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5951__A (.DIODE(_2733_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5984__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5982__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5980__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5978__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5976__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5974__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5958__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5956__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5954__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5952__B (.DIODE(_2734_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5985__A2 (.DIODE(_2743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5983__A2 (.DIODE(_2743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__A2 (.DIODE(_2743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__A2 (.DIODE(_2743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__A2 (.DIODE(_2743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__A2 (.DIODE(_2743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__A2 (.DIODE(_2743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5971__B (.DIODE(_2743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5970__A2 (.DIODE(_2743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5969__B (.DIODE(_2743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5994__C1 (.DIODE(_2746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5992__C1 (.DIODE(_2746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5990__C1 (.DIODE(_2746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5985__C1 (.DIODE(_2746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5983__C1 (.DIODE(_2746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__C1 (.DIODE(_2746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__C1 (.DIODE(_2746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__C1 (.DIODE(_2746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__C1 (.DIODE(_2746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__C1 (.DIODE(_2746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6022__B (.DIODE(_2755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6020__B (.DIODE(_2755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6017__B (.DIODE(_2755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6015__B (.DIODE(_2755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6013__B (.DIODE(_2755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6011__B (.DIODE(_2755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5995__B (.DIODE(_2755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5993__B (.DIODE(_2755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5991__B (.DIODE(_2755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5989__B (.DIODE(_2755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__C1 (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6014__C1 (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__C1 (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6010__C1 (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6008__C1 (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6005__C1 (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6003__C1 (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6001__C1 (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5999__C1 (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__5997__C1 (.DIODE(_2760_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6040__C1 (.DIODE(_2772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6038__C1 (.DIODE(_2772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6036__C1 (.DIODE(_2772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6034__C1 (.DIODE(_2772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6032__C1 (.DIODE(_2772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6030__C1 (.DIODE(_2772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6028__C1 (.DIODE(_2772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6023__C1 (.DIODE(_2772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6021__C1 (.DIODE(_2772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6019__C1 (.DIODE(_2772_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6044__A (.DIODE(_2776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__B (.DIODE(_2776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6039__B (.DIODE(_2776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6037__B (.DIODE(_2776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6035__B (.DIODE(_2776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6026__A (.DIODE(_2776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6059__B (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6057__B (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6055__B (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6053__B (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6051__B (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6049__B (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6033__B (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__B (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6029__B (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6027__B (.DIODE(_2777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6065__C1 (.DIODE(_2786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6060__C1 (.DIODE(_2786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6058__C1 (.DIODE(_2786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6056__C1 (.DIODE(_2786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6054__C1 (.DIODE(_2786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6052__C1 (.DIODE(_2786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__C1 (.DIODE(_2786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6048__C1 (.DIODE(_2786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6046__C1 (.DIODE(_2786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6043__C1 (.DIODE(_2786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6060__A2 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6058__A2 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6056__A2 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6054__A2 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6052__A2 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6050__A2 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6048__A2 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6047__B (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6046__A2 (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6045__B (.DIODE(_2787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6097__B (.DIODE(_2798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6095__B (.DIODE(_2798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6093__B (.DIODE(_2798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6091__B (.DIODE(_2798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6088__B (.DIODE(_2798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6086__B (.DIODE(_2798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6071__B (.DIODE(_2798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__B (.DIODE(_2798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6066__B (.DIODE(_2798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__B (.DIODE(_2798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6085__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6080__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6078__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6076__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6074__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6072__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6070__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6068__C1 (.DIODE(_2801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6510__C1 (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6478__C1 (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6472__C1 (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6469__C1 (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6466__C1 (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__C1 (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6096__C1 (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__C1 (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__C1 (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__C1 (.DIODE(_2813_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6448__A (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6442__A (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6435__A (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6423__A (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6417__A (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6410__A (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6403__A (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6397__A (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6345__A (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6102__B (.DIODE(_2819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6281__B1 (.DIODE(_2822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6172__B1 (.DIODE(_2822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6163__A1 (.DIODE(_2822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6160__B1 (.DIODE(_2822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6105__B1 (.DIODE(_2822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6124__B (.DIODE(_2840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6293__A2 (.DIODE(_2843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__B1 (.DIODE(_2843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__A2 (.DIODE(_2843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6228__A2 (.DIODE(_2843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__A2 (.DIODE(_2843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__C1 (.DIODE(_2843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__C1 (.DIODE(_2843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6144__A (.DIODE(_2843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__B1 (.DIODE(_2843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6135__A2 (.DIODE(_2843_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6284__A2 (.DIODE(_2844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6263__B2 (.DIODE(_2844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6203__B1 (.DIODE(_2844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6174__A2 (.DIODE(_2844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6151__A2 (.DIODE(_2844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6128__A (.DIODE(_2844_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6293__B1 (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__B1 (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6253__B1 (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6239__B1 (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6228__B1 (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6215__B1 (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6190__B1 (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6183__B1 (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6143__A2 (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6135__B1 (.DIODE(_2845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6275__A (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6252__B (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6240__A1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6229__A1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6216__A1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6204__A1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6191__A1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6184__A1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6142__A1 (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6134__A (.DIODE(_2846_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__A1 (.DIODE(_2852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__A1 (.DIODE(_2852_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6176__A2 (.DIODE(_2853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6138__A2 (.DIODE(_2853_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__B (.DIODE(_2973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__B (.DIODE(_2973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6290__B (.DIODE(_2991_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__A3 (.DIODE(_3026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6429__A (.DIODE(_3026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6360__B (.DIODE(_3026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__B (.DIODE(_3026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__B1 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__B1 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__B1 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6632__B1 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6390__A (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6383__A (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6376__A (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6369__A (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6362__A (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6346__C1 (.DIODE(_3029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6447__A1 (.DIODE(_3036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6434__A1 (.DIODE(_3036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__A1 (.DIODE(_3036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6406__A1 (.DIODE(_3036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__A1 (.DIODE(_3036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__A1 (.DIODE(_3036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6386__A1 (.DIODE(_3036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6379__A1 (.DIODE(_3036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6365__A1 (.DIODE(_3036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__A1 (.DIODE(_3036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6438__C1 (.DIODE(_3038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6420__C1 (.DIODE(_3038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6413__C1 (.DIODE(_3038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6406__C1 (.DIODE(_3038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6400__C1 (.DIODE(_3038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6393__C1 (.DIODE(_3038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6386__C1 (.DIODE(_3038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6379__C1 (.DIODE(_3038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6365__C1 (.DIODE(_3038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6357__C1 (.DIODE(_3038_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6408__D (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6407__A3 (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6395__B (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6394__B (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6389__A2 (.DIODE(_3066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6497__A1 (.DIODE(_3119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6496__B (.DIODE(_3119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6474__B1 (.DIODE(_3119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6458__D (.DIODE(_3119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6451__A2 (.DIODE(_3119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6573__A2 (.DIODE(_3164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6569__A2 (.DIODE(_3164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6565__A2 (.DIODE(_3164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6561__A2 (.DIODE(_3164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6557__A2 (.DIODE(_3164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6552__A2 (.DIODE(_3164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6501__A (.DIODE(_3164_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6548__A2 (.DIODE(_3165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6544__A2 (.DIODE(_3165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6540__A2 (.DIODE(_3165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6536__A2 (.DIODE(_3165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__A2 (.DIODE(_3165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6528__A2 (.DIODE(_3165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6523__A2 (.DIODE(_3165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6519__A2 (.DIODE(_3165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__A2 (.DIODE(_3165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6510__A2 (.DIODE(_3165_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6547__A1 (.DIODE(_3166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6543__A1 (.DIODE(_3166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6539__A1 (.DIODE(_3166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6535__A1 (.DIODE(_3166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6531__A1 (.DIODE(_3166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__A1 (.DIODE(_3166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6522__A1 (.DIODE(_3166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6518__A1 (.DIODE(_3166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__A1 (.DIODE(_3166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6509__A1 (.DIODE(_3166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__A1 (.DIODE(_3167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6541__S (.DIODE(_3167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6537__S (.DIODE(_3167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__S (.DIODE(_3167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6529__S (.DIODE(_3167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6524__S (.DIODE(_3167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__S (.DIODE(_3167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6516__S (.DIODE(_3167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6511__S (.DIODE(_3167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6504__S (.DIODE(_3167_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__A1 (.DIODE(_3169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__A1 (.DIODE(_3169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__A1 (.DIODE(_3169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6560__A1 (.DIODE(_3169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6555__A1 (.DIODE(_3169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6551__A1 (.DIODE(_3169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6521__B (.DIODE(_3169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6517__B (.DIODE(_3169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6512__B (.DIODE(_3169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6506__B (.DIODE(_3169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6572__C1 (.DIODE(_3171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6568__C1 (.DIODE(_3171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6564__C1 (.DIODE(_3171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6560__C1 (.DIODE(_3171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6555__C1 (.DIODE(_3171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6551__C1 (.DIODE(_3171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6508__A (.DIODE(_3171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6547__C1 (.DIODE(_3172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6543__C1 (.DIODE(_3172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6539__C1 (.DIODE(_3172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6535__C1 (.DIODE(_3172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6531__C1 (.DIODE(_3172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6527__C1 (.DIODE(_3172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6522__C1 (.DIODE(_3172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6518__C1 (.DIODE(_3172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6513__C1 (.DIODE(_3172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6509__C1 (.DIODE(_3172_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6552__C1 (.DIODE(_3177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6548__C1 (.DIODE(_3177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6544__C1 (.DIODE(_3177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6540__C1 (.DIODE(_3177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6536__C1 (.DIODE(_3177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__C1 (.DIODE(_3177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6528__C1 (.DIODE(_3177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6523__C1 (.DIODE(_3177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6519__C1 (.DIODE(_3177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6515__C1 (.DIODE(_3177_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6563__B (.DIODE(_3185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6559__B (.DIODE(_3185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6554__B (.DIODE(_3185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6550__B (.DIODE(_3185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6546__B (.DIODE(_3185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6542__B (.DIODE(_3185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6538__B (.DIODE(_3185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6534__B (.DIODE(_3185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6530__B (.DIODE(_3185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6526__B (.DIODE(_3185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6543__A2 (.DIODE(_3197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__C1 (.DIODE(_3209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__C1 (.DIODE(_3209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__C1 (.DIODE(_3209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__C1 (.DIODE(_3209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6651__C1 (.DIODE(_3209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6573__C1 (.DIODE(_3209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6569__C1 (.DIODE(_3209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6565__C1 (.DIODE(_3209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6561__C1 (.DIODE(_3209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6557__C1 (.DIODE(_3209_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6629__A2 (.DIODE(_3236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6627__A2 (.DIODE(_3236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6606__A (.DIODE(_3236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6596__A (.DIODE(_3236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6595__A (.DIODE(_3236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6618__A2 (.DIODE(_3237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6616__A2 (.DIODE(_3237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6614__A2 (.DIODE(_3237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6612__A2 (.DIODE(_3237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6610__A2 (.DIODE(_3237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6608__A2 (.DIODE(_3237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6605__A2 (.DIODE(_3237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6603__A2 (.DIODE(_3237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6601__A2 (.DIODE(_3237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6599__A2 (.DIODE(_3237_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6630__A2 (.DIODE(_3238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6628__A2 (.DIODE(_3238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6626__A2 (.DIODE(_3238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6624__A2 (.DIODE(_3238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6622__A2 (.DIODE(_3238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6620__A2 (.DIODE(_3238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__A2 (.DIODE(_3238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6602__A2 (.DIODE(_3238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6600__A2 (.DIODE(_3238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6598__A2 (.DIODE(_3238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6690__C1 (.DIODE(_3239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6615__B1 (.DIODE(_3239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6613__B1 (.DIODE(_3239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__B1 (.DIODE(_3239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__B1 (.DIODE(_3239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__B1 (.DIODE(_3239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6604__B1 (.DIODE(_3239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6602__B1 (.DIODE(_3239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6600__B1 (.DIODE(_3239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6598__B1 (.DIODE(_3239_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6625__A2 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6623__A2 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6621__A2 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6619__A2 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6617__A2 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6615__A2 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6613__A2 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6611__A2 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6609__A2 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6607__A2 (.DIODE(_3244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__C1 (.DIODE(_3257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__C1 (.DIODE(_3257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__C1 (.DIODE(_3257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__C1 (.DIODE(_3257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__C1 (.DIODE(_3257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__C1 (.DIODE(_3257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__A3 (.DIODE(_3257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6637__A2 (.DIODE(_3257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6636__A2 (.DIODE(_3257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6632__A3 (.DIODE(_3257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6693__A2 (.DIODE(_3262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6692__A (.DIODE(_3262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__A2 (.DIODE(_3262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__B1 (.DIODE(_3262_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__B1 (.DIODE(_3264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6689__C1 (.DIODE(_3264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__A2 (.DIODE(_3264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6675__C1 (.DIODE(_3264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__A2 (.DIODE(_3264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6663__C1 (.DIODE(_3264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__A2 (.DIODE(_3264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6657__A (.DIODE(_3264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6651__A2 (.DIODE(_3264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6644__A (.DIODE(_3264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6724__B1 (.DIODE(_3312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6722__A2 (.DIODE(_3312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__A2 (.DIODE(_3312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6716__A2 (.DIODE(_3312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__A2 (.DIODE(_3312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6710__A2 (.DIODE(_3312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__A2 (.DIODE(_3312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6704__A2 (.DIODE(_3312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__6701__A (.DIODE(_3312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__4065__A0 (.DIODE(\core_1.de_jmp_pred ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3934__S (.DIODE(\core_1.de_jmp_pred ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5748__A1 (.DIODE(\core_1.dec_mem_access ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5509__A1 (.DIODE(\core_1.dec_mem_access ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5508__C1 (.DIODE(\core_1.dec_mem_access ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5189__A (.DIODE(\core_1.dec_mem_access ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4067__A0 (.DIODE(\core_1.dec_mem_access ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4902__A1 (.DIODE(\core_1.dec_mem_we ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4069__A0 (.DIODE(\core_1.dec_mem_we ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4371__A (.DIODE(\core_1.dec_r_bus_imm ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4369__C1 (.DIODE(\core_1.dec_r_bus_imm ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__B (.DIODE(\core_1.dec_r_bus_imm ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3992__A (.DIODE(\core_1.dec_r_bus_imm ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5205__A1 (.DIODE(\core_1.dec_sreg_irt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4361__B (.DIODE(\core_1.dec_sreg_irt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4083__A (.DIODE(\core_1.dec_sreg_irt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3910__A (.DIODE(\core_1.dec_sreg_irt ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6698__A2 (.DIODE(\core_1.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__B2 (.DIODE(\core_1.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__B2 (.DIODE(\core_1.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5243__A (.DIODE(\core_1.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5206__D1 (.DIODE(\core_1.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5203__D1 (.DIODE(\core_1.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5186__B (.DIODE(\core_1.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5147__A (.DIODE(\core_1.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5140__C1 (.DIODE(\core_1.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4079__A (.DIODE(\core_1.dec_sreg_jal_over ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6696__A (.DIODE(\core_1.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6639__A (.DIODE(\core_1.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6450__A (.DIODE(\core_1.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6350__B (.DIODE(\core_1.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4359__B (.DIODE(\core_1.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__A2 (.DIODE(\core_1.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3951__A (.DIODE(\core_1.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__B (.DIODE(\core_1.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3912__A1 (.DIODE(\core_1.dec_sreg_store ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4897__A (.DIODE(\core_1.dec_sys ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4087__A1 (.DIODE(\core_1.dec_sys ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4828__A (.DIODE(\core_1.decode.i_flush ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4160__A (.DIODE(\core_1.decode.i_flush ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3896__A (.DIODE(\core_1.decode.i_flush ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3891__A (.DIODE(\core_1.decode.i_flush ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3775__B (.DIODE(\core_1.decode.i_flush ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3724__B (.DIODE(\core_1.decode.i_flush ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__A (.DIODE(\core_1.decode.i_flush ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3522__A (.DIODE(\core_1.decode.i_flush ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4269__A1 (.DIODE(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4021__A1 (.DIODE(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4017__A1 (.DIODE(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4013__A (.DIODE(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3998__A1 (.DIODE(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3720__A1 (.DIODE(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3676__A1 (.DIODE(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__B (.DIODE(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__B (.DIODE(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3623__A (.DIODE(\core_1.decode.i_instr_l[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4290__A1 (.DIODE(\core_1.decode.i_instr_l[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4063__B2 (.DIODE(\core_1.decode.i_instr_l[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__B2 (.DIODE(\core_1.decode.i_instr_l[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__A1 (.DIODE(\core_1.decode.i_instr_l[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4293__A1 (.DIODE(\core_1.decode.i_instr_l[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__B2 (.DIODE(\core_1.decode.i_instr_l[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__A1 (.DIODE(\core_1.decode.i_instr_l[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4296__A1 (.DIODE(\core_1.decode.i_instr_l[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__B2 (.DIODE(\core_1.decode.i_instr_l[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__A1 (.DIODE(\core_1.decode.i_instr_l[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4299__A1 (.DIODE(\core_1.decode.i_instr_l[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4053__A1 (.DIODE(\core_1.decode.i_instr_l[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4022__B2 (.DIODE(\core_1.decode.i_instr_l[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4302__A1 (.DIODE(\core_1.decode.i_instr_l[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4055__A1 (.DIODE(\core_1.decode.i_instr_l[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4024__B2 (.DIODE(\core_1.decode.i_instr_l[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4305__A1 (.DIODE(\core_1.decode.i_instr_l[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4057__A1 (.DIODE(\core_1.decode.i_instr_l[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4026__B2 (.DIODE(\core_1.decode.i_instr_l[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4271__A1 (.DIODE(\core_1.decode.i_instr_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4088__A1 (.DIODE(\core_1.decode.i_instr_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3688__A (.DIODE(\core_1.decode.i_instr_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3672__A (.DIODE(\core_1.decode.i_instr_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3638__A (.DIODE(\core_1.decode.i_instr_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3629__A (.DIODE(\core_1.decode.i_instr_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3626__A (.DIODE(\core_1.decode.i_instr_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3624__A (.DIODE(\core_1.decode.i_instr_l[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4283__A1 (.DIODE(\core_1.decode.i_instr_l[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4060__B2 (.DIODE(\core_1.decode.i_instr_l[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__A2 (.DIODE(\core_1.decode.i_instr_l[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4045__A2 (.DIODE(\core_1.decode.i_instr_l[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4043__A (.DIODE(\core_1.decode.i_instr_l[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__A2 (.DIODE(\core_1.decode.i_instr_l[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4039__A2 (.DIODE(\core_1.decode.i_instr_l[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4036__A_N (.DIODE(\core_1.decode.i_instr_l[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4285__A1 (.DIODE(\core_1.decode.i_instr_l[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4061__B2 (.DIODE(\core_1.decode.i_instr_l[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4047__A1 (.DIODE(\core_1.decode.i_instr_l[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4044__A1_N (.DIODE(\core_1.decode.i_instr_l[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4041__A1 (.DIODE(\core_1.decode.i_instr_l[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4040__B2 (.DIODE(\core_1.decode.i_instr_l[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4037__A (.DIODE(\core_1.decode.i_instr_l[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4287__A1 (.DIODE(\core_1.decode.i_instr_l[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4062__B2 (.DIODE(\core_1.decode.i_instr_l[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4042__A (.DIODE(\core_1.decode.i_instr_l[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4035__A_N (.DIODE(\core_1.decode.i_instr_l[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6309__A (.DIODE(\core_1.decode.o_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6292__C1 (.DIODE(\core_1.decode.o_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6129__A (.DIODE(\core_1.decode.o_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6104__A (.DIODE(\core_1.decode.o_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__A (.DIODE(\core_1.decode.o_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3560__A (.DIODE(\core_1.decode.o_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3521__B (.DIODE(\core_1.decode.o_submit ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__B (.DIODE(\core_1.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4466__A (.DIODE(\core_1.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4441__A (.DIODE(\core_1.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4411__A (.DIODE(\core_1.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4382__A (.DIODE(\core_1.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4381__A1 (.DIODE(\core_1.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4380__A (.DIODE(\core_1.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3665__A (.DIODE(\core_1.decode.oc_alu_mode[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__B2 (.DIODE(\core_1.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__A1 (.DIODE(\core_1.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__B2 (.DIODE(\core_1.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5460__B2 (.DIODE(\core_1.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__B2 (.DIODE(\core_1.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5237__B2 (.DIODE(\core_1.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5158__B1 (.DIODE(\core_1.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__C (.DIODE(\core_1.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3686__A (.DIODE(\core_1.decode.oc_alu_mode[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5458__A (.DIODE(\core_1.decode.oc_alu_mode[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5151__A (.DIODE(\core_1.decode.oc_alu_mode[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4497__A (.DIODE(\core_1.decode.oc_alu_mode[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__C (.DIODE(\core_1.decode.oc_alu_mode[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3719__A1 (.DIODE(\core_1.decode.oc_alu_mode[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5676__B1 (.DIODE(\core_1.decode.oc_alu_mode[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5462__A (.DIODE(\core_1.decode.oc_alu_mode[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__B2 (.DIODE(\core_1.decode.oc_alu_mode[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5233__B2 (.DIODE(\core_1.decode.oc_alu_mode[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5155__A (.DIODE(\core_1.decode.oc_alu_mode[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4500__B2 (.DIODE(\core_1.decode.oc_alu_mode[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4495__A (.DIODE(\core_1.decode.oc_alu_mode[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3621__A (.DIODE(\core_1.decode.oc_alu_mode[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5494__A1 (.DIODE(\core_1.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5388__A (.DIODE(\core_1.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5285__C1 (.DIODE(\core_1.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5235__A (.DIODE(\core_1.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4499__B2 (.DIODE(\core_1.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__B (.DIODE(\core_1.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3677__A (.DIODE(\core_1.decode.oc_alu_mode[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5616__A1 (.DIODE(\core_1.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5589__A1 (.DIODE(\core_1.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5492__A1 (.DIODE(\core_1.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__A1 (.DIODE(\core_1.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__A1 (.DIODE(\core_1.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5236__A1 (.DIODE(\core_1.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4498__A1 (.DIODE(\core_1.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4494__A (.DIODE(\core_1.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3695__A (.DIODE(\core_1.decode.oc_alu_mode[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5617__A1 (.DIODE(\core_1.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5590__B2 (.DIODE(\core_1.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5493__A1 (.DIODE(\core_1.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5459__B2 (.DIODE(\core_1.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5316__C1 (.DIODE(\core_1.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5286__C1 (.DIODE(\core_1.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5153__B2 (.DIODE(\core_1.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4496__A (.DIODE(\core_1.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3656__A (.DIODE(\core_1.decode.oc_alu_mode[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5759__A0 (.DIODE(\core_1.ew_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5192__A0 (.DIODE(\core_1.ew_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__A0 (.DIODE(\core_1.ew_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__A (.DIODE(\core_1.ew_data[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5766__A0 (.DIODE(\core_1.ew_data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5212__A0 (.DIODE(\core_1.ew_data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__A0 (.DIODE(\core_1.ew_data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__A (.DIODE(\core_1.ew_data[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5771__A0 (.DIODE(\core_1.ew_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5257__A0 (.DIODE(\core_1.ew_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3876__A0 (.DIODE(\core_1.ew_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__A (.DIODE(\core_1.ew_data[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5776__A0 (.DIODE(\core_1.ew_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5295__A0 (.DIODE(\core_1.ew_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3878__A0 (.DIODE(\core_1.ew_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__A (.DIODE(\core_1.ew_data[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5782__A0 (.DIODE(\core_1.ew_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5332__A0 (.DIODE(\core_1.ew_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3880__A0 (.DIODE(\core_1.ew_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__A (.DIODE(\core_1.ew_data[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5787__A0 (.DIODE(\core_1.ew_data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5369__A0 (.DIODE(\core_1.ew_data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3882__A0 (.DIODE(\core_1.ew_data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__A (.DIODE(\core_1.ew_data[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5792__A0 (.DIODE(\core_1.ew_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5406__A0 (.DIODE(\core_1.ew_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3884__A0 (.DIODE(\core_1.ew_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__A (.DIODE(\core_1.ew_data[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5797__A0 (.DIODE(\core_1.ew_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5442__A0 (.DIODE(\core_1.ew_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3886__A0 (.DIODE(\core_1.ew_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__A (.DIODE(\core_1.ew_data[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5475__A (.DIODE(\core_1.ew_data[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3874__A1 (.DIODE(\core_1.ew_data[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5802__A_N (.DIODE(\core_1.ew_mem_width ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5750__A0 (.DIODE(\core_1.ew_mem_width ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3888__B_N (.DIODE(\core_1.ew_mem_width ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3853__B (.DIODE(\core_1.ew_mem_width ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6062__A (.DIODE(\core_1.ew_reg_ie[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6061__A (.DIODE(\core_1.ew_reg_ie[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5732__A0 (.DIODE(\core_1.ew_reg_ie[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__A0 (.DIODE(\core_1.ew_reg_ie[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3544__B2 (.DIODE(\core_1.ew_reg_ie[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5987__A (.DIODE(\core_1.ew_reg_ie[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5986__A (.DIODE(\core_1.ew_reg_ie[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5736__A0 (.DIODE(\core_1.ew_reg_ie[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__A2 (.DIODE(\core_1.ew_reg_ie[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3543__B (.DIODE(\core_1.ew_reg_ie[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3529__A (.DIODE(\core_1.ew_reg_ie[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5950__A (.DIODE(\core_1.ew_reg_ie[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5949__A (.DIODE(\core_1.ew_reg_ie[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5738__A0 (.DIODE(\core_1.ew_reg_ie[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3552__A3 (.DIODE(\core_1.ew_reg_ie[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3545__A1 (.DIODE(\core_1.ew_reg_ie[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3534__A2 (.DIODE(\core_1.ew_reg_ie[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5912__A (.DIODE(\core_1.ew_reg_ie[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5911__A (.DIODE(\core_1.ew_reg_ie[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5740__A0 (.DIODE(\core_1.ew_reg_ie[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__A0 (.DIODE(\core_1.ew_reg_ie[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3547__B2 (.DIODE(\core_1.ew_reg_ie[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__A3 (.DIODE(\core_1.ew_reg_ie[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5874__A (.DIODE(\core_1.ew_reg_ie[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5873__A (.DIODE(\core_1.ew_reg_ie[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5742__A0 (.DIODE(\core_1.ew_reg_ie[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__A1 (.DIODE(\core_1.ew_reg_ie[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3547__A1 (.DIODE(\core_1.ew_reg_ie[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__A0 (.DIODE(\core_1.ew_reg_ie[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5837__A (.DIODE(\core_1.ew_reg_ie[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5836__A (.DIODE(\core_1.ew_reg_ie[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5744__A0 (.DIODE(\core_1.ew_reg_ie[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__A2 (.DIODE(\core_1.ew_reg_ie[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3546__B (.DIODE(\core_1.ew_reg_ie[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__A1 (.DIODE(\core_1.ew_reg_ie[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5761__A (.DIODE(\core_1.ew_reg_ie[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5757__A (.DIODE(\core_1.ew_reg_ie[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5746__A0 (.DIODE(\core_1.ew_reg_ie[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3553__A3 (.DIODE(\core_1.ew_reg_ie[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3550__A1 (.DIODE(\core_1.ew_reg_ie[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3538__A2 (.DIODE(\core_1.ew_reg_ie[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6466__A1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__A1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__A2 (.DIODE(\core_1.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__A2 (.DIODE(\core_1.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__A1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3922__A1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__A2 (.DIODE(\core_1.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__A1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6469__A1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5201__A (.DIODE(\core_1.execute.alu_flag_reg.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4480__A (.DIODE(\core_1.execute.alu_flag_reg.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3921__A0 (.DIODE(\core_1.execute.alu_flag_reg.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3918__A1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3915__C1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6472__A1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__A1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3929__A1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3925__A1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3924__A0 (.DIODE(\core_1.execute.alu_flag_reg.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3921__A1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6479__A1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5301__A1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3916__A1 (.DIODE(\core_1.execute.alu_flag_reg.o_d[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6177__S0 (.DIODE(\core_1.execute.alu_mul_div.cbit[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6136__A (.DIODE(\core_1.execute.alu_mul_div.cbit[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6130__A (.DIODE(\core_1.execute.alu_mul_div.cbit[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4819__A (.DIODE(\core_1.execute.alu_mul_div.cbit[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4809__A (.DIODE(\core_1.execute.alu_mul_div.cbit[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4803__A (.DIODE(\core_1.execute.alu_mul_div.cbit[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4154__A (.DIODE(\core_1.execute.alu_mul_div.cbit[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5185__A2 (.DIODE(\core_1.execute.alu_mul_div.div_cur[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4825__A0 (.DIODE(\core_1.execute.alu_mul_div.div_cur[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4704__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4699__A (.DIODE(\core_1.execute.alu_mul_div.div_cur[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4697__A (.DIODE(\core_1.execute.alu_mul_div.div_cur[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4662__B1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4798__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4794__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4788__B (.DIODE(\core_1.execute.alu_mul_div.div_cur[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4686__B_N (.DIODE(\core_1.execute.alu_mul_div.div_cur[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4636__A_N (.DIODE(\core_1.execute.alu_mul_div.div_cur[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5686__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4799__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4688__A (.DIODE(\core_1.execute.alu_mul_div.div_cur[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4635__A (.DIODE(\core_1.execute.alu_mul_div.div_cur[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4715__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4707__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4663__A (.DIODE(\core_1.execute.alu_mul_div.div_cur[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4661__B1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4624__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5242__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4723__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4716__A1 (.DIODE(\core_1.execute.alu_mul_div.div_cur[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4666__A (.DIODE(\core_1.execute.alu_mul_div.div_cur[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4660__A (.DIODE(\core_1.execute.alu_mul_div.div_cur[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5683__B1 (.DIODE(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__C1 (.DIODE(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5536__B1 (.DIODE(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5437__B1 (.DIODE(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5364__B1 (.DIODE(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__A2 (.DIODE(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5183__B1 (.DIODE(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4622__B1 (.DIODE(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3675__A (.DIODE(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__A (.DIODE(\core_1.execute.alu_mul_div.i_div ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5661__A2 (.DIODE(\core_1.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5599__A2 (.DIODE(\core_1.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5538__A2 (.DIODE(\core_1.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5470__A2 (.DIODE(\core_1.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5439__A2 (.DIODE(\core_1.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5403__A2 (.DIODE(\core_1.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5184__C1 (.DIODE(\core_1.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4363__A (.DIODE(\core_1.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3681__A (.DIODE(\core_1.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3559__B (.DIODE(\core_1.execute.alu_mul_div.i_mod ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5215__A (.DIODE(\core_1.execute.alu_mul_div.i_mul ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5181__A (.DIODE(\core_1.execute.alu_mul_div.i_mul ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4367__A (.DIODE(\core_1.execute.alu_mul_div.i_mul ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3709__A (.DIODE(\core_1.execute.alu_mul_div.i_mul ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3561__B (.DIODE(\core_1.execute.alu_mul_div.i_mul ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6253__A1 (.DIODE(\core_1.execute.alu_mul_div.mul_res[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6248__A (.DIODE(\core_1.execute.alu_mul_div.mul_res[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6247__A (.DIODE(\core_1.execute.alu_mul_div.mul_res[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5561__A2 (.DIODE(\core_1.execute.alu_mul_div.mul_res[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6264__A (.DIODE(\core_1.execute.alu_mul_div.mul_res[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6259__A (.DIODE(\core_1.execute.alu_mul_div.mul_res[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6258__A (.DIODE(\core_1.execute.alu_mul_div.mul_res[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5598__A2 (.DIODE(\core_1.execute.alu_mul_div.mul_res[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6276__A1 (.DIODE(\core_1.execute.alu_mul_div.mul_res[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6271__A (.DIODE(\core_1.execute.alu_mul_div.mul_res[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6270__A (.DIODE(\core_1.execute.alu_mul_div.mul_res[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5623__A2 (.DIODE(\core_1.execute.alu_mul_div.mul_res[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6285__A1 (.DIODE(\core_1.execute.alu_mul_div.mul_res[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6277__A (.DIODE(\core_1.execute.alu_mul_div.mul_res[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5659__A2 (.DIODE(\core_1.execute.alu_mul_div.mul_res[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6638__A1 (.DIODE(\core_1.execute.irq_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6632__A1 (.DIODE(\core_1.execute.irq_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6101__B1 (.DIODE(\core_1.execute.irq_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__A1 (.DIODE(\core_1.execute.irq_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3497__B1 (.DIODE(\core_1.execute.irq_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6707__A1 (.DIODE(\core_1.execute.pc_high_buff_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6655__A1 (.DIODE(\core_1.execute.pc_high_buff_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__A (.DIODE(\core_1.execute.pc_high_buff_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6713__A1 (.DIODE(\core_1.execute.pc_high_buff_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6668__A1 (.DIODE(\core_1.execute.pc_high_buff_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__B2 (.DIODE(\core_1.execute.pc_high_buff_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6719__A1 (.DIODE(\core_1.execute.pc_high_buff_out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6680__A1 (.DIODE(\core_1.execute.pc_high_buff_out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5336__B2 (.DIODE(\core_1.execute.pc_high_buff_out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__D (.DIODE(\core_1.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6653__B (.DIODE(\core_1.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__B (.DIODE(\core_1.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6651__A1 (.DIODE(\core_1.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6647__A (.DIODE(\core_1.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5134__B2 (.DIODE(\core_1.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3516__A (.DIODE(\core_1.execute.pc_high_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__C (.DIODE(\core_1.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6658__A1 (.DIODE(\core_1.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6653__A (.DIODE(\core_1.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6652__A (.DIODE(\core_1.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5202__A (.DIODE(\core_1.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3506__A (.DIODE(\core_1.execute.pc_high_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__B (.DIODE(\core_1.execute.pc_high_out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6659__A (.DIODE(\core_1.execute.pc_high_out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5247__A1 (.DIODE(\core_1.execute.pc_high_out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__A (.DIODE(\core_1.execute.pc_high_out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6670__A1 (.DIODE(\core_1.execute.pc_high_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6666__B1_N (.DIODE(\core_1.execute.pc_high_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6665__A (.DIODE(\core_1.execute.pc_high_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5262__B2 (.DIODE(\core_1.execute.pc_high_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__A (.DIODE(\core_1.execute.pc_high_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6682__A1 (.DIODE(\core_1.execute.pc_high_out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6678__B1 (.DIODE(\core_1.execute.pc_high_out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6677__A (.DIODE(\core_1.execute.pc_high_out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__B2 (.DIODE(\core_1.execute.pc_high_out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3509__A (.DIODE(\core_1.execute.pc_high_out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6695__A1 (.DIODE(\core_1.execute.pc_high_out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6691__A (.DIODE(\core_1.execute.pc_high_out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5411__B2 (.DIODE(\core_1.execute.pc_high_out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__A (.DIODE(\core_1.execute.pc_high_out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6029__A (.DIODE(\core_1.execute.rf.reg_outputs[1][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5072__A (.DIODE(\core_1.execute.rf.reg_outputs[1][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__A1 (.DIODE(\core_1.execute.rf.reg_outputs[1][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3475__B2 (.DIODE(\core_1.execute.rf.reg_outputs[1][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6031__A (.DIODE(\core_1.execute.rf.reg_outputs[1][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5084__A1 (.DIODE(\core_1.execute.rf.reg_outputs[1][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4611__A1 (.DIODE(\core_1.execute.rf.reg_outputs[1][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3466__B2 (.DIODE(\core_1.execute.rf.reg_outputs[1][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6035__A (.DIODE(\core_1.execute.rf.reg_outputs[1][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5096__A1 (.DIODE(\core_1.execute.rf.reg_outputs[1][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__A1 (.DIODE(\core_1.execute.rf.reg_outputs[1][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3452__B2 (.DIODE(\core_1.execute.rf.reg_outputs[1][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6041__A (.DIODE(\core_1.execute.rf.reg_outputs[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5115__A1 (.DIODE(\core_1.execute.rf.reg_outputs[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__A1 (.DIODE(\core_1.execute.rf.reg_outputs[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3430__D (.DIODE(\core_1.execute.rf.reg_outputs[1][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6012__A1 (.DIODE(\core_1.execute.rf.reg_outputs[2][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4505__B2 (.DIODE(\core_1.execute.rf.reg_outputs[2][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3408__A1 (.DIODE(\core_1.execute.rf.reg_outputs[2][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6016__A1 (.DIODE(\core_1.execute.rf.reg_outputs[2][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__B2 (.DIODE(\core_1.execute.rf.reg_outputs[2][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3392__A1 (.DIODE(\core_1.execute.rf.reg_outputs[2][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6019__A1 (.DIODE(\core_1.execute.rf.reg_outputs[2][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__B2 (.DIODE(\core_1.execute.rf.reg_outputs[2][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3385__A1 (.DIODE(\core_1.execute.rf.reg_outputs[2][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5995__A (.DIODE(\core_1.execute.rf.reg_outputs[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4601__B2 (.DIODE(\core_1.execute.rf.reg_outputs[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3462__A1 (.DIODE(\core_1.execute.rf.reg_outputs[2][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6002__A (.DIODE(\core_1.execute.rf.reg_outputs[2][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__A1 (.DIODE(\core_1.execute.rf.reg_outputs[2][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3438__A1 (.DIODE(\core_1.execute.rf.reg_outputs[2][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5975__A1 (.DIODE(\core_1.execute.rf.reg_outputs[3][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__B2 (.DIODE(\core_1.execute.rf.reg_outputs[3][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3406__D (.DIODE(\core_1.execute.rf.reg_outputs[3][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5977__A1 (.DIODE(\core_1.execute.rf.reg_outputs[3][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4534__B2 (.DIODE(\core_1.execute.rf.reg_outputs[3][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3398__D (.DIODE(\core_1.execute.rf.reg_outputs[3][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5979__A1 (.DIODE(\core_1.execute.rf.reg_outputs[3][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4524__A (.DIODE(\core_1.execute.rf.reg_outputs[3][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3390__D (.DIODE(\core_1.execute.rf.reg_outputs[3][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5981__A1 (.DIODE(\core_1.execute.rf.reg_outputs[3][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4540__A1 (.DIODE(\core_1.execute.rf.reg_outputs[3][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3381__D (.DIODE(\core_1.execute.rf.reg_outputs[3][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5983__A1 (.DIODE(\core_1.execute.rf.reg_outputs[3][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4549__B2 (.DIODE(\core_1.execute.rf.reg_outputs[3][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3367__A1 (.DIODE(\core_1.execute.rf.reg_outputs[3][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5985__A1 (.DIODE(\core_1.execute.rf.reg_outputs[3][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4438__B2 (.DIODE(\core_1.execute.rf.reg_outputs[3][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3359__B2 (.DIODE(\core_1.execute.rf.reg_outputs[3][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5973__A1 (.DIODE(\core_1.execute.rf.reg_outputs[3][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__B2 (.DIODE(\core_1.execute.rf.reg_outputs[3][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3415__D (.DIODE(\core_1.execute.rf.reg_outputs[3][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5914__A (.DIODE(\core_1.execute.rf.reg_outputs[4][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4389__B2 (.DIODE(\core_1.execute.rf.reg_outputs[4][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3484__A (.DIODE(\core_1.execute.rf.reg_outputs[4][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5937__A1 (.DIODE(\core_1.execute.rf.reg_outputs[4][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4504__A1 (.DIODE(\core_1.execute.rf.reg_outputs[4][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3404__B2 (.DIODE(\core_1.execute.rf.reg_outputs[4][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5941__A1 (.DIODE(\core_1.execute.rf.reg_outputs[4][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4525__A (.DIODE(\core_1.execute.rf.reg_outputs[4][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__B2 (.DIODE(\core_1.execute.rf.reg_outputs[4][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5943__A1 (.DIODE(\core_1.execute.rf.reg_outputs[4][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4541__A1 (.DIODE(\core_1.execute.rf.reg_outputs[4][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3379__A1 (.DIODE(\core_1.execute.rf.reg_outputs[4][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5945__A1 (.DIODE(\core_1.execute.rf.reg_outputs[4][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4547__A (.DIODE(\core_1.execute.rf.reg_outputs[4][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3366__A (.DIODE(\core_1.execute.rf.reg_outputs[4][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5948__A1 (.DIODE(\core_1.execute.rf.reg_outputs[4][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4436__A (.DIODE(\core_1.execute.rf.reg_outputs[4][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3355__A1 (.DIODE(\core_1.execute.rf.reg_outputs[4][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5916__A (.DIODE(\core_1.execute.rf.reg_outputs[4][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4446__B2 (.DIODE(\core_1.execute.rf.reg_outputs[4][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__B2 (.DIODE(\core_1.execute.rf.reg_outputs[4][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5918__A (.DIODE(\core_1.execute.rf.reg_outputs[4][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__B2 (.DIODE(\core_1.execute.rf.reg_outputs[4][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3467__A (.DIODE(\core_1.execute.rf.reg_outputs[4][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5920__A (.DIODE(\core_1.execute.rf.reg_outputs[4][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__B2 (.DIODE(\core_1.execute.rf.reg_outputs[4][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__B2 (.DIODE(\core_1.execute.rf.reg_outputs[4][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5922__A (.DIODE(\core_1.execute.rf.reg_outputs[4][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4593__B2 (.DIODE(\core_1.execute.rf.reg_outputs[4][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__B2 (.DIODE(\core_1.execute.rf.reg_outputs[4][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5924__A (.DIODE(\core_1.execute.rf.reg_outputs[4][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4570__B2 (.DIODE(\core_1.execute.rf.reg_outputs[4][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3444__A1 (.DIODE(\core_1.execute.rf.reg_outputs[4][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5927__A (.DIODE(\core_1.execute.rf.reg_outputs[4][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4560__B2 (.DIODE(\core_1.execute.rf.reg_outputs[4][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__A1 (.DIODE(\core_1.execute.rf.reg_outputs[4][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5929__A (.DIODE(\core_1.execute.rf.reg_outputs[4][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4577__B2 (.DIODE(\core_1.execute.rf.reg_outputs[4][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3431__A1 (.DIODE(\core_1.execute.rf.reg_outputs[4][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5935__A1 (.DIODE(\core_1.execute.rf.reg_outputs[4][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4513__A (.DIODE(\core_1.execute.rf.reg_outputs[4][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3414__A1 (.DIODE(\core_1.execute.rf.reg_outputs[4][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5876__A (.DIODE(\core_1.execute.rf.reg_outputs[5][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4384__C (.DIODE(\core_1.execute.rf.reg_outputs[5][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3487__D (.DIODE(\core_1.execute.rf.reg_outputs[5][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5899__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4503__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3404__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5904__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4527__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3388__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5906__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4542__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3377__D (.DIODE(\core_1.execute.rf.reg_outputs[5][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5878__A (.DIODE(\core_1.execute.rf.reg_outputs[5][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4448__C (.DIODE(\core_1.execute.rf.reg_outputs[5][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3474__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5881__A (.DIODE(\core_1.execute.rf.reg_outputs[5][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4608__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3469__D (.DIODE(\core_1.execute.rf.reg_outputs[5][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5883__A (.DIODE(\core_1.execute.rf.reg_outputs[5][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4600__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3458__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5885__A (.DIODE(\core_1.execute.rf.reg_outputs[5][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4596__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3451__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5887__A (.DIODE(\core_1.execute.rf.reg_outputs[5][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4568__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3445__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5889__A (.DIODE(\core_1.execute.rf.reg_outputs[5][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4564__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3439__A1 (.DIODE(\core_1.execute.rf.reg_outputs[5][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5839__A (.DIODE(\core_1.execute.rf.reg_outputs[6][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4393__B2 (.DIODE(\core_1.execute.rf.reg_outputs[6][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3483__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5862__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__B2 (.DIODE(\core_1.execute.rf.reg_outputs[6][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3405__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5864__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4533__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3397__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5866__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__B2 (.DIODE(\core_1.execute.rf.reg_outputs[6][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3389__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5868__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__B2 (.DIODE(\core_1.execute.rf.reg_outputs[6][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3378__C (.DIODE(\core_1.execute.rf.reg_outputs[6][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5870__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4548__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3363__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5872__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4437__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3345__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5841__A (.DIODE(\core_1.execute.rf.reg_outputs[6][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4452__B2 (.DIODE(\core_1.execute.rf.reg_outputs[6][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3477__C (.DIODE(\core_1.execute.rf.reg_outputs[6][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5843__A (.DIODE(\core_1.execute.rf.reg_outputs[6][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4612__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3468__C (.DIODE(\core_1.execute.rf.reg_outputs[6][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5845__A (.DIODE(\core_1.execute.rf.reg_outputs[6][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4602__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3459__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5847__A (.DIODE(\core_1.execute.rf.reg_outputs[6][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4592__B2 (.DIODE(\core_1.execute.rf.reg_outputs[6][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3452__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5849__A (.DIODE(\core_1.execute.rf.reg_outputs[6][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4571__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3447__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5851__A (.DIODE(\core_1.execute.rf.reg_outputs[6][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4559__B2 (.DIODE(\core_1.execute.rf.reg_outputs[6][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3440__B2 (.DIODE(\core_1.execute.rf.reg_outputs[6][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5853__A (.DIODE(\core_1.execute.rf.reg_outputs[6][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4576__B2 (.DIODE(\core_1.execute.rf.reg_outputs[6][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3428__C (.DIODE(\core_1.execute.rf.reg_outputs[6][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5858__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4586__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3421__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5860__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4514__A1 (.DIODE(\core_1.execute.rf.reg_outputs[6][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3412__C (.DIODE(\core_1.execute.rf.reg_outputs[6][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5814__A1 (.DIODE(\core_1.execute.rf.reg_outputs[7][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4506__A1 (.DIODE(\core_1.execute.rf.reg_outputs[7][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3407__A (.DIODE(\core_1.execute.rf.reg_outputs[7][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5822__A1 (.DIODE(\core_1.execute.rf.reg_outputs[7][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4522__A1 (.DIODE(\core_1.execute.rf.reg_outputs[7][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3391__A (.DIODE(\core_1.execute.rf.reg_outputs[7][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5827__A1 (.DIODE(\core_1.execute.rf.reg_outputs[7][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4543__A1 (.DIODE(\core_1.execute.rf.reg_outputs[7][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3382__A (.DIODE(\core_1.execute.rf.reg_outputs[7][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5768__A (.DIODE(\core_1.execute.rf.reg_outputs[7][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4447__A (.DIODE(\core_1.execute.rf.reg_outputs[7][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3476__A (.DIODE(\core_1.execute.rf.reg_outputs[7][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5778__A (.DIODE(\core_1.execute.rf.reg_outputs[7][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4599__A (.DIODE(\core_1.execute.rf.reg_outputs[7][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3461__A (.DIODE(\core_1.execute.rf.reg_outputs[7][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5810__A1 (.DIODE(\core_1.execute.rf.reg_outputs[7][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4515__A1 (.DIODE(\core_1.execute.rf.reg_outputs[7][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3416__A (.DIODE(\core_1.execute.rf.reg_outputs[7][9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6532__A1 (.DIODE(\core_1.execute.sreg_irq_pc.o_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5338__A (.DIODE(\core_1.execute.sreg_irq_pc.o_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5334__A1 (.DIODE(\core_1.execute.sreg_irq_pc.o_d[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5259__A1 (.DIODE(\core_1.execute.sreg_long_ptr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4108__B2 (.DIODE(\core_1.execute.sreg_long_ptr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3539__A (.DIODE(\core_1.execute.sreg_long_ptr_en ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6575__A1 (.DIODE(\core_1.execute.sreg_priv_control.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6574__A (.DIODE(\core_1.execute.sreg_priv_control.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5142__A1 (.DIODE(\core_1.execute.sreg_priv_control.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4101__A1 (.DIODE(\core_1.execute.sreg_priv_control.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4094__A1 (.DIODE(\core_1.execute.sreg_priv_control.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3952__A (.DIODE(\core_1.execute.sreg_priv_control.o_d[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__6587__B2 (.DIODE(\core_1.execute.trap_flag ));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__B2 (.DIODE(\core_1.execute.trap_flag ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4895__A (.DIODE(\core_1.execute.trap_flag ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3589__S (.DIODE(\core_1.fetch.out_buffer_valid ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3585__S (.DIODE(\core_1.fetch.out_buffer_valid ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3584__S (.DIODE(\core_1.fetch.out_buffer_valid ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3579__S (.DIODE(\core_1.fetch.out_buffer_valid ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3578__S (.DIODE(\core_1.fetch.out_buffer_valid ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3493__A (.DIODE(\core_1.fetch.out_buffer_valid ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__A0 (.DIODE(\core_1.fetch.prev_request_pc[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__C (.DIODE(\core_1.fetch.prev_request_pc[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__A2 (.DIODE(\core_1.fetch.prev_request_pc[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__B (.DIODE(\core_1.fetch.prev_request_pc[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3778__A (.DIODE(\core_1.fetch.prev_request_pc[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3738__A (.DIODE(\core_1.fetch.prev_request_pc[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4238__A0 (.DIODE(\core_1.fetch.prev_request_pc[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__B (.DIODE(\core_1.fetch.prev_request_pc[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__A1 (.DIODE(\core_1.fetch.prev_request_pc[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3782__A (.DIODE(\core_1.fetch.prev_request_pc[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3737__A (.DIODE(\core_1.fetch.prev_request_pc[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__A0 (.DIODE(\core_1.fetch.prev_request_pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3787__A (.DIODE(\core_1.fetch.prev_request_pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3786__B1 (.DIODE(\core_1.fetch.prev_request_pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3736__A (.DIODE(\core_1.fetch.prev_request_pc[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__A0 (.DIODE(\core_1.fetch.prev_request_pc[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__A1 (.DIODE(\core_1.fetch.prev_request_pc[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__B (.DIODE(\core_1.fetch.prev_request_pc[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3797__A (.DIODE(\core_1.fetch.prev_request_pc[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3734__A (.DIODE(\core_1.fetch.prev_request_pc[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__A0 (.DIODE(\core_1.fetch.prev_request_pc[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3802__B1 (.DIODE(\core_1.fetch.prev_request_pc[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3801__A (.DIODE(\core_1.fetch.prev_request_pc[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__3733__A (.DIODE(\core_1.fetch.prev_request_pc[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_i_clk_A (.DIODE(i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(i_core_int_sreg[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(i_core_int_sreg[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(i_core_int_sreg[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(i_core_int_sreg[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(i_core_int_sreg[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(i_core_int_sreg[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(i_core_int_sreg[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(i_core_int_sreg[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(i_core_int_sreg[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(i_core_int_sreg[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(i_core_int_sreg[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(i_core_int_sreg[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(i_core_int_sreg[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(i_core_int_sreg[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(i_core_int_sreg[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(i_core_int_sreg[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(i_disable));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(i_irq));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(i_mc_core_int));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(i_mem_ack));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(i_mem_data[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(i_mem_data[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(i_mem_data[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(i_mem_data[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(i_mem_data[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(i_mem_data[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(i_mem_data[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(i_mem_data[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(i_mem_data[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(i_mem_data[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(i_mem_data[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(i_mem_data[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(i_mem_data[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(i_mem_data[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(i_mem_data[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(i_mem_data[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(i_mem_exception));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(i_req_data[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(i_req_data[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(i_req_data[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(i_req_data[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(i_req_data[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(i_req_data[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(i_req_data[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(i_req_data[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(i_req_data[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(i_req_data[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(i_req_data[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(i_req_data[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(i_req_data[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(i_req_data[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(i_req_data[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(i_req_data[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(i_req_data[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(i_req_data[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(i_req_data[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(i_req_data[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(i_req_data[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(i_req_data[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(i_req_data[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(i_req_data[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(i_req_data[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(i_req_data[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(i_req_data[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(i_req_data[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(i_req_data[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(i_req_data[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(i_req_data[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(i_req_data[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(i_req_data_valid));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(i_rst));
 sky130_fd_sc_hd__diode_2 ANTENNA__5129__B2 (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__5511__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__5565__A1 (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__5576__A1 (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__5626__B2 (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__5638__B2 (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__5688__A1 (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__5200__A1 (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__5245__B2 (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA__5261__A1 (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__5298__A1 (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA__5335__A1 (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__5375__A1 (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA__5413__A1 (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__5445__A1 (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__5501__A1 (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__5755__A1 (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__3557__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__A1 (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__5829__A1_N (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__A0 (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__5833__A1_N (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__A0 (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__A1 (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA__5770__A1 (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA__5775__A1 (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA__5781__A1 (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA__5786__A1 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__5791__A1 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA__5796__A1 (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__5805__A1_N (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__5758__A0 (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA__5808__A1_N (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__5765__A0 (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__6570__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6566__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6562__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6558__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6553__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6549__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6545__S (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__6503__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__4347__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__3498__A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA__4166__A0 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__3571__A0 (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__4187__A0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__3768__A0 (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__4292__A0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__4189__A0 (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA__4230__A0 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__3727__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__3592__A2 (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__4340__B (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__4232__A1 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__4163__D_N (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3892__A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3851__S (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__3570__A2 (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA__4102__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3650__B (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA__3491__A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_output72_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__6504__A0 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__B (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__6343__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5144__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__5128__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__4848__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__4628__A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA__3780__A1 (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_output73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__6549__A0 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__6408__A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__6407__B1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__5513__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__4874__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__3828__A1 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__6553__A0 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__6427__B (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__6415__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__6414__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__5564__A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__4876__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__3833__A1 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__6558__A0 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__6427__A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__6422__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__6421__B2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__5578__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__4878__A1 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__3836__A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_output76_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__6562__A0 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__6431__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__6430__A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__5629__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__4880__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__3842__A1 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_output77_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6642__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6566__A0 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6440__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__6439__A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__5641__A1_N (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__4882__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__3846__A1 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_output78_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__6570__A0 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__6445__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__6444__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__5690__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__4884__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__3850__A1 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_output79_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__6511__A0 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__C (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__B (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5196__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__5195__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4854__A1 (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4630__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__4629__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA__3784__A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_output80_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__6516__A0 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__6359__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__6348__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__6347__A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__5249__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__4856__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__3791__A1 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_output81_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6520__A0 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__B (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6360__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__6358__A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__5264__A1_N (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__4858__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA__3796__A1 (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_output82_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__6524__A0 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__6425__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__B (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__6366__A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__5302__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__4860__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA__3800__A1 (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_output83_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__6529__A0 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__6427__C (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__6372__A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__6371__B1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__5337__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__4862__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA__3805__A1 (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_output84_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__6533__A0 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__6426__C (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__6388__B (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__6381__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__6380__A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__5376__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__4864__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA__3810__A1 (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_output85_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__6537__A0 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__6426__B (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__6388__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__6387__A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__5414__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__4866__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA__3814__A1 (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_output86_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6541__A0 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6426__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6408__C (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6407__A2 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6395__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__6394__A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__5447__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__4868__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA__3819__A1 (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_output87_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6545__A0 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6428__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6408__B (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6407__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__6401__A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__5503__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__4872__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA__3824__A1 (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_output88_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__6064__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__4396__A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__4378__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__4374__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__3489__A1 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_output89_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__6087__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__4507__A1 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA__3409__B2 (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_output90_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__6090__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4801__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__4535__A1 (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA__3401__A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_output91_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__6092__A1 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__4528__B2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__3393__A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_output92_A (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__6094__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__4544__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__3386__A1 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA_output93_A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__6096__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__4812__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__4551__A1 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__3369__A (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA_output94_A (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__6098__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4800__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__4440__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__3361__A1 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA_output95_A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6137__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__6066__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__4454__A1 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__3479__A (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA_output96_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__6069__A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__4613__A1 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA__3472__B2 (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_output97_A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__6071__A (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__4604__A1 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__3463__B2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA_output98_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__6073__A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4916__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__4598__A1 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA__3456__B2 (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_output99_A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__6075__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__4572__B2 (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA__3448__A (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 ANTENNA_output100_A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__6077__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__4912__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__4566__A1 (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA__3441__A (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 ANTENNA_output101_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__6079__A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__4580__A1 (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA__3435__A1_N (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_output102_A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__6083__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4813__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__4588__A1 (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA__3425__A (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 ANTENNA_output103_A (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__6085__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__4516__B2 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA__3418__A1 (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 ANTENNA_output104_A (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA__4844__A1 (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 ANTENNA_output105_A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__5244__B2 (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3507__B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3504__B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3502__A (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA__3501__B (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 ANTENNA_output106_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__6585__A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__5137__B2 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3945__A1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA__3944__B1 (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_output109_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_output110_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_output111_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_output112_A (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 ANTENNA_output113_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_output114_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_output115_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA__6724__A1 (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_output120_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA__5727__A0 (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_output121_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA__5729__A0 (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_output135_A (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA__5102__A1 (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 ANTENNA_output136_A (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA__5107__A0 (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 ANTENNA_output137_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA__5113__A0 (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_output138_A (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA__5119__A0 (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 ANTENNA_output155_A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__5752__A0 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__3894__A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_output156_A (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__3558__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA_output157_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3872__S (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3870__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3868__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3866__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3864__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3862__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3860__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3858__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__3856__B (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_output161_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__A1 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_output168_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__4238__A1 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_output169_A (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__A1 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA_output177_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4341__B1 (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4250__S (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4248__S (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4246__S (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4244__S (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4242__S (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4240__S (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4238__S (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA__4236__S (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout211_A (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__3956__A0 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA_output179_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__4403__A0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3977__A0 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__C (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_output180_A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4640__A (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__A0 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3979__A0 (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__B (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 ANTENNA_output181_A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__4423__A (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__3981__A0 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__B (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA_output182_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__A0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3983__A0 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_output183_A (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__A0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__3985__A0 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__D (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA_output184_A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__A0 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__4408__A (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__3987__A0 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__3906__C (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA_output185_A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__D (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__4368__A (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3958__A0 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__A_N (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA_output186_A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5138__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__B (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__A0 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3960__A0 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__3902__A (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA_output187_A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5131__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5123__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__5121__A_N (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__4416__A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3962__A0 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__3904__A_N (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_output188_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__4419__A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__3964__A0 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__B (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_output189_A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__4412__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__3966__A0 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__A (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA_output190_A (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__A0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3968__A0 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__D (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA_output191_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__A0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3970__A0 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__3903__C (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_output192_A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__5125__A_N (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__4406__A0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3972__A0 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3942__A (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__3907__B_N (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA_output193_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__4405__A0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3974__A0 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__3905__A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_output194_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6703__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6650__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6576__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__6341__A1 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA__5191__A0 (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_output196_A (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__5573__A0 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA__4404__A1 (.DIODE(net196));
 sky130_fd_sc_hd__diode_2 ANTENNA_output198_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__6433__B1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__5634__A0 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA__4422__A1 (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_output199_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__5663__A0 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__4402__A1 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_output200_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__6446__B1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__5695__A0 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__4905__A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_output201_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__6706__A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__6656__A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__6579__A1 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__5210__A0 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_output202_A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6709__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__6582__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__5256__A0 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__4463__A1 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_output203_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__6712__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__6669__A1 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__5294__A0 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_output204_A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6715__A1 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__6496__A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__5331__A0 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_output205_A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6718__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__6681__A1 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__5368__A0 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_output206_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__6721__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__5405__A0 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__4399__A1 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_output207_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__6694__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__5441__A0 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__4398__A1 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_output178_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5198__B (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5197__B (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5141__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5139__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5135__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__5126__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__4377__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__4091__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__3900__A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__6991__CLK (.DIODE(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6989__CLK (.DIODE(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6757__CLK (.DIODE(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6754__CLK (.DIODE(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6751__CLK (.DIODE(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6750__CLK (.DIODE(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6753__CLK (.DIODE(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6849__CLK (.DIODE(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6744__CLK (.DIODE(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6893__CLK (.DIODE(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6887__CLK (.DIODE(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6890__CLK (.DIODE(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7102__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7103__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7099__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7098__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7101__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7097__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6755__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6756__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6992__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6994__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6993__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7100__CLK (.DIODE(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7071__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7072__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7069__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7007__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7006__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7068__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7003__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7066__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7067__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7002__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7065__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7001__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7070__CLK (.DIODE(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7087__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7088__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7081__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7085__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7086__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7008__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7005__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7034__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7038__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7040__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7039__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7036__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7037__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7033__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7049__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7052__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7050__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7004__CLK (.DIODE(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7015__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7064__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7016__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7048__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7024__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7056__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7019__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7020__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7051__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7022__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7017__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7018__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7054__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7021__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7053__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7035__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7082__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7055__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7023__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7083__CLK (.DIODE(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7095__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7046__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7047__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7042__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7014__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7010__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7074__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7026__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7076__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7077__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7030__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7078__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7079__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7031__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7032__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7080__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7063__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7062__CLK (.DIODE(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6855__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6988__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6990__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6995__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6748__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6749__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6747__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6760__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7104__CLK (.DIODE(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7120__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7117__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7115__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7114__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6952__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6954__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7113__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7106__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7118__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7109__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7110__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6758__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6759__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6770__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6951__CLK (.DIODE(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7093__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7108__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7105__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7111__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7112__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7107__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7122__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7125__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7123__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7128__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6861__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6859__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6858__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7116__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7126__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7119__CLK (.DIODE(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7057__CLK (.DIODE(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7058__CLK (.DIODE(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7059__CLK (.DIODE(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7061__CLK (.DIODE(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7028__CLK (.DIODE(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7027__CLK (.DIODE(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7029__CLK (.DIODE(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7075__CLK (.DIODE(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7025__CLK (.DIODE(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7011__CLK (.DIODE(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7012__CLK (.DIODE(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7009__CLK (.DIODE(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7013__CLK (.DIODE(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7043__CLK (.DIODE(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7060__CLK (.DIODE(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7041__CLK (.DIODE(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7045__CLK (.DIODE(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7044__CLK (.DIODE(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7073__CLK (.DIODE(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6808__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6857__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6826__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7121__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7127__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6741__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6868__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6733__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7124__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7092__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7091__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7089__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6740__CLK (.DIODE(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6875__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6736__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6874__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6737__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6739__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6871__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6869__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6734__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6866__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6867__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6732__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6876__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6742__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6809__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6860__CLK (.DIODE(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6816__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6814__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6819__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6817__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6818__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6820__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6823__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6822__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6824__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6821__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6873__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6735__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6870__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6738__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6872__CLK (.DIODE(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6877__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6727__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6863__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6728__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6731__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6864__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6729__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6815__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6813__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6825__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6862__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6845__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6843__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6844__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6810__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6811__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6812__CLK (.DIODE(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6865__CLK (.DIODE(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6984__CLK (.DIODE(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6968__CLK (.DIODE(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6804__CLK (.DIODE(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6730__CLK (.DIODE(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6806__CLK (.DIODE(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6969__CLK (.DIODE(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6807__CLK (.DIODE(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6805__CLK (.DIODE(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6880__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6838__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6839__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6827__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6841__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6840__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6842__CLK (.DIODE(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6985__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6966__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6983__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6964__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6982__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6931__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6963__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6981__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6879__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6972__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6828__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6803__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6802__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6878__CLK (.DIODE(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7195__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6932__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6777__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6953__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6999__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6947__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6965__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6971__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6856__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6970__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6987__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6986__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6967__CLK (.DIODE(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7218__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7147__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6853__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6955__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7217__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7216__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6882__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6766__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6996__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6829__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6883__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6933__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7197__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7196__CLK (.DIODE(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7198__CLK (.DIODE(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7199__CLK (.DIODE(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6790__CLK (.DIODE(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6792__CLK (.DIODE(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6788__CLK (.DIODE(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7221__CLK (.DIODE(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6791__CLK (.DIODE(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6789__CLK (.DIODE(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7219__CLK (.DIODE(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7220__CLK (.DIODE(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6852__CLK (.DIODE(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6850__CLK (.DIODE(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6847__CLK (.DIODE(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7164__CLK (.DIODE(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7192__CLK (.DIODE(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6929__CLK (.DIODE(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7193__CLK (.DIODE(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7129__CLK (.DIODE(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7215__CLK (.DIODE(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7194__CLK (.DIODE(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6935__CLK (.DIODE(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6930__CLK (.DIODE(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6837__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6800__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6801__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6979__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6978__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7176__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7178__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6962__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6881__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6980__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6934__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7177__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7174__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7175__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7173__CLK (.DIODE(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6830__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6794__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6833__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6834__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6796__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6831__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6798__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6961__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6799__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6832__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6835__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6836__CLK (.DIODE(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7189__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6923__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7187__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7166__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7167__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7171__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7172__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6960__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6959__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6797__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6958__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7168__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6795__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6977__CLK (.DIODE(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6924__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6940__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6942__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7242__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6921__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6925__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6946__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6926__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6927__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6948__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6973__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6974__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6928__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6922__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6949__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6975__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6976__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6950__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6956__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7170__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6957__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7169__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7191__CLK (.DIODE(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7235__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7234__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7239__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7241__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7222__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7226__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6938__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6943__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7237__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7240__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7236__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7238__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6939__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6941__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6936__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6937__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6919__CLK (.DIODE(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7188__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7190__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7232__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7230__CLK (.DIODE(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7231__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7233__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7225__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7185__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7186__CLK (.DIODE(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7207__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7209__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7206__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7212__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6945__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6783__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6779__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6781__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7204__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7201__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7200__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6944__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7202__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6918__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7223__CLK (.DIODE(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6920__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7210__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7208__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6782__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6998__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7180__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7179__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7181__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7183__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6780__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6784__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7213__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6907__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7211__CLK (.DIODE(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7182__CLK (.DIODE(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6743__CLK (.DIODE(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7000__CLK (.DIODE(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6774__CLK (.DIODE(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7214__CLK (.DIODE(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6785__CLK (.DIODE(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6778__CLK (.DIODE(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7165__CLK (.DIODE(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6884__CLK (.DIODE(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7184__CLK (.DIODE(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6768__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6851__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6917__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6771__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6787__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6786__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6773__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6745__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6772__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6763__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6762__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6765__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6764__CLK (.DIODE(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6726__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6761__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6775__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6886__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6897__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6896__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6848__CLK (.DIODE(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6902__CLK (.DIODE(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6895__CLK (.DIODE(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6885__CLK (.DIODE(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6888__CLK (.DIODE(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6891__CLK (.DIODE(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6746__CLK (.DIODE(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6889__CLK (.DIODE(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6892__CLK (.DIODE(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6894__CLK (.DIODE(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6910__CLK (.DIODE(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6906__CLK (.DIODE(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6905__CLK (.DIODE(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6904__CLK (.DIODE(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6903__CLK (.DIODE(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6901__CLK (.DIODE(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6900__CLK (.DIODE(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7158__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7152__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7161__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7162__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7154__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6913__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7155__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7160__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7163__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6912__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6911__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6909__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6908__CLK (.DIODE(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7148__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6793__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7153__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7159__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7150__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7157__CLK (.DIODE(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7151__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7130__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7156__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6916__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6914__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7131__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6915__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6898__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__6899__CLK (.DIODE(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7136__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7134__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7141__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7135__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7142__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7143__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7144__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7145__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA__7133__CLK (.DIODE(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1_0_i_clk_A (.DIODE(clknet_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0_0_i_clk_A (.DIODE(clknet_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1_0_i_clk_A (.DIODE(clknet_1_0_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0_0_i_clk_A (.DIODE(clknet_1_0_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3_0_i_clk_A (.DIODE(clknet_1_1_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2_0_i_clk_A (.DIODE(clknet_1_1_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_i_clk_A (.DIODE(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_i_clk_A (.DIODE(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_i_clk_A (.DIODE(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_i_clk_A (.DIODE(clknet_2_3_0_i_clk));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_516 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_803 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_718 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_478 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_815 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_506 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_431 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_621 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_430 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_692 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_368 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_794 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_780 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_723 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_592 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_795 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_638 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_560 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_448 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_440 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_625 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_794 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_665 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_395 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_379 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_345 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_378 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_637 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_659 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_838 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_383 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_659 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_434 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_706 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_602 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_649 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_410 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_518 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_535 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_751 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_718 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_730 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_413 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_789 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_376 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_385 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_448 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_731 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_743 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_820 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_471 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_732 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_518 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_721 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_372 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_733 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_759 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_534 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_499 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_592 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_507 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_463 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_482 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_808 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_800 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_764 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_680 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_519 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_730 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_756 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_710 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_770 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_703 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_734 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_491 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_700 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_778 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_740 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_746 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_736 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_624 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_718 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_649 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_532 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_563 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_591 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_631 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_748 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_507 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_722 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_791 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_810 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_793 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_805 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_743 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_655 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_538 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_821 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_748 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_760 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_661 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_796 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_802 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_497 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_788 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_588 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_815 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_783 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_819 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_604 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_841 ();
 assign dbg_out[0] = net212;
 assign dbg_out[10] = net222;
 assign dbg_out[11] = net223;
 assign dbg_out[12] = net224;
 assign dbg_out[13] = net225;
 assign dbg_out[14] = net226;
 assign dbg_out[15] = net227;
 assign dbg_out[16] = net228;
 assign dbg_out[17] = net229;
 assign dbg_out[18] = net230;
 assign dbg_out[19] = net231;
 assign dbg_out[1] = net213;
 assign dbg_out[20] = net232;
 assign dbg_out[21] = net233;
 assign dbg_out[22] = net234;
 assign dbg_out[23] = net235;
 assign dbg_out[24] = net236;
 assign dbg_out[25] = net237;
 assign dbg_out[26] = net238;
 assign dbg_out[27] = net239;
 assign dbg_out[28] = net240;
 assign dbg_out[29] = net241;
 assign dbg_out[2] = net214;
 assign dbg_out[30] = net242;
 assign dbg_out[31] = net243;
 assign dbg_out[32] = net244;
 assign dbg_out[33] = net245;
 assign dbg_out[34] = net246;
 assign dbg_out[35] = net247;
 assign dbg_out[3] = net215;
 assign dbg_out[4] = net216;
 assign dbg_out[5] = net217;
 assign dbg_out[6] = net218;
 assign dbg_out[7] = net219;
 assign dbg_out[8] = net220;
 assign dbg_out[9] = net221;
 assign o_mem_addr_high[7] = net248;
endmodule

