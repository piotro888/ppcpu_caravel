VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO core
  CLASS BLOCK ;
  FOREIGN core ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.000 BY 800.000 ;
  PIN dbg_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 12.960 200.000 13.560 ;
    END
  END dbg_in[0]
  PIN dbg_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 23.840 200.000 24.440 ;
    END
  END dbg_in[1]
  PIN dbg_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 34.720 200.000 35.320 ;
    END
  END dbg_in[2]
  PIN dbg_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 45.600 200.000 46.200 ;
    END
  END dbg_in[3]
  PIN dbg_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 56.480 200.000 57.080 ;
    END
  END dbg_out[0]
  PIN dbg_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 165.280 200.000 165.880 ;
    END
  END dbg_out[10]
  PIN dbg_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 176.160 200.000 176.760 ;
    END
  END dbg_out[11]
  PIN dbg_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 187.040 200.000 187.640 ;
    END
  END dbg_out[12]
  PIN dbg_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 197.920 200.000 198.520 ;
    END
  END dbg_out[13]
  PIN dbg_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 208.800 200.000 209.400 ;
    END
  END dbg_out[14]
  PIN dbg_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 219.680 200.000 220.280 ;
    END
  END dbg_out[15]
  PIN dbg_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 230.560 200.000 231.160 ;
    END
  END dbg_out[16]
  PIN dbg_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 241.440 200.000 242.040 ;
    END
  END dbg_out[17]
  PIN dbg_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 252.320 200.000 252.920 ;
    END
  END dbg_out[18]
  PIN dbg_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 263.200 200.000 263.800 ;
    END
  END dbg_out[19]
  PIN dbg_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 67.360 200.000 67.960 ;
    END
  END dbg_out[1]
  PIN dbg_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 274.080 200.000 274.680 ;
    END
  END dbg_out[20]
  PIN dbg_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 284.960 200.000 285.560 ;
    END
  END dbg_out[21]
  PIN dbg_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 295.840 200.000 296.440 ;
    END
  END dbg_out[22]
  PIN dbg_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 306.720 200.000 307.320 ;
    END
  END dbg_out[23]
  PIN dbg_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 317.600 200.000 318.200 ;
    END
  END dbg_out[24]
  PIN dbg_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 328.480 200.000 329.080 ;
    END
  END dbg_out[25]
  PIN dbg_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 339.360 200.000 339.960 ;
    END
  END dbg_out[26]
  PIN dbg_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 350.240 200.000 350.840 ;
    END
  END dbg_out[27]
  PIN dbg_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 361.120 200.000 361.720 ;
    END
  END dbg_out[28]
  PIN dbg_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 372.000 200.000 372.600 ;
    END
  END dbg_out[29]
  PIN dbg_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 78.240 200.000 78.840 ;
    END
  END dbg_out[2]
  PIN dbg_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 382.880 200.000 383.480 ;
    END
  END dbg_out[30]
  PIN dbg_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 393.760 200.000 394.360 ;
    END
  END dbg_out[31]
  PIN dbg_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 404.640 200.000 405.240 ;
    END
  END dbg_out[32]
  PIN dbg_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 415.520 200.000 416.120 ;
    END
  END dbg_out[33]
  PIN dbg_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 426.400 200.000 427.000 ;
    END
  END dbg_out[34]
  PIN dbg_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 437.280 200.000 437.880 ;
    END
  END dbg_out[35]
  PIN dbg_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 89.120 200.000 89.720 ;
    END
  END dbg_out[3]
  PIN dbg_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 100.000 200.000 100.600 ;
    END
  END dbg_out[4]
  PIN dbg_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 110.880 200.000 111.480 ;
    END
  END dbg_out[5]
  PIN dbg_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 121.760 200.000 122.360 ;
    END
  END dbg_out[6]
  PIN dbg_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 132.640 200.000 133.240 ;
    END
  END dbg_out[7]
  PIN dbg_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 143.520 200.000 144.120 ;
    END
  END dbg_out[8]
  PIN dbg_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 154.400 200.000 155.000 ;
    END
  END dbg_out[9]
  PIN dbg_pc[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 448.160 200.000 448.760 ;
    END
  END dbg_pc[0]
  PIN dbg_pc[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 556.960 200.000 557.560 ;
    END
  END dbg_pc[10]
  PIN dbg_pc[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 567.840 200.000 568.440 ;
    END
  END dbg_pc[11]
  PIN dbg_pc[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 578.720 200.000 579.320 ;
    END
  END dbg_pc[12]
  PIN dbg_pc[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 589.600 200.000 590.200 ;
    END
  END dbg_pc[13]
  PIN dbg_pc[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 600.480 200.000 601.080 ;
    END
  END dbg_pc[14]
  PIN dbg_pc[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 611.360 200.000 611.960 ;
    END
  END dbg_pc[15]
  PIN dbg_pc[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 459.040 200.000 459.640 ;
    END
  END dbg_pc[1]
  PIN dbg_pc[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 469.920 200.000 470.520 ;
    END
  END dbg_pc[2]
  PIN dbg_pc[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 480.800 200.000 481.400 ;
    END
  END dbg_pc[3]
  PIN dbg_pc[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 491.680 200.000 492.280 ;
    END
  END dbg_pc[4]
  PIN dbg_pc[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 502.560 200.000 503.160 ;
    END
  END dbg_pc[5]
  PIN dbg_pc[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 513.440 200.000 514.040 ;
    END
  END dbg_pc[6]
  PIN dbg_pc[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 524.320 200.000 524.920 ;
    END
  END dbg_pc[7]
  PIN dbg_pc[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 535.200 200.000 535.800 ;
    END
  END dbg_pc[8]
  PIN dbg_pc[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 546.080 200.000 546.680 ;
    END
  END dbg_pc[9]
  PIN dbg_r0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 622.240 200.000 622.840 ;
    END
  END dbg_r0[0]
  PIN dbg_r0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 731.040 200.000 731.640 ;
    END
  END dbg_r0[10]
  PIN dbg_r0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 741.920 200.000 742.520 ;
    END
  END dbg_r0[11]
  PIN dbg_r0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 752.800 200.000 753.400 ;
    END
  END dbg_r0[12]
  PIN dbg_r0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 763.680 200.000 764.280 ;
    END
  END dbg_r0[13]
  PIN dbg_r0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 774.560 200.000 775.160 ;
    END
  END dbg_r0[14]
  PIN dbg_r0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 785.440 200.000 786.040 ;
    END
  END dbg_r0[15]
  PIN dbg_r0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 633.120 200.000 633.720 ;
    END
  END dbg_r0[1]
  PIN dbg_r0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 644.000 200.000 644.600 ;
    END
  END dbg_r0[2]
  PIN dbg_r0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 654.880 200.000 655.480 ;
    END
  END dbg_r0[3]
  PIN dbg_r0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 665.760 200.000 666.360 ;
    END
  END dbg_r0[4]
  PIN dbg_r0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 676.640 200.000 677.240 ;
    END
  END dbg_r0[5]
  PIN dbg_r0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 687.520 200.000 688.120 ;
    END
  END dbg_r0[6]
  PIN dbg_r0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 698.400 200.000 699.000 ;
    END
  END dbg_r0[7]
  PIN dbg_r0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 709.280 200.000 709.880 ;
    END
  END dbg_r0[8]
  PIN dbg_r0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 196.000 720.160 200.000 720.760 ;
    END
  END dbg_r0[9]
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.770 796.000 4.050 800.000 ;
    END
  END i_clk
  PIN i_irq
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 13.890 796.000 14.170 800.000 ;
    END
  END i_irq
  PIN i_mem_ack
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END i_mem_ack
  PIN i_mem_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END i_mem_data[0]
  PIN i_mem_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 92.520 4.000 93.120 ;
    END
  END i_mem_data[10]
  PIN i_mem_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 100.000 4.000 100.600 ;
    END
  END i_mem_data[11]
  PIN i_mem_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 107.480 4.000 108.080 ;
    END
  END i_mem_data[12]
  PIN i_mem_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 114.960 4.000 115.560 ;
    END
  END i_mem_data[13]
  PIN i_mem_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END i_mem_data[14]
  PIN i_mem_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.920 4.000 130.520 ;
    END
  END i_mem_data[15]
  PIN i_mem_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 25.200 4.000 25.800 ;
    END
  END i_mem_data[1]
  PIN i_mem_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 32.680 4.000 33.280 ;
    END
  END i_mem_data[2]
  PIN i_mem_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.160 4.000 40.760 ;
    END
  END i_mem_data[3]
  PIN i_mem_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END i_mem_data[4]
  PIN i_mem_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 55.120 4.000 55.720 ;
    END
  END i_mem_data[5]
  PIN i_mem_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 62.600 4.000 63.200 ;
    END
  END i_mem_data[6]
  PIN i_mem_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END i_mem_data[7]
  PIN i_mem_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 77.560 4.000 78.160 ;
    END
  END i_mem_data[8]
  PIN i_mem_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END i_mem_data[9]
  PIN i_mem_exception
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 137.400 4.000 138.000 ;
    END
  END i_mem_exception
  PIN i_req_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.160 4.000 414.760 ;
    END
  END i_req_data[0]
  PIN i_req_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.960 4.000 489.560 ;
    END
  END i_req_data[10]
  PIN i_req_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 496.440 4.000 497.040 ;
    END
  END i_req_data[11]
  PIN i_req_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.920 4.000 504.520 ;
    END
  END i_req_data[12]
  PIN i_req_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 511.400 4.000 512.000 ;
    END
  END i_req_data[13]
  PIN i_req_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 518.880 4.000 519.480 ;
    END
  END i_req_data[14]
  PIN i_req_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 526.360 4.000 526.960 ;
    END
  END i_req_data[15]
  PIN i_req_data[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END i_req_data[16]
  PIN i_req_data[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 541.320 4.000 541.920 ;
    END
  END i_req_data[17]
  PIN i_req_data[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 548.800 4.000 549.400 ;
    END
  END i_req_data[18]
  PIN i_req_data[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 556.280 4.000 556.880 ;
    END
  END i_req_data[19]
  PIN i_req_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END i_req_data[1]
  PIN i_req_data[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 563.760 4.000 564.360 ;
    END
  END i_req_data[20]
  PIN i_req_data[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END i_req_data[21]
  PIN i_req_data[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.720 4.000 579.320 ;
    END
  END i_req_data[22]
  PIN i_req_data[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 586.200 4.000 586.800 ;
    END
  END i_req_data[23]
  PIN i_req_data[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 593.680 4.000 594.280 ;
    END
  END i_req_data[24]
  PIN i_req_data[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 601.160 4.000 601.760 ;
    END
  END i_req_data[25]
  PIN i_req_data[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 608.640 4.000 609.240 ;
    END
  END i_req_data[26]
  PIN i_req_data[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 616.120 4.000 616.720 ;
    END
  END i_req_data[27]
  PIN i_req_data[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 623.600 4.000 624.200 ;
    END
  END i_req_data[28]
  PIN i_req_data[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 631.080 4.000 631.680 ;
    END
  END i_req_data[29]
  PIN i_req_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.120 4.000 429.720 ;
    END
  END i_req_data[2]
  PIN i_req_data[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 638.560 4.000 639.160 ;
    END
  END i_req_data[30]
  PIN i_req_data[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 646.040 4.000 646.640 ;
    END
  END i_req_data[31]
  PIN i_req_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 436.600 4.000 437.200 ;
    END
  END i_req_data[3]
  PIN i_req_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.080 4.000 444.680 ;
    END
  END i_req_data[4]
  PIN i_req_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 451.560 4.000 452.160 ;
    END
  END i_req_data[5]
  PIN i_req_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END i_req_data[6]
  PIN i_req_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 466.520 4.000 467.120 ;
    END
  END i_req_data[7]
  PIN i_req_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.000 4.000 474.600 ;
    END
  END i_req_data[8]
  PIN i_req_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 481.480 4.000 482.080 ;
    END
  END i_req_data[9]
  PIN i_req_data_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 653.520 4.000 654.120 ;
    END
  END i_req_data_valid
  PIN i_rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.830 796.000 9.110 800.000 ;
    END
  END i_rst
  PIN o_c_data_page
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 796.000 19.230 800.000 ;
    END
  END o_c_data_page
  PIN o_c_instr_page
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 24.010 796.000 24.290 800.000 ;
    END
  END o_c_instr_page
  PIN o_icache_flush
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 796.000 196.330 800.000 ;
    END
  END o_icache_flush
  PIN o_mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 144.880 4.000 145.480 ;
    END
  END o_mem_addr[0]
  PIN o_mem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END o_mem_addr[10]
  PIN o_mem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.160 4.000 227.760 ;
    END
  END o_mem_addr[11]
  PIN o_mem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END o_mem_addr[12]
  PIN o_mem_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 242.120 4.000 242.720 ;
    END
  END o_mem_addr[13]
  PIN o_mem_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END o_mem_addr[14]
  PIN o_mem_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 257.080 4.000 257.680 ;
    END
  END o_mem_addr[15]
  PIN o_mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 152.360 4.000 152.960 ;
    END
  END o_mem_addr[1]
  PIN o_mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END o_mem_addr[2]
  PIN o_mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 167.320 4.000 167.920 ;
    END
  END o_mem_addr[3]
  PIN o_mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.800 4.000 175.400 ;
    END
  END o_mem_addr[4]
  PIN o_mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 182.280 4.000 182.880 ;
    END
  END o_mem_addr[5]
  PIN o_mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.760 4.000 190.360 ;
    END
  END o_mem_addr[6]
  PIN o_mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END o_mem_addr[7]
  PIN o_mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.720 4.000 205.320 ;
    END
  END o_mem_addr[8]
  PIN o_mem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END o_mem_addr[9]
  PIN o_mem_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 4.000 265.160 ;
    END
  END o_mem_data[0]
  PIN o_mem_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 339.360 4.000 339.960 ;
    END
  END o_mem_data[10]
  PIN o_mem_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 346.840 4.000 347.440 ;
    END
  END o_mem_data[11]
  PIN o_mem_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 354.320 4.000 354.920 ;
    END
  END o_mem_data[12]
  PIN o_mem_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 361.800 4.000 362.400 ;
    END
  END o_mem_data[13]
  PIN o_mem_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.280 4.000 369.880 ;
    END
  END o_mem_data[14]
  PIN o_mem_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 376.760 4.000 377.360 ;
    END
  END o_mem_data[15]
  PIN o_mem_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END o_mem_data[1]
  PIN o_mem_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 279.520 4.000 280.120 ;
    END
  END o_mem_data[2]
  PIN o_mem_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END o_mem_data[3]
  PIN o_mem_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 294.480 4.000 295.080 ;
    END
  END o_mem_data[4]
  PIN o_mem_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END o_mem_data[5]
  PIN o_mem_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END o_mem_data[6]
  PIN o_mem_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.920 4.000 317.520 ;
    END
  END o_mem_data[7]
  PIN o_mem_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 324.400 4.000 325.000 ;
    END
  END o_mem_data[8]
  PIN o_mem_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 331.880 4.000 332.480 ;
    END
  END o_mem_data[9]
  PIN o_mem_req
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 384.240 4.000 384.840 ;
    END
  END o_mem_req
  PIN o_mem_sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.720 4.000 392.320 ;
    END
  END o_mem_sel[0]
  PIN o_mem_sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 399.200 4.000 399.800 ;
    END
  END o_mem_sel[1]
  PIN o_mem_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.680 4.000 407.280 ;
    END
  END o_mem_we
  PIN o_req_active
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 661.000 4.000 661.600 ;
    END
  END o_req_active
  PIN o_req_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 668.480 4.000 669.080 ;
    END
  END o_req_addr[0]
  PIN o_req_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 743.280 4.000 743.880 ;
    END
  END o_req_addr[10]
  PIN o_req_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 750.760 4.000 751.360 ;
    END
  END o_req_addr[11]
  PIN o_req_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 758.240 4.000 758.840 ;
    END
  END o_req_addr[12]
  PIN o_req_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.720 4.000 766.320 ;
    END
  END o_req_addr[13]
  PIN o_req_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 773.200 4.000 773.800 ;
    END
  END o_req_addr[14]
  PIN o_req_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.680 4.000 781.280 ;
    END
  END o_req_addr[15]
  PIN o_req_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 675.960 4.000 676.560 ;
    END
  END o_req_addr[1]
  PIN o_req_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 683.440 4.000 684.040 ;
    END
  END o_req_addr[2]
  PIN o_req_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 690.920 4.000 691.520 ;
    END
  END o_req_addr[3]
  PIN o_req_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 698.400 4.000 699.000 ;
    END
  END o_req_addr[4]
  PIN o_req_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 705.880 4.000 706.480 ;
    END
  END o_req_addr[5]
  PIN o_req_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 713.360 4.000 713.960 ;
    END
  END o_req_addr[6]
  PIN o_req_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 720.840 4.000 721.440 ;
    END
  END o_req_addr[7]
  PIN o_req_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 728.320 4.000 728.920 ;
    END
  END o_req_addr[8]
  PIN o_req_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 735.800 4.000 736.400 ;
    END
  END o_req_addr[9]
  PIN o_req_ppl_submit
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 788.160 4.000 788.760 ;
    END
  END o_req_ppl_submit
  PIN sr_bus_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 796.000 29.350 800.000 ;
    END
  END sr_bus_addr[0]
  PIN sr_bus_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.670 796.000 79.950 800.000 ;
    END
  END sr_bus_addr[10]
  PIN sr_bus_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.730 796.000 85.010 800.000 ;
    END
  END sr_bus_addr[11]
  PIN sr_bus_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 89.790 796.000 90.070 800.000 ;
    END
  END sr_bus_addr[12]
  PIN sr_bus_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 796.000 95.130 800.000 ;
    END
  END sr_bus_addr[13]
  PIN sr_bus_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 796.000 100.190 800.000 ;
    END
  END sr_bus_addr[14]
  PIN sr_bus_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.970 796.000 105.250 800.000 ;
    END
  END sr_bus_addr[15]
  PIN sr_bus_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 34.130 796.000 34.410 800.000 ;
    END
  END sr_bus_addr[1]
  PIN sr_bus_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.190 796.000 39.470 800.000 ;
    END
  END sr_bus_addr[2]
  PIN sr_bus_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 796.000 44.530 800.000 ;
    END
  END sr_bus_addr[3]
  PIN sr_bus_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 796.000 49.590 800.000 ;
    END
  END sr_bus_addr[4]
  PIN sr_bus_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 796.000 54.650 800.000 ;
    END
  END sr_bus_addr[5]
  PIN sr_bus_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 796.000 59.710 800.000 ;
    END
  END sr_bus_addr[6]
  PIN sr_bus_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 796.000 64.770 800.000 ;
    END
  END sr_bus_addr[7]
  PIN sr_bus_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 796.000 69.830 800.000 ;
    END
  END sr_bus_addr[8]
  PIN sr_bus_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.610 796.000 74.890 800.000 ;
    END
  END sr_bus_addr[9]
  PIN sr_bus_data_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.030 796.000 110.310 800.000 ;
    END
  END sr_bus_data_o[0]
  PIN sr_bus_data_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.630 796.000 160.910 800.000 ;
    END
  END sr_bus_data_o[10]
  PIN sr_bus_data_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 165.690 796.000 165.970 800.000 ;
    END
  END sr_bus_data_o[11]
  PIN sr_bus_data_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 796.000 171.030 800.000 ;
    END
  END sr_bus_data_o[12]
  PIN sr_bus_data_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.810 796.000 176.090 800.000 ;
    END
  END sr_bus_data_o[13]
  PIN sr_bus_data_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.870 796.000 181.150 800.000 ;
    END
  END sr_bus_data_o[14]
  PIN sr_bus_data_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.930 796.000 186.210 800.000 ;
    END
  END sr_bus_data_o[15]
  PIN sr_bus_data_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.090 796.000 115.370 800.000 ;
    END
  END sr_bus_data_o[1]
  PIN sr_bus_data_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 796.000 120.430 800.000 ;
    END
  END sr_bus_data_o[2]
  PIN sr_bus_data_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 796.000 125.490 800.000 ;
    END
  END sr_bus_data_o[3]
  PIN sr_bus_data_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 130.270 796.000 130.550 800.000 ;
    END
  END sr_bus_data_o[4]
  PIN sr_bus_data_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 796.000 135.610 800.000 ;
    END
  END sr_bus_data_o[5]
  PIN sr_bus_data_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.390 796.000 140.670 800.000 ;
    END
  END sr_bus_data_o[6]
  PIN sr_bus_data_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 796.000 145.730 800.000 ;
    END
  END sr_bus_data_o[7]
  PIN sr_bus_data_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 796.000 150.790 800.000 ;
    END
  END sr_bus_data_o[8]
  PIN sr_bus_data_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.570 796.000 155.850 800.000 ;
    END
  END sr_bus_data_o[9]
  PIN sr_bus_we
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.990 796.000 191.270 800.000 ;
    END
  END sr_bus_we
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 789.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 789.040 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 789.040 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 194.120 788.885 ;
      LAYER met1 ;
        RECT 0.990 10.640 199.570 789.440 ;
      LAYER met2 ;
        RECT 1.010 795.720 3.490 796.690 ;
        RECT 4.330 795.720 8.550 796.690 ;
        RECT 9.390 795.720 13.610 796.690 ;
        RECT 14.450 795.720 18.670 796.690 ;
        RECT 19.510 795.720 23.730 796.690 ;
        RECT 24.570 795.720 28.790 796.690 ;
        RECT 29.630 795.720 33.850 796.690 ;
        RECT 34.690 795.720 38.910 796.690 ;
        RECT 39.750 795.720 43.970 796.690 ;
        RECT 44.810 795.720 49.030 796.690 ;
        RECT 49.870 795.720 54.090 796.690 ;
        RECT 54.930 795.720 59.150 796.690 ;
        RECT 59.990 795.720 64.210 796.690 ;
        RECT 65.050 795.720 69.270 796.690 ;
        RECT 70.110 795.720 74.330 796.690 ;
        RECT 75.170 795.720 79.390 796.690 ;
        RECT 80.230 795.720 84.450 796.690 ;
        RECT 85.290 795.720 89.510 796.690 ;
        RECT 90.350 795.720 94.570 796.690 ;
        RECT 95.410 795.720 99.630 796.690 ;
        RECT 100.470 795.720 104.690 796.690 ;
        RECT 105.530 795.720 109.750 796.690 ;
        RECT 110.590 795.720 114.810 796.690 ;
        RECT 115.650 795.720 119.870 796.690 ;
        RECT 120.710 795.720 124.930 796.690 ;
        RECT 125.770 795.720 129.990 796.690 ;
        RECT 130.830 795.720 135.050 796.690 ;
        RECT 135.890 795.720 140.110 796.690 ;
        RECT 140.950 795.720 145.170 796.690 ;
        RECT 146.010 795.720 150.230 796.690 ;
        RECT 151.070 795.720 155.290 796.690 ;
        RECT 156.130 795.720 160.350 796.690 ;
        RECT 161.190 795.720 165.410 796.690 ;
        RECT 166.250 795.720 170.470 796.690 ;
        RECT 171.310 795.720 175.530 796.690 ;
        RECT 176.370 795.720 180.590 796.690 ;
        RECT 181.430 795.720 185.650 796.690 ;
        RECT 186.490 795.720 190.710 796.690 ;
        RECT 191.550 795.720 195.770 796.690 ;
        RECT 196.610 795.720 199.940 796.690 ;
        RECT 1.010 10.355 199.940 795.720 ;
      LAYER met3 ;
        RECT 4.400 787.760 199.575 788.965 ;
        RECT 0.270 786.440 199.575 787.760 ;
        RECT 0.270 785.040 195.600 786.440 ;
        RECT 0.270 781.680 199.575 785.040 ;
        RECT 4.400 780.280 199.575 781.680 ;
        RECT 0.270 775.560 199.575 780.280 ;
        RECT 0.270 774.200 195.600 775.560 ;
        RECT 4.400 774.160 195.600 774.200 ;
        RECT 4.400 772.800 199.575 774.160 ;
        RECT 0.270 766.720 199.575 772.800 ;
        RECT 4.400 765.320 199.575 766.720 ;
        RECT 0.270 764.680 199.575 765.320 ;
        RECT 0.270 763.280 195.600 764.680 ;
        RECT 0.270 759.240 199.575 763.280 ;
        RECT 4.400 757.840 199.575 759.240 ;
        RECT 0.270 753.800 199.575 757.840 ;
        RECT 0.270 752.400 195.600 753.800 ;
        RECT 0.270 751.760 199.575 752.400 ;
        RECT 4.400 750.360 199.575 751.760 ;
        RECT 0.270 744.280 199.575 750.360 ;
        RECT 4.400 742.920 199.575 744.280 ;
        RECT 4.400 742.880 195.600 742.920 ;
        RECT 0.270 741.520 195.600 742.880 ;
        RECT 0.270 736.800 199.575 741.520 ;
        RECT 4.400 735.400 199.575 736.800 ;
        RECT 0.270 732.040 199.575 735.400 ;
        RECT 0.270 730.640 195.600 732.040 ;
        RECT 0.270 729.320 199.575 730.640 ;
        RECT 4.400 727.920 199.575 729.320 ;
        RECT 0.270 721.840 199.575 727.920 ;
        RECT 4.400 721.160 199.575 721.840 ;
        RECT 4.400 720.440 195.600 721.160 ;
        RECT 0.270 719.760 195.600 720.440 ;
        RECT 0.270 714.360 199.575 719.760 ;
        RECT 4.400 712.960 199.575 714.360 ;
        RECT 0.270 710.280 199.575 712.960 ;
        RECT 0.270 708.880 195.600 710.280 ;
        RECT 0.270 706.880 199.575 708.880 ;
        RECT 4.400 705.480 199.575 706.880 ;
        RECT 0.270 699.400 199.575 705.480 ;
        RECT 4.400 698.000 195.600 699.400 ;
        RECT 0.270 691.920 199.575 698.000 ;
        RECT 4.400 690.520 199.575 691.920 ;
        RECT 0.270 688.520 199.575 690.520 ;
        RECT 0.270 687.120 195.600 688.520 ;
        RECT 0.270 684.440 199.575 687.120 ;
        RECT 4.400 683.040 199.575 684.440 ;
        RECT 0.270 677.640 199.575 683.040 ;
        RECT 0.270 676.960 195.600 677.640 ;
        RECT 4.400 676.240 195.600 676.960 ;
        RECT 4.400 675.560 199.575 676.240 ;
        RECT 0.270 669.480 199.575 675.560 ;
        RECT 4.400 668.080 199.575 669.480 ;
        RECT 0.270 666.760 199.575 668.080 ;
        RECT 0.270 665.360 195.600 666.760 ;
        RECT 0.270 662.000 199.575 665.360 ;
        RECT 4.400 660.600 199.575 662.000 ;
        RECT 0.270 655.880 199.575 660.600 ;
        RECT 0.270 654.520 195.600 655.880 ;
        RECT 4.400 654.480 195.600 654.520 ;
        RECT 4.400 653.120 199.575 654.480 ;
        RECT 0.270 647.040 199.575 653.120 ;
        RECT 4.400 645.640 199.575 647.040 ;
        RECT 0.270 645.000 199.575 645.640 ;
        RECT 0.270 643.600 195.600 645.000 ;
        RECT 0.270 639.560 199.575 643.600 ;
        RECT 4.400 638.160 199.575 639.560 ;
        RECT 0.270 634.120 199.575 638.160 ;
        RECT 0.270 632.720 195.600 634.120 ;
        RECT 0.270 632.080 199.575 632.720 ;
        RECT 4.400 630.680 199.575 632.080 ;
        RECT 0.270 624.600 199.575 630.680 ;
        RECT 4.400 623.240 199.575 624.600 ;
        RECT 4.400 623.200 195.600 623.240 ;
        RECT 0.270 621.840 195.600 623.200 ;
        RECT 0.270 617.120 199.575 621.840 ;
        RECT 4.400 615.720 199.575 617.120 ;
        RECT 0.270 612.360 199.575 615.720 ;
        RECT 0.270 610.960 195.600 612.360 ;
        RECT 0.270 609.640 199.575 610.960 ;
        RECT 4.400 608.240 199.575 609.640 ;
        RECT 0.270 602.160 199.575 608.240 ;
        RECT 4.400 601.480 199.575 602.160 ;
        RECT 4.400 600.760 195.600 601.480 ;
        RECT 0.270 600.080 195.600 600.760 ;
        RECT 0.270 594.680 199.575 600.080 ;
        RECT 4.400 593.280 199.575 594.680 ;
        RECT 0.270 590.600 199.575 593.280 ;
        RECT 0.270 589.200 195.600 590.600 ;
        RECT 0.270 587.200 199.575 589.200 ;
        RECT 4.400 585.800 199.575 587.200 ;
        RECT 0.270 579.720 199.575 585.800 ;
        RECT 4.400 578.320 195.600 579.720 ;
        RECT 0.270 572.240 199.575 578.320 ;
        RECT 4.400 570.840 199.575 572.240 ;
        RECT 0.270 568.840 199.575 570.840 ;
        RECT 0.270 567.440 195.600 568.840 ;
        RECT 0.270 564.760 199.575 567.440 ;
        RECT 4.400 563.360 199.575 564.760 ;
        RECT 0.270 557.960 199.575 563.360 ;
        RECT 0.270 557.280 195.600 557.960 ;
        RECT 4.400 556.560 195.600 557.280 ;
        RECT 4.400 555.880 199.575 556.560 ;
        RECT 0.270 549.800 199.575 555.880 ;
        RECT 4.400 548.400 199.575 549.800 ;
        RECT 0.270 547.080 199.575 548.400 ;
        RECT 0.270 545.680 195.600 547.080 ;
        RECT 0.270 542.320 199.575 545.680 ;
        RECT 4.400 540.920 199.575 542.320 ;
        RECT 0.270 536.200 199.575 540.920 ;
        RECT 0.270 534.840 195.600 536.200 ;
        RECT 4.400 534.800 195.600 534.840 ;
        RECT 4.400 533.440 199.575 534.800 ;
        RECT 0.270 527.360 199.575 533.440 ;
        RECT 4.400 525.960 199.575 527.360 ;
        RECT 0.270 525.320 199.575 525.960 ;
        RECT 0.270 523.920 195.600 525.320 ;
        RECT 0.270 519.880 199.575 523.920 ;
        RECT 4.400 518.480 199.575 519.880 ;
        RECT 0.270 514.440 199.575 518.480 ;
        RECT 0.270 513.040 195.600 514.440 ;
        RECT 0.270 512.400 199.575 513.040 ;
        RECT 4.400 511.000 199.575 512.400 ;
        RECT 0.270 504.920 199.575 511.000 ;
        RECT 4.400 503.560 199.575 504.920 ;
        RECT 4.400 503.520 195.600 503.560 ;
        RECT 0.270 502.160 195.600 503.520 ;
        RECT 0.270 497.440 199.575 502.160 ;
        RECT 4.400 496.040 199.575 497.440 ;
        RECT 0.270 492.680 199.575 496.040 ;
        RECT 0.270 491.280 195.600 492.680 ;
        RECT 0.270 489.960 199.575 491.280 ;
        RECT 4.400 488.560 199.575 489.960 ;
        RECT 0.270 482.480 199.575 488.560 ;
        RECT 4.400 481.800 199.575 482.480 ;
        RECT 4.400 481.080 195.600 481.800 ;
        RECT 0.270 480.400 195.600 481.080 ;
        RECT 0.270 475.000 199.575 480.400 ;
        RECT 4.400 473.600 199.575 475.000 ;
        RECT 0.270 470.920 199.575 473.600 ;
        RECT 0.270 469.520 195.600 470.920 ;
        RECT 0.270 467.520 199.575 469.520 ;
        RECT 4.400 466.120 199.575 467.520 ;
        RECT 0.270 460.040 199.575 466.120 ;
        RECT 4.400 458.640 195.600 460.040 ;
        RECT 0.270 452.560 199.575 458.640 ;
        RECT 4.400 451.160 199.575 452.560 ;
        RECT 0.270 449.160 199.575 451.160 ;
        RECT 0.270 447.760 195.600 449.160 ;
        RECT 0.270 445.080 199.575 447.760 ;
        RECT 4.400 443.680 199.575 445.080 ;
        RECT 0.270 438.280 199.575 443.680 ;
        RECT 0.270 437.600 195.600 438.280 ;
        RECT 4.400 436.880 195.600 437.600 ;
        RECT 4.400 436.200 199.575 436.880 ;
        RECT 0.270 430.120 199.575 436.200 ;
        RECT 4.400 428.720 199.575 430.120 ;
        RECT 0.270 427.400 199.575 428.720 ;
        RECT 0.270 426.000 195.600 427.400 ;
        RECT 0.270 422.640 199.575 426.000 ;
        RECT 4.400 421.240 199.575 422.640 ;
        RECT 0.270 416.520 199.575 421.240 ;
        RECT 0.270 415.160 195.600 416.520 ;
        RECT 4.400 415.120 195.600 415.160 ;
        RECT 4.400 413.760 199.575 415.120 ;
        RECT 0.270 407.680 199.575 413.760 ;
        RECT 4.400 406.280 199.575 407.680 ;
        RECT 0.270 405.640 199.575 406.280 ;
        RECT 0.270 404.240 195.600 405.640 ;
        RECT 0.270 400.200 199.575 404.240 ;
        RECT 4.400 398.800 199.575 400.200 ;
        RECT 0.270 394.760 199.575 398.800 ;
        RECT 0.270 393.360 195.600 394.760 ;
        RECT 0.270 392.720 199.575 393.360 ;
        RECT 4.400 391.320 199.575 392.720 ;
        RECT 0.270 385.240 199.575 391.320 ;
        RECT 4.400 383.880 199.575 385.240 ;
        RECT 4.400 383.840 195.600 383.880 ;
        RECT 0.270 382.480 195.600 383.840 ;
        RECT 0.270 377.760 199.575 382.480 ;
        RECT 4.400 376.360 199.575 377.760 ;
        RECT 0.270 373.000 199.575 376.360 ;
        RECT 0.270 371.600 195.600 373.000 ;
        RECT 0.270 370.280 199.575 371.600 ;
        RECT 4.400 368.880 199.575 370.280 ;
        RECT 0.270 362.800 199.575 368.880 ;
        RECT 4.400 362.120 199.575 362.800 ;
        RECT 4.400 361.400 195.600 362.120 ;
        RECT 0.270 360.720 195.600 361.400 ;
        RECT 0.270 355.320 199.575 360.720 ;
        RECT 4.400 353.920 199.575 355.320 ;
        RECT 0.270 351.240 199.575 353.920 ;
        RECT 0.270 349.840 195.600 351.240 ;
        RECT 0.270 347.840 199.575 349.840 ;
        RECT 4.400 346.440 199.575 347.840 ;
        RECT 0.270 340.360 199.575 346.440 ;
        RECT 4.400 338.960 195.600 340.360 ;
        RECT 0.270 332.880 199.575 338.960 ;
        RECT 4.400 331.480 199.575 332.880 ;
        RECT 0.270 329.480 199.575 331.480 ;
        RECT 0.270 328.080 195.600 329.480 ;
        RECT 0.270 325.400 199.575 328.080 ;
        RECT 4.400 324.000 199.575 325.400 ;
        RECT 0.270 318.600 199.575 324.000 ;
        RECT 0.270 317.920 195.600 318.600 ;
        RECT 4.400 317.200 195.600 317.920 ;
        RECT 4.400 316.520 199.575 317.200 ;
        RECT 0.270 310.440 199.575 316.520 ;
        RECT 4.400 309.040 199.575 310.440 ;
        RECT 0.270 307.720 199.575 309.040 ;
        RECT 0.270 306.320 195.600 307.720 ;
        RECT 0.270 302.960 199.575 306.320 ;
        RECT 4.400 301.560 199.575 302.960 ;
        RECT 0.270 296.840 199.575 301.560 ;
        RECT 0.270 295.480 195.600 296.840 ;
        RECT 4.400 295.440 195.600 295.480 ;
        RECT 4.400 294.080 199.575 295.440 ;
        RECT 0.270 288.000 199.575 294.080 ;
        RECT 4.400 286.600 199.575 288.000 ;
        RECT 0.270 285.960 199.575 286.600 ;
        RECT 0.270 284.560 195.600 285.960 ;
        RECT 0.270 280.520 199.575 284.560 ;
        RECT 4.400 279.120 199.575 280.520 ;
        RECT 0.270 275.080 199.575 279.120 ;
        RECT 0.270 273.680 195.600 275.080 ;
        RECT 0.270 273.040 199.575 273.680 ;
        RECT 4.400 271.640 199.575 273.040 ;
        RECT 0.270 265.560 199.575 271.640 ;
        RECT 4.400 264.200 199.575 265.560 ;
        RECT 4.400 264.160 195.600 264.200 ;
        RECT 0.270 262.800 195.600 264.160 ;
        RECT 0.270 258.080 199.575 262.800 ;
        RECT 4.400 256.680 199.575 258.080 ;
        RECT 0.270 253.320 199.575 256.680 ;
        RECT 0.270 251.920 195.600 253.320 ;
        RECT 0.270 250.600 199.575 251.920 ;
        RECT 4.400 249.200 199.575 250.600 ;
        RECT 0.270 243.120 199.575 249.200 ;
        RECT 4.400 242.440 199.575 243.120 ;
        RECT 4.400 241.720 195.600 242.440 ;
        RECT 0.270 241.040 195.600 241.720 ;
        RECT 0.270 235.640 199.575 241.040 ;
        RECT 4.400 234.240 199.575 235.640 ;
        RECT 0.270 231.560 199.575 234.240 ;
        RECT 0.270 230.160 195.600 231.560 ;
        RECT 0.270 228.160 199.575 230.160 ;
        RECT 4.400 226.760 199.575 228.160 ;
        RECT 0.270 220.680 199.575 226.760 ;
        RECT 4.400 219.280 195.600 220.680 ;
        RECT 0.270 213.200 199.575 219.280 ;
        RECT 4.400 211.800 199.575 213.200 ;
        RECT 0.270 209.800 199.575 211.800 ;
        RECT 0.270 208.400 195.600 209.800 ;
        RECT 0.270 205.720 199.575 208.400 ;
        RECT 4.400 204.320 199.575 205.720 ;
        RECT 0.270 198.920 199.575 204.320 ;
        RECT 0.270 198.240 195.600 198.920 ;
        RECT 4.400 197.520 195.600 198.240 ;
        RECT 4.400 196.840 199.575 197.520 ;
        RECT 0.270 190.760 199.575 196.840 ;
        RECT 4.400 189.360 199.575 190.760 ;
        RECT 0.270 188.040 199.575 189.360 ;
        RECT 0.270 186.640 195.600 188.040 ;
        RECT 0.270 183.280 199.575 186.640 ;
        RECT 4.400 181.880 199.575 183.280 ;
        RECT 0.270 177.160 199.575 181.880 ;
        RECT 0.270 175.800 195.600 177.160 ;
        RECT 4.400 175.760 195.600 175.800 ;
        RECT 4.400 174.400 199.575 175.760 ;
        RECT 0.270 168.320 199.575 174.400 ;
        RECT 4.400 166.920 199.575 168.320 ;
        RECT 0.270 166.280 199.575 166.920 ;
        RECT 0.270 164.880 195.600 166.280 ;
        RECT 0.270 160.840 199.575 164.880 ;
        RECT 4.400 159.440 199.575 160.840 ;
        RECT 0.270 155.400 199.575 159.440 ;
        RECT 0.270 154.000 195.600 155.400 ;
        RECT 0.270 153.360 199.575 154.000 ;
        RECT 4.400 151.960 199.575 153.360 ;
        RECT 0.270 145.880 199.575 151.960 ;
        RECT 4.400 144.520 199.575 145.880 ;
        RECT 4.400 144.480 195.600 144.520 ;
        RECT 0.270 143.120 195.600 144.480 ;
        RECT 0.270 138.400 199.575 143.120 ;
        RECT 4.400 137.000 199.575 138.400 ;
        RECT 0.270 133.640 199.575 137.000 ;
        RECT 0.270 132.240 195.600 133.640 ;
        RECT 0.270 130.920 199.575 132.240 ;
        RECT 4.400 129.520 199.575 130.920 ;
        RECT 0.270 123.440 199.575 129.520 ;
        RECT 4.400 122.760 199.575 123.440 ;
        RECT 4.400 122.040 195.600 122.760 ;
        RECT 0.270 121.360 195.600 122.040 ;
        RECT 0.270 115.960 199.575 121.360 ;
        RECT 4.400 114.560 199.575 115.960 ;
        RECT 0.270 111.880 199.575 114.560 ;
        RECT 0.270 110.480 195.600 111.880 ;
        RECT 0.270 108.480 199.575 110.480 ;
        RECT 4.400 107.080 199.575 108.480 ;
        RECT 0.270 101.000 199.575 107.080 ;
        RECT 4.400 99.600 195.600 101.000 ;
        RECT 0.270 93.520 199.575 99.600 ;
        RECT 4.400 92.120 199.575 93.520 ;
        RECT 0.270 90.120 199.575 92.120 ;
        RECT 0.270 88.720 195.600 90.120 ;
        RECT 0.270 86.040 199.575 88.720 ;
        RECT 4.400 84.640 199.575 86.040 ;
        RECT 0.270 79.240 199.575 84.640 ;
        RECT 0.270 78.560 195.600 79.240 ;
        RECT 4.400 77.840 195.600 78.560 ;
        RECT 4.400 77.160 199.575 77.840 ;
        RECT 0.270 71.080 199.575 77.160 ;
        RECT 4.400 69.680 199.575 71.080 ;
        RECT 0.270 68.360 199.575 69.680 ;
        RECT 0.270 66.960 195.600 68.360 ;
        RECT 0.270 63.600 199.575 66.960 ;
        RECT 4.400 62.200 199.575 63.600 ;
        RECT 0.270 57.480 199.575 62.200 ;
        RECT 0.270 56.120 195.600 57.480 ;
        RECT 4.400 56.080 195.600 56.120 ;
        RECT 4.400 54.720 199.575 56.080 ;
        RECT 0.270 48.640 199.575 54.720 ;
        RECT 4.400 47.240 199.575 48.640 ;
        RECT 0.270 46.600 199.575 47.240 ;
        RECT 0.270 45.200 195.600 46.600 ;
        RECT 0.270 41.160 199.575 45.200 ;
        RECT 4.400 39.760 199.575 41.160 ;
        RECT 0.270 35.720 199.575 39.760 ;
        RECT 0.270 34.320 195.600 35.720 ;
        RECT 0.270 33.680 199.575 34.320 ;
        RECT 4.400 32.280 199.575 33.680 ;
        RECT 0.270 26.200 199.575 32.280 ;
        RECT 4.400 24.840 199.575 26.200 ;
        RECT 4.400 24.800 195.600 24.840 ;
        RECT 0.270 23.440 195.600 24.800 ;
        RECT 0.270 18.720 199.575 23.440 ;
        RECT 4.400 17.320 199.575 18.720 ;
        RECT 0.270 13.960 199.575 17.320 ;
        RECT 0.270 12.560 195.600 13.960 ;
        RECT 0.270 11.240 199.575 12.560 ;
        RECT 4.400 10.375 199.575 11.240 ;
      LAYER met4 ;
        RECT 0.295 12.415 20.640 787.945 ;
        RECT 23.040 12.415 97.440 787.945 ;
        RECT 99.840 12.415 174.240 787.945 ;
        RECT 176.640 12.415 185.545 787.945 ;
  END
END core
END LIBRARY

