magic
tech sky130B
magscale 1 2
timestamp 1662672245
<< obsli1 >>
rect 1104 2159 161368 162129
<< obsm1 >>
rect 14 1708 161722 162580
<< metal2 >>
rect 2594 163845 2650 164645
rect 5814 163845 5870 164645
rect 9678 163845 9734 164645
rect 13542 163845 13598 164645
rect 16762 163845 16818 164645
rect 20626 163845 20682 164645
rect 24490 163845 24546 164645
rect 28354 163845 28410 164645
rect 31574 163845 31630 164645
rect 35438 163845 35494 164645
rect 39302 163845 39358 164645
rect 43166 163845 43222 164645
rect 46386 163845 46442 164645
rect 50250 163845 50306 164645
rect 54114 163845 54170 164645
rect 57334 163845 57390 164645
rect 61198 163845 61254 164645
rect 65062 163845 65118 164645
rect 68926 163845 68982 164645
rect 72146 163845 72202 164645
rect 76010 163845 76066 164645
rect 79874 163845 79930 164645
rect 83094 163845 83150 164645
rect 86958 163845 87014 164645
rect 90822 163845 90878 164645
rect 94686 163845 94742 164645
rect 97906 163845 97962 164645
rect 101770 163845 101826 164645
rect 105634 163845 105690 164645
rect 109498 163845 109554 164645
rect 112718 163845 112774 164645
rect 116582 163845 116638 164645
rect 120446 163845 120502 164645
rect 123666 163845 123722 164645
rect 127530 163845 127586 164645
rect 131394 163845 131450 164645
rect 135258 163845 135314 164645
rect 138478 163845 138534 164645
rect 142342 163845 142398 164645
rect 146206 163845 146262 164645
rect 149426 163845 149482 164645
rect 153290 163845 153346 164645
rect 157154 163845 157210 164645
rect 161018 163845 161074 164645
rect 18 0 74 800
rect 3238 0 3294 800
rect 7102 0 7158 800
rect 10966 0 11022 800
rect 14186 0 14242 800
rect 18050 0 18106 800
rect 21914 0 21970 800
rect 25778 0 25834 800
rect 28998 0 29054 800
rect 32862 0 32918 800
rect 36726 0 36782 800
rect 39946 0 40002 800
rect 43810 0 43866 800
rect 47674 0 47730 800
rect 51538 0 51594 800
rect 54758 0 54814 800
rect 58622 0 58678 800
rect 62486 0 62542 800
rect 66350 0 66406 800
rect 69570 0 69626 800
rect 73434 0 73490 800
rect 77298 0 77354 800
rect 80518 0 80574 800
rect 84382 0 84438 800
rect 88246 0 88302 800
rect 92110 0 92166 800
rect 95330 0 95386 800
rect 99194 0 99250 800
rect 103058 0 103114 800
rect 106278 0 106334 800
rect 110142 0 110198 800
rect 114006 0 114062 800
rect 117870 0 117926 800
rect 121090 0 121146 800
rect 124954 0 125010 800
rect 128818 0 128874 800
rect 132682 0 132738 800
rect 135902 0 135958 800
rect 139766 0 139822 800
rect 143630 0 143686 800
rect 146850 0 146906 800
rect 150714 0 150770 800
rect 154578 0 154634 800
rect 158442 0 158498 800
rect 161662 0 161718 800
<< obsm2 >>
rect 20 163789 2538 163962
rect 2706 163789 5758 163962
rect 5926 163789 9622 163962
rect 9790 163789 13486 163962
rect 13654 163789 16706 163962
rect 16874 163789 20570 163962
rect 20738 163789 24434 163962
rect 24602 163789 28298 163962
rect 28466 163789 31518 163962
rect 31686 163789 35382 163962
rect 35550 163789 39246 163962
rect 39414 163789 43110 163962
rect 43278 163789 46330 163962
rect 46498 163789 50194 163962
rect 50362 163789 54058 163962
rect 54226 163789 57278 163962
rect 57446 163789 61142 163962
rect 61310 163789 65006 163962
rect 65174 163789 68870 163962
rect 69038 163789 72090 163962
rect 72258 163789 75954 163962
rect 76122 163789 79818 163962
rect 79986 163789 83038 163962
rect 83206 163789 86902 163962
rect 87070 163789 90766 163962
rect 90934 163789 94630 163962
rect 94798 163789 97850 163962
rect 98018 163789 101714 163962
rect 101882 163789 105578 163962
rect 105746 163789 109442 163962
rect 109610 163789 112662 163962
rect 112830 163789 116526 163962
rect 116694 163789 120390 163962
rect 120558 163789 123610 163962
rect 123778 163789 127474 163962
rect 127642 163789 131338 163962
rect 131506 163789 135202 163962
rect 135370 163789 138422 163962
rect 138590 163789 142286 163962
rect 142454 163789 146150 163962
rect 146318 163789 149370 163962
rect 149538 163789 153234 163962
rect 153402 163789 157098 163962
rect 157266 163789 160962 163962
rect 161130 163789 161716 163962
rect 20 856 161716 163789
rect 130 734 3182 856
rect 3350 734 7046 856
rect 7214 734 10910 856
rect 11078 734 14130 856
rect 14298 734 17994 856
rect 18162 734 21858 856
rect 22026 734 25722 856
rect 25890 734 28942 856
rect 29110 734 32806 856
rect 32974 734 36670 856
rect 36838 734 39890 856
rect 40058 734 43754 856
rect 43922 734 47618 856
rect 47786 734 51482 856
rect 51650 734 54702 856
rect 54870 734 58566 856
rect 58734 734 62430 856
rect 62598 734 66294 856
rect 66462 734 69514 856
rect 69682 734 73378 856
rect 73546 734 77242 856
rect 77410 734 80462 856
rect 80630 734 84326 856
rect 84494 734 88190 856
rect 88358 734 92054 856
rect 92222 734 95274 856
rect 95442 734 99138 856
rect 99306 734 103002 856
rect 103170 734 106222 856
rect 106390 734 110086 856
rect 110254 734 113950 856
rect 114118 734 117814 856
rect 117982 734 121034 856
rect 121202 734 124898 856
rect 125066 734 128762 856
rect 128930 734 132626 856
rect 132794 734 135846 856
rect 136014 734 139710 856
rect 139878 734 143574 856
rect 143742 734 146794 856
rect 146962 734 150658 856
rect 150826 734 154522 856
rect 154690 734 158386 856
rect 158554 734 161606 856
<< metal3 >>
rect 0 163208 800 163328
rect 161701 162528 162501 162648
rect 0 159128 800 159248
rect 161701 158448 162501 158568
rect 0 155048 800 155168
rect 161701 154368 162501 154488
rect 0 151648 800 151768
rect 161701 150288 162501 150408
rect 0 147568 800 147688
rect 161701 146888 162501 147008
rect 0 143488 800 143608
rect 161701 142808 162501 142928
rect 0 140088 800 140208
rect 161701 138728 162501 138848
rect 0 136008 800 136128
rect 161701 135328 162501 135448
rect 0 131928 800 132048
rect 161701 131248 162501 131368
rect 0 127848 800 127968
rect 161701 127168 162501 127288
rect 0 124448 800 124568
rect 161701 123088 162501 123208
rect 0 120368 800 120488
rect 161701 119688 162501 119808
rect 0 116288 800 116408
rect 161701 115608 162501 115728
rect 0 112208 800 112328
rect 161701 111528 162501 111648
rect 0 108808 800 108928
rect 161701 108128 162501 108248
rect 0 104728 800 104848
rect 161701 104048 162501 104168
rect 0 100648 800 100768
rect 161701 99968 162501 100088
rect 0 97248 800 97368
rect 161701 95888 162501 96008
rect 0 93168 800 93288
rect 161701 92488 162501 92608
rect 0 89088 800 89208
rect 161701 88408 162501 88528
rect 0 85008 800 85128
rect 161701 84328 162501 84448
rect 0 81608 800 81728
rect 161701 80248 162501 80368
rect 0 77528 800 77648
rect 161701 76848 162501 76968
rect 0 73448 800 73568
rect 161701 72768 162501 72888
rect 0 70048 800 70168
rect 161701 68688 162501 68808
rect 0 65968 800 66088
rect 161701 65288 162501 65408
rect 0 61888 800 62008
rect 161701 61208 162501 61328
rect 0 57808 800 57928
rect 161701 57128 162501 57248
rect 0 54408 800 54528
rect 161701 53048 162501 53168
rect 0 50328 800 50448
rect 161701 49648 162501 49768
rect 0 46248 800 46368
rect 161701 45568 162501 45688
rect 0 42168 800 42288
rect 161701 41488 162501 41608
rect 0 38768 800 38888
rect 161701 38088 162501 38208
rect 0 34688 800 34808
rect 161701 34008 162501 34128
rect 0 30608 800 30728
rect 161701 29928 162501 30048
rect 0 27208 800 27328
rect 161701 25848 162501 25968
rect 0 23128 800 23248
rect 161701 22448 162501 22568
rect 0 19048 800 19168
rect 161701 18368 162501 18488
rect 0 14968 800 15088
rect 161701 14288 162501 14408
rect 0 11568 800 11688
rect 161701 10208 162501 10328
rect 0 7488 800 7608
rect 161701 6808 162501 6928
rect 0 3408 800 3528
rect 161701 2728 162501 2848
<< obsm3 >>
rect 880 163128 161701 163301
rect 800 162728 161701 163128
rect 800 162448 161621 162728
rect 800 159328 161701 162448
rect 880 159048 161701 159328
rect 800 158648 161701 159048
rect 800 158368 161621 158648
rect 800 155248 161701 158368
rect 880 154968 161701 155248
rect 800 154568 161701 154968
rect 800 154288 161621 154568
rect 800 151848 161701 154288
rect 880 151568 161701 151848
rect 800 150488 161701 151568
rect 800 150208 161621 150488
rect 800 147768 161701 150208
rect 880 147488 161701 147768
rect 800 147088 161701 147488
rect 800 146808 161621 147088
rect 800 143688 161701 146808
rect 880 143408 161701 143688
rect 800 143008 161701 143408
rect 800 142728 161621 143008
rect 800 140288 161701 142728
rect 880 140008 161701 140288
rect 800 138928 161701 140008
rect 800 138648 161621 138928
rect 800 136208 161701 138648
rect 880 135928 161701 136208
rect 800 135528 161701 135928
rect 800 135248 161621 135528
rect 800 132128 161701 135248
rect 880 131848 161701 132128
rect 800 131448 161701 131848
rect 800 131168 161621 131448
rect 800 128048 161701 131168
rect 880 127768 161701 128048
rect 800 127368 161701 127768
rect 800 127088 161621 127368
rect 800 124648 161701 127088
rect 880 124368 161701 124648
rect 800 123288 161701 124368
rect 800 123008 161621 123288
rect 800 120568 161701 123008
rect 880 120288 161701 120568
rect 800 119888 161701 120288
rect 800 119608 161621 119888
rect 800 116488 161701 119608
rect 880 116208 161701 116488
rect 800 115808 161701 116208
rect 800 115528 161621 115808
rect 800 112408 161701 115528
rect 880 112128 161701 112408
rect 800 111728 161701 112128
rect 800 111448 161621 111728
rect 800 109008 161701 111448
rect 880 108728 161701 109008
rect 800 108328 161701 108728
rect 800 108048 161621 108328
rect 800 104928 161701 108048
rect 880 104648 161701 104928
rect 800 104248 161701 104648
rect 800 103968 161621 104248
rect 800 100848 161701 103968
rect 880 100568 161701 100848
rect 800 100168 161701 100568
rect 800 99888 161621 100168
rect 800 97448 161701 99888
rect 880 97168 161701 97448
rect 800 96088 161701 97168
rect 800 95808 161621 96088
rect 800 93368 161701 95808
rect 880 93088 161701 93368
rect 800 92688 161701 93088
rect 800 92408 161621 92688
rect 800 89288 161701 92408
rect 880 89008 161701 89288
rect 800 88608 161701 89008
rect 800 88328 161621 88608
rect 800 85208 161701 88328
rect 880 84928 161701 85208
rect 800 84528 161701 84928
rect 800 84248 161621 84528
rect 800 81808 161701 84248
rect 880 81528 161701 81808
rect 800 80448 161701 81528
rect 800 80168 161621 80448
rect 800 77728 161701 80168
rect 880 77448 161701 77728
rect 800 77048 161701 77448
rect 800 76768 161621 77048
rect 800 73648 161701 76768
rect 880 73368 161701 73648
rect 800 72968 161701 73368
rect 800 72688 161621 72968
rect 800 70248 161701 72688
rect 880 69968 161701 70248
rect 800 68888 161701 69968
rect 800 68608 161621 68888
rect 800 66168 161701 68608
rect 880 65888 161701 66168
rect 800 65488 161701 65888
rect 800 65208 161621 65488
rect 800 62088 161701 65208
rect 880 61808 161701 62088
rect 800 61408 161701 61808
rect 800 61128 161621 61408
rect 800 58008 161701 61128
rect 880 57728 161701 58008
rect 800 57328 161701 57728
rect 800 57048 161621 57328
rect 800 54608 161701 57048
rect 880 54328 161701 54608
rect 800 53248 161701 54328
rect 800 52968 161621 53248
rect 800 50528 161701 52968
rect 880 50248 161701 50528
rect 800 49848 161701 50248
rect 800 49568 161621 49848
rect 800 46448 161701 49568
rect 880 46168 161701 46448
rect 800 45768 161701 46168
rect 800 45488 161621 45768
rect 800 42368 161701 45488
rect 880 42088 161701 42368
rect 800 41688 161701 42088
rect 800 41408 161621 41688
rect 800 38968 161701 41408
rect 880 38688 161701 38968
rect 800 38288 161701 38688
rect 800 38008 161621 38288
rect 800 34888 161701 38008
rect 880 34608 161701 34888
rect 800 34208 161701 34608
rect 800 33928 161621 34208
rect 800 30808 161701 33928
rect 880 30528 161701 30808
rect 800 30128 161701 30528
rect 800 29848 161621 30128
rect 800 27408 161701 29848
rect 880 27128 161701 27408
rect 800 26048 161701 27128
rect 800 25768 161621 26048
rect 800 23328 161701 25768
rect 880 23048 161701 23328
rect 800 22648 161701 23048
rect 800 22368 161621 22648
rect 800 19248 161701 22368
rect 880 18968 161701 19248
rect 800 18568 161701 18968
rect 800 18288 161621 18568
rect 800 15168 161701 18288
rect 880 14888 161701 15168
rect 800 14488 161701 14888
rect 800 14208 161621 14488
rect 800 11768 161701 14208
rect 880 11488 161701 11768
rect 800 10408 161701 11488
rect 800 10128 161621 10408
rect 800 7688 161701 10128
rect 880 7408 161701 7688
rect 800 7008 161701 7408
rect 800 6728 161621 7008
rect 800 3608 161701 6728
rect 880 3328 161701 3608
rect 800 2928 161701 3328
rect 800 2648 161621 2928
rect 800 1939 161701 2648
<< metal4 >>
rect 4208 2128 4528 162160
rect 19568 2128 19888 162160
rect 34928 2128 35248 162160
rect 50288 2128 50608 162160
rect 65648 2128 65968 162160
rect 81008 2128 81328 162160
rect 96368 2128 96688 162160
rect 111728 2128 112048 162160
rect 127088 2128 127408 162160
rect 142448 2128 142768 162160
rect 157808 2128 158128 162160
<< obsm4 >>
rect 1715 162240 159653 162485
rect 1715 2048 4128 162240
rect 4608 2048 19488 162240
rect 19968 2048 34848 162240
rect 35328 2048 50208 162240
rect 50688 2048 65568 162240
rect 66048 2048 80928 162240
rect 81408 2048 96288 162240
rect 96768 2048 111648 162240
rect 112128 2048 127008 162240
rect 127488 2048 142368 162240
rect 142848 2048 157728 162240
rect 158208 2048 159653 162240
rect 1715 1939 159653 2048
<< metal5 >>
rect 1056 158526 161416 158846
rect 1056 143208 161416 143528
rect 1056 127890 161416 128210
rect 1056 112572 161416 112892
rect 1056 97254 161416 97574
rect 1056 81936 161416 82256
rect 1056 66618 161416 66938
rect 1056 51300 161416 51620
rect 1056 35982 161416 36302
rect 1056 20664 161416 20984
rect 1056 5346 161416 5666
<< labels >>
rlabel metal4 s 19568 2128 19888 162160 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 162160 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 162160 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 162160 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 162160 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 20664 161416 20984 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 51300 161416 51620 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 81936 161416 82256 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 112572 161416 112892 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 143208 161416 143528 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 162160 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 162160 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 162160 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 162160 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 162160 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 162160 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5346 161416 5666 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 35982 161416 36302 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 66618 161416 66938 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 97254 161416 97574 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 127890 161416 128210 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 158526 161416 158846 6 VPWR
port 2 nsew power bidirectional
rlabel metal2 s 157154 163845 157210 164645 6 i_addr[0]
port 3 nsew signal input
rlabel metal2 s 65062 163845 65118 164645 6 i_addr[1]
port 4 nsew signal input
rlabel metal3 s 161701 22448 162501 22568 6 i_addr[2]
port 5 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 i_addr[3]
port 6 nsew signal input
rlabel metal3 s 0 131928 800 132048 6 i_addr[4]
port 7 nsew signal input
rlabel metal2 s 20626 163845 20682 164645 6 i_addr[5]
port 8 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 i_clk
port 9 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 i_data[0]
port 10 nsew signal input
rlabel metal2 s 132682 0 132738 800 6 i_data[10]
port 11 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 i_data[11]
port 12 nsew signal input
rlabel metal3 s 161701 154368 162501 154488 6 i_data[12]
port 13 nsew signal input
rlabel metal2 s 105634 163845 105690 164645 6 i_data[13]
port 14 nsew signal input
rlabel metal2 s 97906 163845 97962 164645 6 i_data[14]
port 15 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 i_data[15]
port 16 nsew signal input
rlabel metal2 s 76010 163845 76066 164645 6 i_data[16]
port 17 nsew signal input
rlabel metal2 s 36726 0 36782 800 6 i_data[17]
port 18 nsew signal input
rlabel metal2 s 13542 163845 13598 164645 6 i_data[18]
port 19 nsew signal input
rlabel metal3 s 0 163208 800 163328 6 i_data[19]
port 20 nsew signal input
rlabel metal2 s 94686 163845 94742 164645 6 i_data[1]
port 21 nsew signal input
rlabel metal3 s 161701 25848 162501 25968 6 i_data[20]
port 22 nsew signal input
rlabel metal2 s 35438 163845 35494 164645 6 i_data[21]
port 23 nsew signal input
rlabel metal2 s 72146 163845 72202 164645 6 i_data[22]
port 24 nsew signal input
rlabel metal3 s 161701 72768 162501 72888 6 i_data[23]
port 25 nsew signal input
rlabel metal2 s 39302 163845 39358 164645 6 i_data[24]
port 26 nsew signal input
rlabel metal3 s 161701 146888 162501 147008 6 i_data[25]
port 27 nsew signal input
rlabel metal3 s 161701 14288 162501 14408 6 i_data[26]
port 28 nsew signal input
rlabel metal2 s 123666 163845 123722 164645 6 i_data[27]
port 29 nsew signal input
rlabel metal3 s 161701 10208 162501 10328 6 i_data[28]
port 30 nsew signal input
rlabel metal2 s 128818 0 128874 800 6 i_data[29]
port 31 nsew signal input
rlabel metal3 s 0 85008 800 85128 6 i_data[2]
port 32 nsew signal input
rlabel metal2 s 9678 163845 9734 164645 6 i_data[30]
port 33 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 i_data[31]
port 34 nsew signal input
rlabel metal3 s 161701 138728 162501 138848 6 i_data[32]
port 35 nsew signal input
rlabel metal2 s 51538 0 51594 800 6 i_data[33]
port 36 nsew signal input
rlabel metal2 s 31574 163845 31630 164645 6 i_data[34]
port 37 nsew signal input
rlabel metal3 s 0 57808 800 57928 6 i_data[35]
port 38 nsew signal input
rlabel metal2 s 146206 163845 146262 164645 6 i_data[36]
port 39 nsew signal input
rlabel metal2 s 5814 163845 5870 164645 6 i_data[37]
port 40 nsew signal input
rlabel metal2 s 50250 163845 50306 164645 6 i_data[38]
port 41 nsew signal input
rlabel metal3 s 161701 131248 162501 131368 6 i_data[39]
port 42 nsew signal input
rlabel metal3 s 161701 104048 162501 104168 6 i_data[3]
port 43 nsew signal input
rlabel metal3 s 161701 68688 162501 68808 6 i_data[40]
port 44 nsew signal input
rlabel metal2 s 131394 163845 131450 164645 6 i_data[41]
port 45 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 i_data[42]
port 46 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 i_data[43]
port 47 nsew signal input
rlabel metal2 s 161662 0 161718 800 6 i_data[44]
port 48 nsew signal input
rlabel metal3 s 161701 127168 162501 127288 6 i_data[45]
port 49 nsew signal input
rlabel metal2 s 103058 0 103114 800 6 i_data[46]
port 50 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 i_data[47]
port 51 nsew signal input
rlabel metal3 s 161701 88408 162501 88528 6 i_data[48]
port 52 nsew signal input
rlabel metal2 s 153290 163845 153346 164645 6 i_data[49]
port 53 nsew signal input
rlabel metal2 s 68926 163845 68982 164645 6 i_data[4]
port 54 nsew signal input
rlabel metal3 s 161701 80248 162501 80368 6 i_data[50]
port 55 nsew signal input
rlabel metal2 s 149426 163845 149482 164645 6 i_data[51]
port 56 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 i_data[52]
port 57 nsew signal input
rlabel metal3 s 161701 34008 162501 34128 6 i_data[53]
port 58 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 i_data[54]
port 59 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 i_data[55]
port 60 nsew signal input
rlabel metal2 s 142342 163845 142398 164645 6 i_data[56]
port 61 nsew signal input
rlabel metal3 s 161701 162528 162501 162648 6 i_data[57]
port 62 nsew signal input
rlabel metal2 s 61198 163845 61254 164645 6 i_data[58]
port 63 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 i_data[59]
port 64 nsew signal input
rlabel metal2 s 101770 163845 101826 164645 6 i_data[5]
port 65 nsew signal input
rlabel metal2 s 16762 163845 16818 164645 6 i_data[60]
port 66 nsew signal input
rlabel metal2 s 139766 0 139822 800 6 i_data[61]
port 67 nsew signal input
rlabel metal3 s 0 159128 800 159248 6 i_data[62]
port 68 nsew signal input
rlabel metal3 s 0 143488 800 143608 6 i_data[63]
port 69 nsew signal input
rlabel metal3 s 0 116288 800 116408 6 i_data[64]
port 70 nsew signal input
rlabel metal2 s 138478 163845 138534 164645 6 i_data[65]
port 71 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 i_data[66]
port 72 nsew signal input
rlabel metal3 s 161701 41488 162501 41608 6 i_data[67]
port 73 nsew signal input
rlabel metal3 s 161701 61208 162501 61328 6 i_data[68]
port 74 nsew signal input
rlabel metal3 s 0 155048 800 155168 6 i_data[69]
port 75 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 i_data[6]
port 76 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 i_data[70]
port 77 nsew signal input
rlabel metal2 s 158442 0 158498 800 6 i_data[71]
port 78 nsew signal input
rlabel metal3 s 0 127848 800 127968 6 i_data[72]
port 79 nsew signal input
rlabel metal3 s 0 46248 800 46368 6 i_data[73]
port 80 nsew signal input
rlabel metal3 s 0 65968 800 66088 6 i_data[74]
port 81 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 i_data[75]
port 82 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 i_data[76]
port 83 nsew signal input
rlabel metal2 s 46386 163845 46442 164645 6 i_data[77]
port 84 nsew signal input
rlabel metal2 s 57334 163845 57390 164645 6 i_data[78]
port 85 nsew signal input
rlabel metal3 s 0 124448 800 124568 6 i_data[79]
port 86 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 i_data[7]
port 87 nsew signal input
rlabel metal2 s 121090 0 121146 800 6 i_data[80]
port 88 nsew signal input
rlabel metal3 s 161701 135328 162501 135448 6 i_data[81]
port 89 nsew signal input
rlabel metal2 s 54758 0 54814 800 6 i_data[8]
port 90 nsew signal input
rlabel metal3 s 0 147568 800 147688 6 i_data[9]
port 91 nsew signal input
rlabel metal3 s 161701 115608 162501 115728 6 i_rst
port 92 nsew signal input
rlabel metal2 s 43166 163845 43222 164645 6 i_we
port 93 nsew signal input
rlabel metal3 s 161701 45568 162501 45688 6 o_data[0]
port 94 nsew signal output
rlabel metal3 s 0 19048 800 19168 6 o_data[10]
port 95 nsew signal output
rlabel metal3 s 0 3408 800 3528 6 o_data[11]
port 96 nsew signal output
rlabel metal2 s 150714 0 150770 800 6 o_data[12]
port 97 nsew signal output
rlabel metal2 s 84382 0 84438 800 6 o_data[13]
port 98 nsew signal output
rlabel metal3 s 161701 84328 162501 84448 6 o_data[14]
port 99 nsew signal output
rlabel metal3 s 0 70048 800 70168 6 o_data[15]
port 100 nsew signal output
rlabel metal3 s 0 50328 800 50448 6 o_data[16]
port 101 nsew signal output
rlabel metal2 s 86958 163845 87014 164645 6 o_data[17]
port 102 nsew signal output
rlabel metal2 s 110142 0 110198 800 6 o_data[18]
port 103 nsew signal output
rlabel metal3 s 0 151648 800 151768 6 o_data[19]
port 104 nsew signal output
rlabel metal3 s 161701 150288 162501 150408 6 o_data[1]
port 105 nsew signal output
rlabel metal3 s 161701 53048 162501 53168 6 o_data[20]
port 106 nsew signal output
rlabel metal2 s 90822 163845 90878 164645 6 o_data[21]
port 107 nsew signal output
rlabel metal3 s 0 30608 800 30728 6 o_data[22]
port 108 nsew signal output
rlabel metal2 s 109498 163845 109554 164645 6 o_data[23]
port 109 nsew signal output
rlabel metal2 s 3238 0 3294 800 6 o_data[24]
port 110 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 o_data[25]
port 111 nsew signal output
rlabel metal3 s 161701 18368 162501 18488 6 o_data[26]
port 112 nsew signal output
rlabel metal3 s 0 23128 800 23248 6 o_data[27]
port 113 nsew signal output
rlabel metal3 s 161701 123088 162501 123208 6 o_data[28]
port 114 nsew signal output
rlabel metal3 s 161701 92488 162501 92608 6 o_data[29]
port 115 nsew signal output
rlabel metal2 s 120446 163845 120502 164645 6 o_data[2]
port 116 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 o_data[30]
port 117 nsew signal output
rlabel metal3 s 161701 38088 162501 38208 6 o_data[31]
port 118 nsew signal output
rlabel metal3 s 161701 95888 162501 96008 6 o_data[32]
port 119 nsew signal output
rlabel metal2 s 54114 163845 54170 164645 6 o_data[33]
port 120 nsew signal output
rlabel metal3 s 161701 65288 162501 65408 6 o_data[34]
port 121 nsew signal output
rlabel metal3 s 161701 2728 162501 2848 6 o_data[35]
port 122 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 o_data[36]
port 123 nsew signal output
rlabel metal3 s 161701 119688 162501 119808 6 o_data[37]
port 124 nsew signal output
rlabel metal2 s 127530 163845 127586 164645 6 o_data[38]
port 125 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 o_data[39]
port 126 nsew signal output
rlabel metal3 s 161701 49648 162501 49768 6 o_data[3]
port 127 nsew signal output
rlabel metal2 s 106278 0 106334 800 6 o_data[40]
port 128 nsew signal output
rlabel metal3 s 161701 6808 162501 6928 6 o_data[41]
port 129 nsew signal output
rlabel metal3 s 0 97248 800 97368 6 o_data[42]
port 130 nsew signal output
rlabel metal2 s 135902 0 135958 800 6 o_data[43]
port 131 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 o_data[44]
port 132 nsew signal output
rlabel metal2 s 66350 0 66406 800 6 o_data[45]
port 133 nsew signal output
rlabel metal3 s 0 61888 800 62008 6 o_data[46]
port 134 nsew signal output
rlabel metal3 s 161701 142808 162501 142928 6 o_data[47]
port 135 nsew signal output
rlabel metal3 s 161701 99968 162501 100088 6 o_data[48]
port 136 nsew signal output
rlabel metal2 s 143630 0 143686 800 6 o_data[49]
port 137 nsew signal output
rlabel metal3 s 0 81608 800 81728 6 o_data[4]
port 138 nsew signal output
rlabel metal3 s 161701 57128 162501 57248 6 o_data[50]
port 139 nsew signal output
rlabel metal3 s 0 108808 800 108928 6 o_data[51]
port 140 nsew signal output
rlabel metal3 s 161701 108128 162501 108248 6 o_data[52]
port 141 nsew signal output
rlabel metal3 s 161701 158448 162501 158568 6 o_data[53]
port 142 nsew signal output
rlabel metal2 s 154578 0 154634 800 6 o_data[54]
port 143 nsew signal output
rlabel metal2 s 161018 163845 161074 164645 6 o_data[55]
port 144 nsew signal output
rlabel metal3 s 0 112208 800 112328 6 o_data[56]
port 145 nsew signal output
rlabel metal3 s 0 120368 800 120488 6 o_data[57]
port 146 nsew signal output
rlabel metal2 s 95330 0 95386 800 6 o_data[58]
port 147 nsew signal output
rlabel metal2 s 18 0 74 800 6 o_data[59]
port 148 nsew signal output
rlabel metal3 s 0 14968 800 15088 6 o_data[5]
port 149 nsew signal output
rlabel metal3 s 0 136008 800 136128 6 o_data[60]
port 150 nsew signal output
rlabel metal2 s 24490 163845 24546 164645 6 o_data[61]
port 151 nsew signal output
rlabel metal2 s 83094 163845 83150 164645 6 o_data[62]
port 152 nsew signal output
rlabel metal3 s 0 104728 800 104848 6 o_data[63]
port 153 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 o_data[64]
port 154 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 o_data[65]
port 155 nsew signal output
rlabel metal2 s 112718 163845 112774 164645 6 o_data[66]
port 156 nsew signal output
rlabel metal2 s 79874 163845 79930 164645 6 o_data[67]
port 157 nsew signal output
rlabel metal2 s 80518 0 80574 800 6 o_data[68]
port 158 nsew signal output
rlabel metal2 s 135258 163845 135314 164645 6 o_data[69]
port 159 nsew signal output
rlabel metal3 s 161701 29928 162501 30048 6 o_data[6]
port 160 nsew signal output
rlabel metal3 s 0 7488 800 7608 6 o_data[70]
port 161 nsew signal output
rlabel metal3 s 0 38768 800 38888 6 o_data[71]
port 162 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 o_data[72]
port 163 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 o_data[73]
port 164 nsew signal output
rlabel metal3 s 0 34688 800 34808 6 o_data[74]
port 165 nsew signal output
rlabel metal3 s 161701 111528 162501 111648 6 o_data[75]
port 166 nsew signal output
rlabel metal2 s 92110 0 92166 800 6 o_data[76]
port 167 nsew signal output
rlabel metal3 s 0 27208 800 27328 6 o_data[77]
port 168 nsew signal output
rlabel metal2 s 116582 163845 116638 164645 6 o_data[78]
port 169 nsew signal output
rlabel metal2 s 2594 163845 2650 164645 6 o_data[79]
port 170 nsew signal output
rlabel metal2 s 28354 163845 28410 164645 6 o_data[7]
port 171 nsew signal output
rlabel metal2 s 114006 0 114062 800 6 o_data[80]
port 172 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 o_data[81]
port 173 nsew signal output
rlabel metal3 s 0 140088 800 140208 6 o_data[8]
port 174 nsew signal output
rlabel metal3 s 161701 76848 162501 76968 6 o_data[9]
port 175 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 162501 164645
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 70933492
string GDS_FILE /home/piotro/ppcpu_caravel/openlane/dffram_rst/runs/22_09_08_23_10/results/signoff/d_dffram_rst.magic.gds
string GDS_START 344736
<< end >>

