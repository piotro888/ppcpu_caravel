// This is the unpowered netlist.
module int_ram (i_clk,
    i_we,
    i_addr,
    i_data,
    o_data);
 input i_clk;
 input i_we;
 input [6:0] i_addr;
 input [15:0] i_data;
 output [15:0] o_data;

 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01676_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04348_;
 wire _04349_;
 wire _04350_;
 wire _04351_;
 wire _04352_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire _04688_;
 wire _04689_;
 wire _04690_;
 wire _04691_;
 wire _04692_;
 wire _04693_;
 wire _04694_;
 wire _04695_;
 wire _04696_;
 wire _04697_;
 wire _04698_;
 wire _04699_;
 wire _04700_;
 wire _04701_;
 wire _04702_;
 wire _04703_;
 wire _04704_;
 wire _04705_;
 wire _04706_;
 wire _04707_;
 wire _04708_;
 wire _04709_;
 wire _04710_;
 wire _04711_;
 wire _04712_;
 wire _04713_;
 wire _04714_;
 wire _04715_;
 wire _04716_;
 wire _04717_;
 wire _04718_;
 wire _04719_;
 wire _04720_;
 wire _04721_;
 wire _04722_;
 wire _04723_;
 wire _04724_;
 wire _04725_;
 wire _04726_;
 wire _04727_;
 wire _04728_;
 wire _04729_;
 wire _04730_;
 wire _04731_;
 wire _04732_;
 wire _04733_;
 wire _04734_;
 wire _04735_;
 wire _04736_;
 wire _04737_;
 wire _04738_;
 wire _04739_;
 wire _04740_;
 wire _04741_;
 wire _04742_;
 wire _04743_;
 wire _04744_;
 wire _04745_;
 wire _04746_;
 wire _04747_;
 wire _04748_;
 wire _04749_;
 wire _04750_;
 wire _04751_;
 wire _04752_;
 wire _04753_;
 wire _04754_;
 wire _04755_;
 wire _04756_;
 wire _04757_;
 wire _04758_;
 wire _04759_;
 wire _04760_;
 wire _04761_;
 wire _04762_;
 wire _04763_;
 wire _04764_;
 wire _04765_;
 wire _04766_;
 wire _04767_;
 wire _04768_;
 wire _04769_;
 wire _04770_;
 wire _04771_;
 wire _04772_;
 wire _04773_;
 wire _04774_;
 wire _04775_;
 wire _04776_;
 wire _04777_;
 wire _04778_;
 wire _04779_;
 wire _04780_;
 wire _04781_;
 wire _04782_;
 wire _04783_;
 wire _04784_;
 wire _04785_;
 wire _04786_;
 wire _04787_;
 wire _04788_;
 wire _04789_;
 wire _04790_;
 wire _04791_;
 wire _04792_;
 wire _04793_;
 wire _04794_;
 wire _04795_;
 wire _04796_;
 wire _04797_;
 wire _04798_;
 wire _04799_;
 wire _04800_;
 wire _04801_;
 wire _04802_;
 wire _04803_;
 wire _04804_;
 wire _04805_;
 wire _04806_;
 wire _04807_;
 wire _04808_;
 wire _04809_;
 wire _04810_;
 wire _04811_;
 wire _04812_;
 wire _04813_;
 wire _04814_;
 wire _04815_;
 wire _04816_;
 wire _04817_;
 wire _04818_;
 wire _04819_;
 wire _04820_;
 wire _04821_;
 wire _04822_;
 wire _04823_;
 wire _04824_;
 wire _04825_;
 wire _04826_;
 wire _04827_;
 wire _04828_;
 wire _04829_;
 wire _04830_;
 wire _04831_;
 wire _04832_;
 wire _04833_;
 wire _04834_;
 wire _04835_;
 wire _04836_;
 wire _04837_;
 wire _04838_;
 wire _04839_;
 wire _04840_;
 wire _04841_;
 wire _04842_;
 wire _04843_;
 wire _04844_;
 wire _04845_;
 wire _04846_;
 wire _04847_;
 wire _04848_;
 wire _04849_;
 wire _04850_;
 wire _04851_;
 wire _04852_;
 wire _04853_;
 wire _04854_;
 wire _04855_;
 wire _04856_;
 wire _04857_;
 wire _04858_;
 wire _04859_;
 wire _04860_;
 wire _04861_;
 wire _04862_;
 wire _04863_;
 wire _04864_;
 wire _04865_;
 wire _04866_;
 wire _04867_;
 wire _04868_;
 wire _04869_;
 wire _04870_;
 wire _04871_;
 wire _04872_;
 wire _04873_;
 wire _04874_;
 wire _04875_;
 wire _04876_;
 wire _04877_;
 wire _04878_;
 wire _04879_;
 wire _04880_;
 wire _04881_;
 wire _04882_;
 wire _04883_;
 wire _04884_;
 wire _04885_;
 wire _04886_;
 wire _04887_;
 wire _04888_;
 wire _04889_;
 wire _04890_;
 wire _04891_;
 wire _04892_;
 wire _04893_;
 wire _04894_;
 wire _04895_;
 wire _04896_;
 wire _04897_;
 wire _04898_;
 wire _04899_;
 wire _04900_;
 wire _04901_;
 wire _04902_;
 wire _04903_;
 wire _04904_;
 wire _04905_;
 wire _04906_;
 wire _04907_;
 wire _04908_;
 wire _04909_;
 wire _04910_;
 wire _04911_;
 wire _04912_;
 wire _04913_;
 wire _04914_;
 wire _04915_;
 wire _04916_;
 wire _04917_;
 wire _04918_;
 wire _04919_;
 wire _04920_;
 wire _04921_;
 wire _04922_;
 wire _04923_;
 wire _04924_;
 wire _04925_;
 wire _04926_;
 wire _04927_;
 wire _04928_;
 wire _04929_;
 wire _04930_;
 wire _04931_;
 wire _04932_;
 wire _04933_;
 wire _04934_;
 wire _04935_;
 wire _04936_;
 wire _04937_;
 wire _04938_;
 wire _04939_;
 wire _04940_;
 wire _04941_;
 wire _04942_;
 wire _04943_;
 wire _04944_;
 wire _04945_;
 wire _04946_;
 wire _04947_;
 wire _04948_;
 wire _04949_;
 wire _04950_;
 wire _04951_;
 wire _04952_;
 wire _04953_;
 wire _04954_;
 wire _04955_;
 wire _04956_;
 wire _04957_;
 wire _04958_;
 wire _04959_;
 wire _04960_;
 wire _04961_;
 wire _04962_;
 wire _04963_;
 wire _04964_;
 wire _04965_;
 wire _04966_;
 wire _04967_;
 wire _04968_;
 wire _04969_;
 wire _04970_;
 wire _04971_;
 wire _04972_;
 wire _04973_;
 wire _04974_;
 wire _04975_;
 wire _04976_;
 wire _04977_;
 wire _04978_;
 wire _04979_;
 wire _04980_;
 wire _04981_;
 wire _04982_;
 wire _04983_;
 wire _04984_;
 wire _04985_;
 wire _04986_;
 wire _04987_;
 wire _04988_;
 wire _04989_;
 wire _04990_;
 wire _04991_;
 wire _04992_;
 wire _04993_;
 wire _04994_;
 wire _04995_;
 wire _04996_;
 wire _04997_;
 wire _04998_;
 wire _04999_;
 wire _05000_;
 wire _05001_;
 wire _05002_;
 wire _05003_;
 wire _05004_;
 wire _05005_;
 wire _05006_;
 wire _05007_;
 wire _05008_;
 wire _05009_;
 wire _05010_;
 wire _05011_;
 wire _05012_;
 wire _05013_;
 wire _05014_;
 wire _05015_;
 wire _05016_;
 wire _05017_;
 wire _05018_;
 wire _05019_;
 wire _05020_;
 wire _05021_;
 wire _05022_;
 wire _05023_;
 wire _05024_;
 wire _05025_;
 wire _05026_;
 wire _05027_;
 wire _05028_;
 wire _05029_;
 wire _05030_;
 wire _05031_;
 wire _05032_;
 wire _05033_;
 wire _05034_;
 wire _05035_;
 wire _05036_;
 wire _05037_;
 wire _05038_;
 wire _05039_;
 wire _05040_;
 wire _05041_;
 wire _05042_;
 wire _05043_;
 wire _05044_;
 wire _05045_;
 wire _05046_;
 wire _05047_;
 wire _05048_;
 wire _05049_;
 wire _05050_;
 wire _05051_;
 wire _05052_;
 wire _05053_;
 wire _05054_;
 wire _05055_;
 wire _05056_;
 wire _05057_;
 wire _05058_;
 wire _05059_;
 wire _05060_;
 wire _05061_;
 wire _05062_;
 wire _05063_;
 wire _05064_;
 wire _05065_;
 wire _05066_;
 wire _05067_;
 wire _05068_;
 wire _05069_;
 wire _05070_;
 wire _05071_;
 wire _05072_;
 wire _05073_;
 wire _05074_;
 wire _05075_;
 wire _05076_;
 wire _05077_;
 wire _05078_;
 wire _05079_;
 wire _05080_;
 wire _05081_;
 wire _05082_;
 wire _05083_;
 wire _05084_;
 wire _05085_;
 wire _05086_;
 wire _05087_;
 wire _05088_;
 wire _05089_;
 wire _05090_;
 wire _05091_;
 wire _05092_;
 wire _05093_;
 wire _05094_;
 wire _05095_;
 wire _05096_;
 wire _05097_;
 wire _05098_;
 wire _05099_;
 wire _05100_;
 wire _05101_;
 wire _05102_;
 wire _05103_;
 wire _05104_;
 wire _05105_;
 wire _05106_;
 wire _05107_;
 wire _05108_;
 wire _05109_;
 wire _05110_;
 wire _05111_;
 wire _05112_;
 wire _05113_;
 wire _05114_;
 wire _05115_;
 wire _05116_;
 wire _05117_;
 wire _05118_;
 wire _05119_;
 wire _05120_;
 wire _05121_;
 wire _05122_;
 wire _05123_;
 wire _05124_;
 wire _05125_;
 wire _05126_;
 wire _05127_;
 wire _05128_;
 wire _05129_;
 wire _05130_;
 wire _05131_;
 wire _05132_;
 wire _05133_;
 wire _05134_;
 wire _05135_;
 wire _05136_;
 wire _05137_;
 wire _05138_;
 wire _05139_;
 wire _05140_;
 wire _05141_;
 wire _05142_;
 wire _05143_;
 wire _05144_;
 wire _05145_;
 wire _05146_;
 wire _05147_;
 wire _05148_;
 wire _05149_;
 wire _05150_;
 wire _05151_;
 wire _05152_;
 wire _05153_;
 wire _05154_;
 wire _05155_;
 wire _05156_;
 wire _05157_;
 wire _05158_;
 wire _05159_;
 wire _05160_;
 wire _05161_;
 wire _05162_;
 wire _05163_;
 wire _05164_;
 wire _05165_;
 wire _05166_;
 wire _05167_;
 wire _05168_;
 wire _05169_;
 wire _05170_;
 wire _05171_;
 wire _05172_;
 wire _05173_;
 wire _05174_;
 wire _05175_;
 wire _05176_;
 wire _05177_;
 wire _05178_;
 wire _05179_;
 wire _05180_;
 wire _05181_;
 wire _05182_;
 wire _05183_;
 wire _05184_;
 wire _05185_;
 wire _05186_;
 wire _05187_;
 wire _05188_;
 wire _05189_;
 wire _05190_;
 wire _05191_;
 wire _05192_;
 wire _05193_;
 wire _05194_;
 wire _05195_;
 wire _05196_;
 wire _05197_;
 wire _05198_;
 wire _05199_;
 wire _05200_;
 wire _05201_;
 wire _05202_;
 wire _05203_;
 wire _05204_;
 wire _05205_;
 wire _05206_;
 wire _05207_;
 wire _05208_;
 wire _05209_;
 wire _05210_;
 wire _05211_;
 wire _05212_;
 wire _05213_;
 wire _05214_;
 wire _05215_;
 wire _05216_;
 wire _05217_;
 wire _05218_;
 wire _05219_;
 wire _05220_;
 wire _05221_;
 wire _05222_;
 wire _05223_;
 wire _05224_;
 wire _05225_;
 wire _05226_;
 wire _05227_;
 wire _05228_;
 wire _05229_;
 wire _05230_;
 wire _05231_;
 wire _05232_;
 wire _05233_;
 wire _05234_;
 wire _05235_;
 wire _05236_;
 wire _05237_;
 wire _05238_;
 wire _05239_;
 wire _05240_;
 wire _05241_;
 wire _05242_;
 wire _05243_;
 wire _05244_;
 wire _05245_;
 wire _05246_;
 wire _05247_;
 wire _05248_;
 wire _05249_;
 wire _05250_;
 wire _05251_;
 wire _05252_;
 wire _05253_;
 wire _05254_;
 wire _05255_;
 wire _05256_;
 wire _05257_;
 wire _05258_;
 wire _05259_;
 wire _05260_;
 wire _05261_;
 wire _05262_;
 wire _05263_;
 wire _05264_;
 wire _05265_;
 wire _05266_;
 wire _05267_;
 wire _05268_;
 wire _05269_;
 wire _05270_;
 wire _05271_;
 wire _05272_;
 wire _05273_;
 wire _05274_;
 wire _05275_;
 wire _05276_;
 wire _05277_;
 wire _05278_;
 wire _05279_;
 wire _05280_;
 wire _05281_;
 wire _05282_;
 wire _05283_;
 wire _05284_;
 wire _05285_;
 wire _05286_;
 wire _05287_;
 wire _05288_;
 wire _05289_;
 wire _05290_;
 wire _05291_;
 wire _05292_;
 wire _05293_;
 wire _05294_;
 wire _05295_;
 wire _05296_;
 wire _05297_;
 wire _05298_;
 wire _05299_;
 wire _05300_;
 wire _05301_;
 wire _05302_;
 wire _05303_;
 wire _05304_;
 wire _05305_;
 wire _05306_;
 wire _05307_;
 wire _05308_;
 wire _05309_;
 wire _05310_;
 wire _05311_;
 wire _05312_;
 wire _05313_;
 wire _05314_;
 wire _05315_;
 wire _05316_;
 wire _05317_;
 wire _05318_;
 wire _05319_;
 wire _05320_;
 wire _05321_;
 wire _05322_;
 wire _05323_;
 wire _05324_;
 wire _05325_;
 wire _05326_;
 wire _05327_;
 wire _05328_;
 wire _05329_;
 wire _05330_;
 wire _05331_;
 wire _05332_;
 wire _05333_;
 wire _05334_;
 wire _05335_;
 wire _05336_;
 wire _05337_;
 wire _05338_;
 wire _05339_;
 wire _05340_;
 wire _05341_;
 wire _05342_;
 wire _05343_;
 wire _05344_;
 wire _05345_;
 wire _05346_;
 wire _05347_;
 wire _05348_;
 wire _05349_;
 wire _05350_;
 wire _05351_;
 wire _05352_;
 wire _05353_;
 wire _05354_;
 wire _05355_;
 wire _05356_;
 wire _05357_;
 wire _05358_;
 wire _05359_;
 wire _05360_;
 wire _05361_;
 wire _05362_;
 wire _05363_;
 wire _05364_;
 wire _05365_;
 wire _05366_;
 wire _05367_;
 wire _05368_;
 wire _05369_;
 wire _05370_;
 wire _05371_;
 wire _05372_;
 wire _05373_;
 wire _05374_;
 wire _05375_;
 wire _05376_;
 wire _05377_;
 wire _05378_;
 wire _05379_;
 wire _05380_;
 wire _05381_;
 wire _05382_;
 wire _05383_;
 wire _05384_;
 wire _05385_;
 wire _05386_;
 wire _05387_;
 wire _05388_;
 wire _05389_;
 wire _05390_;
 wire _05391_;
 wire _05392_;
 wire _05393_;
 wire _05394_;
 wire _05395_;
 wire _05396_;
 wire _05397_;
 wire _05398_;
 wire _05399_;
 wire _05400_;
 wire _05401_;
 wire _05402_;
 wire _05403_;
 wire _05404_;
 wire _05405_;
 wire _05406_;
 wire _05407_;
 wire _05408_;
 wire _05409_;
 wire _05410_;
 wire _05411_;
 wire _05412_;
 wire _05413_;
 wire _05414_;
 wire _05415_;
 wire _05416_;
 wire _05417_;
 wire _05418_;
 wire _05419_;
 wire _05420_;
 wire _05421_;
 wire _05422_;
 wire _05423_;
 wire _05424_;
 wire _05425_;
 wire _05426_;
 wire _05427_;
 wire _05428_;
 wire _05429_;
 wire _05430_;
 wire _05431_;
 wire _05432_;
 wire _05433_;
 wire _05434_;
 wire _05435_;
 wire _05436_;
 wire _05437_;
 wire _05438_;
 wire _05439_;
 wire _05440_;
 wire _05441_;
 wire _05442_;
 wire _05443_;
 wire _05444_;
 wire _05445_;
 wire _05446_;
 wire _05447_;
 wire _05448_;
 wire _05449_;
 wire _05450_;
 wire _05451_;
 wire _05452_;
 wire _05453_;
 wire _05454_;
 wire _05455_;
 wire _05456_;
 wire _05457_;
 wire _05458_;
 wire _05459_;
 wire _05460_;
 wire _05461_;
 wire _05462_;
 wire _05463_;
 wire _05464_;
 wire _05465_;
 wire _05466_;
 wire _05467_;
 wire _05468_;
 wire _05469_;
 wire _05470_;
 wire _05471_;
 wire _05472_;
 wire _05473_;
 wire _05474_;
 wire _05475_;
 wire _05476_;
 wire _05477_;
 wire _05478_;
 wire _05479_;
 wire _05480_;
 wire _05481_;
 wire _05482_;
 wire _05483_;
 wire _05484_;
 wire _05485_;
 wire _05486_;
 wire _05487_;
 wire _05488_;
 wire _05489_;
 wire _05490_;
 wire _05491_;
 wire _05492_;
 wire _05493_;
 wire _05494_;
 wire _05495_;
 wire _05496_;
 wire _05497_;
 wire _05498_;
 wire _05499_;
 wire _05500_;
 wire _05501_;
 wire _05502_;
 wire _05503_;
 wire _05504_;
 wire _05505_;
 wire _05506_;
 wire _05507_;
 wire _05508_;
 wire _05509_;
 wire _05510_;
 wire _05511_;
 wire _05512_;
 wire _05513_;
 wire _05514_;
 wire _05515_;
 wire _05516_;
 wire _05517_;
 wire _05518_;
 wire _05519_;
 wire _05520_;
 wire _05521_;
 wire _05522_;
 wire _05523_;
 wire _05524_;
 wire _05525_;
 wire _05526_;
 wire _05527_;
 wire _05528_;
 wire _05529_;
 wire _05530_;
 wire _05531_;
 wire _05532_;
 wire _05533_;
 wire _05534_;
 wire _05535_;
 wire _05536_;
 wire _05537_;
 wire _05538_;
 wire _05539_;
 wire _05540_;
 wire _05541_;
 wire _05542_;
 wire _05543_;
 wire _05544_;
 wire _05545_;
 wire _05546_;
 wire _05547_;
 wire _05548_;
 wire _05549_;
 wire _05550_;
 wire _05551_;
 wire _05552_;
 wire _05553_;
 wire _05554_;
 wire _05555_;
 wire _05556_;
 wire _05557_;
 wire _05558_;
 wire _05559_;
 wire _05560_;
 wire _05561_;
 wire _05562_;
 wire _05563_;
 wire _05564_;
 wire _05565_;
 wire _05566_;
 wire _05567_;
 wire _05568_;
 wire _05569_;
 wire _05570_;
 wire _05571_;
 wire _05572_;
 wire _05573_;
 wire _05574_;
 wire _05575_;
 wire _05576_;
 wire _05577_;
 wire _05578_;
 wire _05579_;
 wire _05580_;
 wire _05581_;
 wire _05582_;
 wire _05583_;
 wire _05584_;
 wire _05585_;
 wire _05586_;
 wire _05587_;
 wire _05588_;
 wire _05589_;
 wire _05590_;
 wire _05591_;
 wire _05592_;
 wire _05593_;
 wire _05594_;
 wire _05595_;
 wire _05596_;
 wire _05597_;
 wire _05598_;
 wire _05599_;
 wire _05600_;
 wire _05601_;
 wire _05602_;
 wire _05603_;
 wire _05604_;
 wire _05605_;
 wire _05606_;
 wire _05607_;
 wire _05608_;
 wire _05609_;
 wire _05610_;
 wire _05611_;
 wire _05612_;
 wire _05613_;
 wire _05614_;
 wire _05615_;
 wire _05616_;
 wire _05617_;
 wire _05618_;
 wire _05619_;
 wire _05620_;
 wire _05621_;
 wire _05622_;
 wire _05623_;
 wire _05624_;
 wire _05625_;
 wire _05626_;
 wire _05627_;
 wire _05628_;
 wire _05629_;
 wire _05630_;
 wire _05631_;
 wire _05632_;
 wire _05633_;
 wire _05634_;
 wire _05635_;
 wire _05636_;
 wire _05637_;
 wire _05638_;
 wire _05639_;
 wire _05640_;
 wire _05641_;
 wire _05642_;
 wire _05643_;
 wire _05644_;
 wire _05645_;
 wire _05646_;
 wire _05647_;
 wire _05648_;
 wire _05649_;
 wire _05650_;
 wire _05651_;
 wire _05652_;
 wire _05653_;
 wire _05654_;
 wire _05655_;
 wire _05656_;
 wire _05657_;
 wire _05658_;
 wire _05659_;
 wire _05660_;
 wire _05661_;
 wire _05662_;
 wire _05663_;
 wire _05664_;
 wire _05665_;
 wire _05666_;
 wire _05667_;
 wire _05668_;
 wire _05669_;
 wire _05670_;
 wire _05671_;
 wire _05672_;
 wire _05673_;
 wire _05674_;
 wire _05675_;
 wire _05676_;
 wire _05677_;
 wire _05678_;
 wire _05679_;
 wire _05680_;
 wire _05681_;
 wire _05682_;
 wire _05683_;
 wire _05684_;
 wire _05685_;
 wire _05686_;
 wire _05687_;
 wire _05688_;
 wire _05689_;
 wire _05690_;
 wire _05691_;
 wire _05692_;
 wire _05693_;
 wire _05694_;
 wire _05695_;
 wire _05696_;
 wire _05697_;
 wire _05698_;
 wire _05699_;
 wire _05700_;
 wire _05701_;
 wire _05702_;
 wire _05703_;
 wire _05704_;
 wire _05705_;
 wire _05706_;
 wire _05707_;
 wire _05708_;
 wire _05709_;
 wire _05710_;
 wire _05711_;
 wire _05712_;
 wire _05713_;
 wire _05714_;
 wire _05715_;
 wire _05716_;
 wire _05717_;
 wire _05718_;
 wire _05719_;
 wire _05720_;
 wire _05721_;
 wire _05722_;
 wire _05723_;
 wire _05724_;
 wire _05725_;
 wire _05726_;
 wire _05727_;
 wire _05728_;
 wire _05729_;
 wire _05730_;
 wire _05731_;
 wire _05732_;
 wire _05733_;
 wire _05734_;
 wire _05735_;
 wire _05736_;
 wire _05737_;
 wire _05738_;
 wire _05739_;
 wire _05740_;
 wire _05741_;
 wire _05742_;
 wire _05743_;
 wire _05744_;
 wire _05745_;
 wire _05746_;
 wire _05747_;
 wire _05748_;
 wire _05749_;
 wire _05750_;
 wire _05751_;
 wire _05752_;
 wire _05753_;
 wire _05754_;
 wire _05755_;
 wire _05756_;
 wire _05757_;
 wire _05758_;
 wire _05759_;
 wire _05760_;
 wire _05761_;
 wire _05762_;
 wire _05763_;
 wire _05764_;
 wire _05765_;
 wire _05766_;
 wire _05767_;
 wire _05768_;
 wire _05769_;
 wire _05770_;
 wire _05771_;
 wire _05772_;
 wire _05773_;
 wire _05774_;
 wire _05775_;
 wire _05776_;
 wire _05777_;
 wire _05778_;
 wire _05779_;
 wire _05780_;
 wire _05781_;
 wire _05782_;
 wire _05783_;
 wire _05784_;
 wire _05785_;
 wire _05786_;
 wire _05787_;
 wire _05788_;
 wire _05789_;
 wire _05790_;
 wire _05791_;
 wire _05792_;
 wire _05793_;
 wire _05794_;
 wire _05795_;
 wire _05796_;
 wire _05797_;
 wire _05798_;
 wire _05799_;
 wire _05800_;
 wire _05801_;
 wire _05802_;
 wire _05803_;
 wire _05804_;
 wire _05805_;
 wire _05806_;
 wire _05807_;
 wire _05808_;
 wire _05809_;
 wire _05810_;
 wire _05811_;
 wire _05812_;
 wire _05813_;
 wire _05814_;
 wire _05815_;
 wire _05816_;
 wire _05817_;
 wire _05818_;
 wire _05819_;
 wire _05820_;
 wire _05821_;
 wire _05822_;
 wire _05823_;
 wire _05824_;
 wire _05825_;
 wire _05826_;
 wire _05827_;
 wire _05828_;
 wire _05829_;
 wire _05830_;
 wire _05831_;
 wire _05832_;
 wire _05833_;
 wire _05834_;
 wire _05835_;
 wire _05836_;
 wire _05837_;
 wire _05838_;
 wire _05839_;
 wire _05840_;
 wire _05841_;
 wire _05842_;
 wire _05843_;
 wire _05844_;
 wire _05845_;
 wire _05846_;
 wire _05847_;
 wire _05848_;
 wire _05849_;
 wire _05850_;
 wire _05851_;
 wire _05852_;
 wire _05853_;
 wire _05854_;
 wire _05855_;
 wire _05856_;
 wire _05857_;
 wire _05858_;
 wire _05859_;
 wire _05860_;
 wire _05861_;
 wire _05862_;
 wire _05863_;
 wire _05864_;
 wire _05865_;
 wire _05866_;
 wire _05867_;
 wire _05868_;
 wire _05869_;
 wire _05870_;
 wire _05871_;
 wire _05872_;
 wire _05873_;
 wire _05874_;
 wire _05875_;
 wire _05876_;
 wire _05877_;
 wire _05878_;
 wire _05879_;
 wire _05880_;
 wire _05881_;
 wire _05882_;
 wire _05883_;
 wire _05884_;
 wire _05885_;
 wire _05886_;
 wire _05887_;
 wire _05888_;
 wire _05889_;
 wire _05890_;
 wire _05891_;
 wire _05892_;
 wire _05893_;
 wire _05894_;
 wire _05895_;
 wire _05896_;
 wire _05897_;
 wire _05898_;
 wire _05899_;
 wire _05900_;
 wire _05901_;
 wire _05902_;
 wire _05903_;
 wire _05904_;
 wire _05905_;
 wire _05906_;
 wire _05907_;
 wire _05908_;
 wire _05909_;
 wire _05910_;
 wire _05911_;
 wire _05912_;
 wire _05913_;
 wire _05914_;
 wire _05915_;
 wire _05916_;
 wire _05917_;
 wire _05918_;
 wire _05919_;
 wire _05920_;
 wire _05921_;
 wire _05922_;
 wire _05923_;
 wire _05924_;
 wire _05925_;
 wire _05926_;
 wire _05927_;
 wire _05928_;
 wire _05929_;
 wire _05930_;
 wire _05931_;
 wire _05932_;
 wire _05933_;
 wire _05934_;
 wire _05935_;
 wire _05936_;
 wire _05937_;
 wire _05938_;
 wire _05939_;
 wire _05940_;
 wire _05941_;
 wire _05942_;
 wire _05943_;
 wire _05944_;
 wire _05945_;
 wire _05946_;
 wire _05947_;
 wire _05948_;
 wire _05949_;
 wire _05950_;
 wire _05951_;
 wire _05952_;
 wire _05953_;
 wire _05954_;
 wire _05955_;
 wire _05956_;
 wire _05957_;
 wire _05958_;
 wire _05959_;
 wire _05960_;
 wire _05961_;
 wire _05962_;
 wire _05963_;
 wire _05964_;
 wire _05965_;
 wire _05966_;
 wire _05967_;
 wire _05968_;
 wire _05969_;
 wire _05970_;
 wire _05971_;
 wire _05972_;
 wire _05973_;
 wire _05974_;
 wire _05975_;
 wire _05976_;
 wire _05977_;
 wire _05978_;
 wire _05979_;
 wire _05980_;
 wire _05981_;
 wire _05982_;
 wire _05983_;
 wire _05984_;
 wire _05985_;
 wire _05986_;
 wire _05987_;
 wire _05988_;
 wire _05989_;
 wire _05990_;
 wire _05991_;
 wire _05992_;
 wire _05993_;
 wire _05994_;
 wire _05995_;
 wire _05996_;
 wire _05997_;
 wire _05998_;
 wire _05999_;
 wire _06000_;
 wire _06001_;
 wire _06002_;
 wire _06003_;
 wire _06004_;
 wire _06005_;
 wire _06006_;
 wire _06007_;
 wire _06008_;
 wire _06009_;
 wire _06010_;
 wire _06011_;
 wire _06012_;
 wire _06013_;
 wire _06014_;
 wire _06015_;
 wire _06016_;
 wire _06017_;
 wire _06018_;
 wire _06019_;
 wire _06020_;
 wire _06021_;
 wire _06022_;
 wire _06023_;
 wire _06024_;
 wire _06025_;
 wire _06026_;
 wire _06027_;
 wire _06028_;
 wire _06029_;
 wire _06030_;
 wire _06031_;
 wire _06032_;
 wire _06033_;
 wire _06034_;
 wire _06035_;
 wire _06036_;
 wire _06037_;
 wire _06038_;
 wire _06039_;
 wire _06040_;
 wire _06041_;
 wire _06042_;
 wire _06043_;
 wire _06044_;
 wire _06045_;
 wire _06046_;
 wire _06047_;
 wire _06048_;
 wire _06049_;
 wire _06050_;
 wire _06051_;
 wire _06052_;
 wire _06053_;
 wire _06054_;
 wire _06055_;
 wire _06056_;
 wire _06057_;
 wire _06058_;
 wire _06059_;
 wire _06060_;
 wire _06061_;
 wire _06062_;
 wire _06063_;
 wire _06064_;
 wire _06065_;
 wire _06066_;
 wire _06067_;
 wire _06068_;
 wire _06069_;
 wire _06070_;
 wire _06071_;
 wire _06072_;
 wire _06073_;
 wire _06074_;
 wire _06075_;
 wire _06076_;
 wire _06077_;
 wire _06078_;
 wire _06079_;
 wire _06080_;
 wire _06081_;
 wire _06082_;
 wire _06083_;
 wire _06084_;
 wire _06085_;
 wire _06086_;
 wire _06087_;
 wire _06088_;
 wire _06089_;
 wire _06090_;
 wire _06091_;
 wire _06092_;
 wire _06093_;
 wire _06094_;
 wire _06095_;
 wire _06096_;
 wire _06097_;
 wire _06098_;
 wire _06099_;
 wire _06100_;
 wire _06101_;
 wire _06102_;
 wire _06103_;
 wire _06104_;
 wire _06105_;
 wire _06106_;
 wire _06107_;
 wire _06108_;
 wire _06109_;
 wire _06110_;
 wire _06111_;
 wire _06112_;
 wire _06113_;
 wire _06114_;
 wire _06115_;
 wire _06116_;
 wire _06117_;
 wire _06118_;
 wire _06119_;
 wire _06120_;
 wire _06121_;
 wire _06122_;
 wire _06123_;
 wire _06124_;
 wire _06125_;
 wire _06126_;
 wire _06127_;
 wire _06128_;
 wire _06129_;
 wire _06130_;
 wire _06131_;
 wire _06132_;
 wire _06133_;
 wire _06134_;
 wire _06135_;
 wire _06136_;
 wire _06137_;
 wire _06138_;
 wire _06139_;
 wire _06140_;
 wire _06141_;
 wire _06142_;
 wire _06143_;
 wire _06144_;
 wire _06145_;
 wire _06146_;
 wire _06147_;
 wire _06148_;
 wire _06149_;
 wire _06150_;
 wire _06151_;
 wire _06152_;
 wire _06153_;
 wire _06154_;
 wire _06155_;
 wire _06156_;
 wire _06157_;
 wire _06158_;
 wire _06159_;
 wire _06160_;
 wire _06161_;
 wire _06162_;
 wire _06163_;
 wire _06164_;
 wire _06165_;
 wire _06166_;
 wire _06167_;
 wire _06168_;
 wire _06169_;
 wire _06170_;
 wire _06171_;
 wire _06172_;
 wire _06173_;
 wire _06174_;
 wire _06175_;
 wire _06176_;
 wire _06177_;
 wire _06178_;
 wire _06179_;
 wire _06180_;
 wire _06181_;
 wire _06182_;
 wire _06183_;
 wire _06184_;
 wire _06185_;
 wire _06186_;
 wire _06187_;
 wire _06188_;
 wire _06189_;
 wire _06190_;
 wire _06191_;
 wire _06192_;
 wire _06193_;
 wire _06194_;
 wire _06195_;
 wire _06196_;
 wire _06197_;
 wire _06198_;
 wire _06199_;
 wire _06200_;
 wire _06201_;
 wire _06202_;
 wire _06203_;
 wire _06204_;
 wire _06205_;
 wire _06206_;
 wire _06207_;
 wire _06208_;
 wire _06209_;
 wire _06210_;
 wire _06211_;
 wire _06212_;
 wire _06213_;
 wire _06214_;
 wire _06215_;
 wire _06216_;
 wire _06217_;
 wire _06218_;
 wire _06219_;
 wire _06220_;
 wire _06221_;
 wire _06222_;
 wire _06223_;
 wire _06224_;
 wire _06225_;
 wire _06226_;
 wire _06227_;
 wire _06228_;
 wire _06229_;
 wire _06230_;
 wire _06231_;
 wire _06232_;
 wire _06233_;
 wire _06234_;
 wire _06235_;
 wire _06236_;
 wire _06237_;
 wire _06238_;
 wire _06239_;
 wire _06240_;
 wire _06241_;
 wire _06242_;
 wire _06243_;
 wire _06244_;
 wire _06245_;
 wire _06246_;
 wire _06247_;
 wire _06248_;
 wire _06249_;
 wire _06250_;
 wire _06251_;
 wire _06252_;
 wire _06253_;
 wire _06254_;
 wire _06255_;
 wire _06256_;
 wire _06257_;
 wire _06258_;
 wire _06259_;
 wire _06260_;
 wire _06261_;
 wire _06262_;
 wire _06263_;
 wire _06264_;
 wire _06265_;
 wire _06266_;
 wire _06267_;
 wire _06268_;
 wire _06269_;
 wire _06270_;
 wire _06271_;
 wire _06272_;
 wire _06273_;
 wire _06274_;
 wire _06275_;
 wire _06276_;
 wire _06277_;
 wire _06278_;
 wire _06279_;
 wire _06280_;
 wire _06281_;
 wire _06282_;
 wire _06283_;
 wire _06284_;
 wire _06285_;
 wire _06286_;
 wire _06287_;
 wire _06288_;
 wire _06289_;
 wire _06290_;
 wire _06291_;
 wire _06292_;
 wire _06293_;
 wire _06294_;
 wire _06295_;
 wire _06296_;
 wire _06297_;
 wire _06298_;
 wire _06299_;
 wire _06300_;
 wire _06301_;
 wire _06302_;
 wire _06303_;
 wire _06304_;
 wire _06305_;
 wire _06306_;
 wire _06307_;
 wire _06308_;
 wire _06309_;
 wire _06310_;
 wire _06311_;
 wire _06312_;
 wire _06313_;
 wire _06314_;
 wire _06315_;
 wire _06316_;
 wire _06317_;
 wire _06318_;
 wire _06319_;
 wire _06320_;
 wire _06321_;
 wire _06322_;
 wire _06323_;
 wire _06324_;
 wire _06325_;
 wire _06326_;
 wire _06327_;
 wire _06328_;
 wire _06329_;
 wire _06330_;
 wire _06331_;
 wire _06332_;
 wire _06333_;
 wire _06334_;
 wire _06335_;
 wire _06336_;
 wire _06337_;
 wire _06338_;
 wire _06339_;
 wire _06340_;
 wire _06341_;
 wire _06342_;
 wire _06343_;
 wire _06344_;
 wire _06345_;
 wire _06346_;
 wire _06347_;
 wire _06348_;
 wire _06349_;
 wire _06350_;
 wire _06351_;
 wire _06352_;
 wire _06353_;
 wire _06354_;
 wire _06355_;
 wire _06356_;
 wire _06357_;
 wire _06358_;
 wire _06359_;
 wire _06360_;
 wire _06361_;
 wire _06362_;
 wire _06363_;
 wire _06364_;
 wire _06365_;
 wire _06366_;
 wire _06367_;
 wire _06368_;
 wire _06369_;
 wire _06370_;
 wire _06371_;
 wire _06372_;
 wire _06373_;
 wire _06374_;
 wire _06375_;
 wire _06376_;
 wire _06377_;
 wire _06378_;
 wire _06379_;
 wire _06380_;
 wire _06381_;
 wire _06382_;
 wire _06383_;
 wire _06384_;
 wire _06385_;
 wire _06386_;
 wire _06387_;
 wire _06388_;
 wire _06389_;
 wire _06390_;
 wire _06391_;
 wire _06392_;
 wire _06393_;
 wire _06394_;
 wire _06395_;
 wire _06396_;
 wire _06397_;
 wire _06398_;
 wire _06399_;
 wire _06400_;
 wire _06401_;
 wire _06402_;
 wire _06403_;
 wire _06404_;
 wire _06405_;
 wire \mem[0][0] ;
 wire \mem[0][10] ;
 wire \mem[0][11] ;
 wire \mem[0][12] ;
 wire \mem[0][13] ;
 wire \mem[0][14] ;
 wire \mem[0][15] ;
 wire \mem[0][1] ;
 wire \mem[0][2] ;
 wire \mem[0][3] ;
 wire \mem[0][4] ;
 wire \mem[0][5] ;
 wire \mem[0][6] ;
 wire \mem[0][7] ;
 wire \mem[0][8] ;
 wire \mem[0][9] ;
 wire \mem[100][0] ;
 wire \mem[100][10] ;
 wire \mem[100][11] ;
 wire \mem[100][12] ;
 wire \mem[100][13] ;
 wire \mem[100][14] ;
 wire \mem[100][15] ;
 wire \mem[100][1] ;
 wire \mem[100][2] ;
 wire \mem[100][3] ;
 wire \mem[100][4] ;
 wire \mem[100][5] ;
 wire \mem[100][6] ;
 wire \mem[100][7] ;
 wire \mem[100][8] ;
 wire \mem[100][9] ;
 wire \mem[101][0] ;
 wire \mem[101][10] ;
 wire \mem[101][11] ;
 wire \mem[101][12] ;
 wire \mem[101][13] ;
 wire \mem[101][14] ;
 wire \mem[101][15] ;
 wire \mem[101][1] ;
 wire \mem[101][2] ;
 wire \mem[101][3] ;
 wire \mem[101][4] ;
 wire \mem[101][5] ;
 wire \mem[101][6] ;
 wire \mem[101][7] ;
 wire \mem[101][8] ;
 wire \mem[101][9] ;
 wire \mem[102][0] ;
 wire \mem[102][10] ;
 wire \mem[102][11] ;
 wire \mem[102][12] ;
 wire \mem[102][13] ;
 wire \mem[102][14] ;
 wire \mem[102][15] ;
 wire \mem[102][1] ;
 wire \mem[102][2] ;
 wire \mem[102][3] ;
 wire \mem[102][4] ;
 wire \mem[102][5] ;
 wire \mem[102][6] ;
 wire \mem[102][7] ;
 wire \mem[102][8] ;
 wire \mem[102][9] ;
 wire \mem[103][0] ;
 wire \mem[103][10] ;
 wire \mem[103][11] ;
 wire \mem[103][12] ;
 wire \mem[103][13] ;
 wire \mem[103][14] ;
 wire \mem[103][15] ;
 wire \mem[103][1] ;
 wire \mem[103][2] ;
 wire \mem[103][3] ;
 wire \mem[103][4] ;
 wire \mem[103][5] ;
 wire \mem[103][6] ;
 wire \mem[103][7] ;
 wire \mem[103][8] ;
 wire \mem[103][9] ;
 wire \mem[104][0] ;
 wire \mem[104][10] ;
 wire \mem[104][11] ;
 wire \mem[104][12] ;
 wire \mem[104][13] ;
 wire \mem[104][14] ;
 wire \mem[104][15] ;
 wire \mem[104][1] ;
 wire \mem[104][2] ;
 wire \mem[104][3] ;
 wire \mem[104][4] ;
 wire \mem[104][5] ;
 wire \mem[104][6] ;
 wire \mem[104][7] ;
 wire \mem[104][8] ;
 wire \mem[104][9] ;
 wire \mem[105][0] ;
 wire \mem[105][10] ;
 wire \mem[105][11] ;
 wire \mem[105][12] ;
 wire \mem[105][13] ;
 wire \mem[105][14] ;
 wire \mem[105][15] ;
 wire \mem[105][1] ;
 wire \mem[105][2] ;
 wire \mem[105][3] ;
 wire \mem[105][4] ;
 wire \mem[105][5] ;
 wire \mem[105][6] ;
 wire \mem[105][7] ;
 wire \mem[105][8] ;
 wire \mem[105][9] ;
 wire \mem[106][0] ;
 wire \mem[106][10] ;
 wire \mem[106][11] ;
 wire \mem[106][12] ;
 wire \mem[106][13] ;
 wire \mem[106][14] ;
 wire \mem[106][15] ;
 wire \mem[106][1] ;
 wire \mem[106][2] ;
 wire \mem[106][3] ;
 wire \mem[106][4] ;
 wire \mem[106][5] ;
 wire \mem[106][6] ;
 wire \mem[106][7] ;
 wire \mem[106][8] ;
 wire \mem[106][9] ;
 wire \mem[107][0] ;
 wire \mem[107][10] ;
 wire \mem[107][11] ;
 wire \mem[107][12] ;
 wire \mem[107][13] ;
 wire \mem[107][14] ;
 wire \mem[107][15] ;
 wire \mem[107][1] ;
 wire \mem[107][2] ;
 wire \mem[107][3] ;
 wire \mem[107][4] ;
 wire \mem[107][5] ;
 wire \mem[107][6] ;
 wire \mem[107][7] ;
 wire \mem[107][8] ;
 wire \mem[107][9] ;
 wire \mem[108][0] ;
 wire \mem[108][10] ;
 wire \mem[108][11] ;
 wire \mem[108][12] ;
 wire \mem[108][13] ;
 wire \mem[108][14] ;
 wire \mem[108][15] ;
 wire \mem[108][1] ;
 wire \mem[108][2] ;
 wire \mem[108][3] ;
 wire \mem[108][4] ;
 wire \mem[108][5] ;
 wire \mem[108][6] ;
 wire \mem[108][7] ;
 wire \mem[108][8] ;
 wire \mem[108][9] ;
 wire \mem[109][0] ;
 wire \mem[109][10] ;
 wire \mem[109][11] ;
 wire \mem[109][12] ;
 wire \mem[109][13] ;
 wire \mem[109][14] ;
 wire \mem[109][15] ;
 wire \mem[109][1] ;
 wire \mem[109][2] ;
 wire \mem[109][3] ;
 wire \mem[109][4] ;
 wire \mem[109][5] ;
 wire \mem[109][6] ;
 wire \mem[109][7] ;
 wire \mem[109][8] ;
 wire \mem[109][9] ;
 wire \mem[10][0] ;
 wire \mem[10][10] ;
 wire \mem[10][11] ;
 wire \mem[10][12] ;
 wire \mem[10][13] ;
 wire \mem[10][14] ;
 wire \mem[10][15] ;
 wire \mem[10][1] ;
 wire \mem[10][2] ;
 wire \mem[10][3] ;
 wire \mem[10][4] ;
 wire \mem[10][5] ;
 wire \mem[10][6] ;
 wire \mem[10][7] ;
 wire \mem[10][8] ;
 wire \mem[10][9] ;
 wire \mem[110][0] ;
 wire \mem[110][10] ;
 wire \mem[110][11] ;
 wire \mem[110][12] ;
 wire \mem[110][13] ;
 wire \mem[110][14] ;
 wire \mem[110][15] ;
 wire \mem[110][1] ;
 wire \mem[110][2] ;
 wire \mem[110][3] ;
 wire \mem[110][4] ;
 wire \mem[110][5] ;
 wire \mem[110][6] ;
 wire \mem[110][7] ;
 wire \mem[110][8] ;
 wire \mem[110][9] ;
 wire \mem[111][0] ;
 wire \mem[111][10] ;
 wire \mem[111][11] ;
 wire \mem[111][12] ;
 wire \mem[111][13] ;
 wire \mem[111][14] ;
 wire \mem[111][15] ;
 wire \mem[111][1] ;
 wire \mem[111][2] ;
 wire \mem[111][3] ;
 wire \mem[111][4] ;
 wire \mem[111][5] ;
 wire \mem[111][6] ;
 wire \mem[111][7] ;
 wire \mem[111][8] ;
 wire \mem[111][9] ;
 wire \mem[112][0] ;
 wire \mem[112][10] ;
 wire \mem[112][11] ;
 wire \mem[112][12] ;
 wire \mem[112][13] ;
 wire \mem[112][14] ;
 wire \mem[112][15] ;
 wire \mem[112][1] ;
 wire \mem[112][2] ;
 wire \mem[112][3] ;
 wire \mem[112][4] ;
 wire \mem[112][5] ;
 wire \mem[112][6] ;
 wire \mem[112][7] ;
 wire \mem[112][8] ;
 wire \mem[112][9] ;
 wire \mem[113][0] ;
 wire \mem[113][10] ;
 wire \mem[113][11] ;
 wire \mem[113][12] ;
 wire \mem[113][13] ;
 wire \mem[113][14] ;
 wire \mem[113][15] ;
 wire \mem[113][1] ;
 wire \mem[113][2] ;
 wire \mem[113][3] ;
 wire \mem[113][4] ;
 wire \mem[113][5] ;
 wire \mem[113][6] ;
 wire \mem[113][7] ;
 wire \mem[113][8] ;
 wire \mem[113][9] ;
 wire \mem[114][0] ;
 wire \mem[114][10] ;
 wire \mem[114][11] ;
 wire \mem[114][12] ;
 wire \mem[114][13] ;
 wire \mem[114][14] ;
 wire \mem[114][15] ;
 wire \mem[114][1] ;
 wire \mem[114][2] ;
 wire \mem[114][3] ;
 wire \mem[114][4] ;
 wire \mem[114][5] ;
 wire \mem[114][6] ;
 wire \mem[114][7] ;
 wire \mem[114][8] ;
 wire \mem[114][9] ;
 wire \mem[115][0] ;
 wire \mem[115][10] ;
 wire \mem[115][11] ;
 wire \mem[115][12] ;
 wire \mem[115][13] ;
 wire \mem[115][14] ;
 wire \mem[115][15] ;
 wire \mem[115][1] ;
 wire \mem[115][2] ;
 wire \mem[115][3] ;
 wire \mem[115][4] ;
 wire \mem[115][5] ;
 wire \mem[115][6] ;
 wire \mem[115][7] ;
 wire \mem[115][8] ;
 wire \mem[115][9] ;
 wire \mem[116][0] ;
 wire \mem[116][10] ;
 wire \mem[116][11] ;
 wire \mem[116][12] ;
 wire \mem[116][13] ;
 wire \mem[116][14] ;
 wire \mem[116][15] ;
 wire \mem[116][1] ;
 wire \mem[116][2] ;
 wire \mem[116][3] ;
 wire \mem[116][4] ;
 wire \mem[116][5] ;
 wire \mem[116][6] ;
 wire \mem[116][7] ;
 wire \mem[116][8] ;
 wire \mem[116][9] ;
 wire \mem[117][0] ;
 wire \mem[117][10] ;
 wire \mem[117][11] ;
 wire \mem[117][12] ;
 wire \mem[117][13] ;
 wire \mem[117][14] ;
 wire \mem[117][15] ;
 wire \mem[117][1] ;
 wire \mem[117][2] ;
 wire \mem[117][3] ;
 wire \mem[117][4] ;
 wire \mem[117][5] ;
 wire \mem[117][6] ;
 wire \mem[117][7] ;
 wire \mem[117][8] ;
 wire \mem[117][9] ;
 wire \mem[118][0] ;
 wire \mem[118][10] ;
 wire \mem[118][11] ;
 wire \mem[118][12] ;
 wire \mem[118][13] ;
 wire \mem[118][14] ;
 wire \mem[118][15] ;
 wire \mem[118][1] ;
 wire \mem[118][2] ;
 wire \mem[118][3] ;
 wire \mem[118][4] ;
 wire \mem[118][5] ;
 wire \mem[118][6] ;
 wire \mem[118][7] ;
 wire \mem[118][8] ;
 wire \mem[118][9] ;
 wire \mem[119][0] ;
 wire \mem[119][10] ;
 wire \mem[119][11] ;
 wire \mem[119][12] ;
 wire \mem[119][13] ;
 wire \mem[119][14] ;
 wire \mem[119][15] ;
 wire \mem[119][1] ;
 wire \mem[119][2] ;
 wire \mem[119][3] ;
 wire \mem[119][4] ;
 wire \mem[119][5] ;
 wire \mem[119][6] ;
 wire \mem[119][7] ;
 wire \mem[119][8] ;
 wire \mem[119][9] ;
 wire \mem[11][0] ;
 wire \mem[11][10] ;
 wire \mem[11][11] ;
 wire \mem[11][12] ;
 wire \mem[11][13] ;
 wire \mem[11][14] ;
 wire \mem[11][15] ;
 wire \mem[11][1] ;
 wire \mem[11][2] ;
 wire \mem[11][3] ;
 wire \mem[11][4] ;
 wire \mem[11][5] ;
 wire \mem[11][6] ;
 wire \mem[11][7] ;
 wire \mem[11][8] ;
 wire \mem[11][9] ;
 wire \mem[120][0] ;
 wire \mem[120][10] ;
 wire \mem[120][11] ;
 wire \mem[120][12] ;
 wire \mem[120][13] ;
 wire \mem[120][14] ;
 wire \mem[120][15] ;
 wire \mem[120][1] ;
 wire \mem[120][2] ;
 wire \mem[120][3] ;
 wire \mem[120][4] ;
 wire \mem[120][5] ;
 wire \mem[120][6] ;
 wire \mem[120][7] ;
 wire \mem[120][8] ;
 wire \mem[120][9] ;
 wire \mem[121][0] ;
 wire \mem[121][10] ;
 wire \mem[121][11] ;
 wire \mem[121][12] ;
 wire \mem[121][13] ;
 wire \mem[121][14] ;
 wire \mem[121][15] ;
 wire \mem[121][1] ;
 wire \mem[121][2] ;
 wire \mem[121][3] ;
 wire \mem[121][4] ;
 wire \mem[121][5] ;
 wire \mem[121][6] ;
 wire \mem[121][7] ;
 wire \mem[121][8] ;
 wire \mem[121][9] ;
 wire \mem[122][0] ;
 wire \mem[122][10] ;
 wire \mem[122][11] ;
 wire \mem[122][12] ;
 wire \mem[122][13] ;
 wire \mem[122][14] ;
 wire \mem[122][15] ;
 wire \mem[122][1] ;
 wire \mem[122][2] ;
 wire \mem[122][3] ;
 wire \mem[122][4] ;
 wire \mem[122][5] ;
 wire \mem[122][6] ;
 wire \mem[122][7] ;
 wire \mem[122][8] ;
 wire \mem[122][9] ;
 wire \mem[123][0] ;
 wire \mem[123][10] ;
 wire \mem[123][11] ;
 wire \mem[123][12] ;
 wire \mem[123][13] ;
 wire \mem[123][14] ;
 wire \mem[123][15] ;
 wire \mem[123][1] ;
 wire \mem[123][2] ;
 wire \mem[123][3] ;
 wire \mem[123][4] ;
 wire \mem[123][5] ;
 wire \mem[123][6] ;
 wire \mem[123][7] ;
 wire \mem[123][8] ;
 wire \mem[123][9] ;
 wire \mem[124][0] ;
 wire \mem[124][10] ;
 wire \mem[124][11] ;
 wire \mem[124][12] ;
 wire \mem[124][13] ;
 wire \mem[124][14] ;
 wire \mem[124][15] ;
 wire \mem[124][1] ;
 wire \mem[124][2] ;
 wire \mem[124][3] ;
 wire \mem[124][4] ;
 wire \mem[124][5] ;
 wire \mem[124][6] ;
 wire \mem[124][7] ;
 wire \mem[124][8] ;
 wire \mem[124][9] ;
 wire \mem[125][0] ;
 wire \mem[125][10] ;
 wire \mem[125][11] ;
 wire \mem[125][12] ;
 wire \mem[125][13] ;
 wire \mem[125][14] ;
 wire \mem[125][15] ;
 wire \mem[125][1] ;
 wire \mem[125][2] ;
 wire \mem[125][3] ;
 wire \mem[125][4] ;
 wire \mem[125][5] ;
 wire \mem[125][6] ;
 wire \mem[125][7] ;
 wire \mem[125][8] ;
 wire \mem[125][9] ;
 wire \mem[126][0] ;
 wire \mem[126][10] ;
 wire \mem[126][11] ;
 wire \mem[126][12] ;
 wire \mem[126][13] ;
 wire \mem[126][14] ;
 wire \mem[126][15] ;
 wire \mem[126][1] ;
 wire \mem[126][2] ;
 wire \mem[126][3] ;
 wire \mem[126][4] ;
 wire \mem[126][5] ;
 wire \mem[126][6] ;
 wire \mem[126][7] ;
 wire \mem[126][8] ;
 wire \mem[126][9] ;
 wire \mem[127][0] ;
 wire \mem[127][10] ;
 wire \mem[127][11] ;
 wire \mem[127][12] ;
 wire \mem[127][13] ;
 wire \mem[127][14] ;
 wire \mem[127][15] ;
 wire \mem[127][1] ;
 wire \mem[127][2] ;
 wire \mem[127][3] ;
 wire \mem[127][4] ;
 wire \mem[127][5] ;
 wire \mem[127][6] ;
 wire \mem[127][7] ;
 wire \mem[127][8] ;
 wire \mem[127][9] ;
 wire \mem[12][0] ;
 wire \mem[12][10] ;
 wire \mem[12][11] ;
 wire \mem[12][12] ;
 wire \mem[12][13] ;
 wire \mem[12][14] ;
 wire \mem[12][15] ;
 wire \mem[12][1] ;
 wire \mem[12][2] ;
 wire \mem[12][3] ;
 wire \mem[12][4] ;
 wire \mem[12][5] ;
 wire \mem[12][6] ;
 wire \mem[12][7] ;
 wire \mem[12][8] ;
 wire \mem[12][9] ;
 wire \mem[13][0] ;
 wire \mem[13][10] ;
 wire \mem[13][11] ;
 wire \mem[13][12] ;
 wire \mem[13][13] ;
 wire \mem[13][14] ;
 wire \mem[13][15] ;
 wire \mem[13][1] ;
 wire \mem[13][2] ;
 wire \mem[13][3] ;
 wire \mem[13][4] ;
 wire \mem[13][5] ;
 wire \mem[13][6] ;
 wire \mem[13][7] ;
 wire \mem[13][8] ;
 wire \mem[13][9] ;
 wire \mem[14][0] ;
 wire \mem[14][10] ;
 wire \mem[14][11] ;
 wire \mem[14][12] ;
 wire \mem[14][13] ;
 wire \mem[14][14] ;
 wire \mem[14][15] ;
 wire \mem[14][1] ;
 wire \mem[14][2] ;
 wire \mem[14][3] ;
 wire \mem[14][4] ;
 wire \mem[14][5] ;
 wire \mem[14][6] ;
 wire \mem[14][7] ;
 wire \mem[14][8] ;
 wire \mem[14][9] ;
 wire \mem[15][0] ;
 wire \mem[15][10] ;
 wire \mem[15][11] ;
 wire \mem[15][12] ;
 wire \mem[15][13] ;
 wire \mem[15][14] ;
 wire \mem[15][15] ;
 wire \mem[15][1] ;
 wire \mem[15][2] ;
 wire \mem[15][3] ;
 wire \mem[15][4] ;
 wire \mem[15][5] ;
 wire \mem[15][6] ;
 wire \mem[15][7] ;
 wire \mem[15][8] ;
 wire \mem[15][9] ;
 wire \mem[16][0] ;
 wire \mem[16][10] ;
 wire \mem[16][11] ;
 wire \mem[16][12] ;
 wire \mem[16][13] ;
 wire \mem[16][14] ;
 wire \mem[16][15] ;
 wire \mem[16][1] ;
 wire \mem[16][2] ;
 wire \mem[16][3] ;
 wire \mem[16][4] ;
 wire \mem[16][5] ;
 wire \mem[16][6] ;
 wire \mem[16][7] ;
 wire \mem[16][8] ;
 wire \mem[16][9] ;
 wire \mem[17][0] ;
 wire \mem[17][10] ;
 wire \mem[17][11] ;
 wire \mem[17][12] ;
 wire \mem[17][13] ;
 wire \mem[17][14] ;
 wire \mem[17][15] ;
 wire \mem[17][1] ;
 wire \mem[17][2] ;
 wire \mem[17][3] ;
 wire \mem[17][4] ;
 wire \mem[17][5] ;
 wire \mem[17][6] ;
 wire \mem[17][7] ;
 wire \mem[17][8] ;
 wire \mem[17][9] ;
 wire \mem[18][0] ;
 wire \mem[18][10] ;
 wire \mem[18][11] ;
 wire \mem[18][12] ;
 wire \mem[18][13] ;
 wire \mem[18][14] ;
 wire \mem[18][15] ;
 wire \mem[18][1] ;
 wire \mem[18][2] ;
 wire \mem[18][3] ;
 wire \mem[18][4] ;
 wire \mem[18][5] ;
 wire \mem[18][6] ;
 wire \mem[18][7] ;
 wire \mem[18][8] ;
 wire \mem[18][9] ;
 wire \mem[19][0] ;
 wire \mem[19][10] ;
 wire \mem[19][11] ;
 wire \mem[19][12] ;
 wire \mem[19][13] ;
 wire \mem[19][14] ;
 wire \mem[19][15] ;
 wire \mem[19][1] ;
 wire \mem[19][2] ;
 wire \mem[19][3] ;
 wire \mem[19][4] ;
 wire \mem[19][5] ;
 wire \mem[19][6] ;
 wire \mem[19][7] ;
 wire \mem[19][8] ;
 wire \mem[19][9] ;
 wire \mem[1][0] ;
 wire \mem[1][10] ;
 wire \mem[1][11] ;
 wire \mem[1][12] ;
 wire \mem[1][13] ;
 wire \mem[1][14] ;
 wire \mem[1][15] ;
 wire \mem[1][1] ;
 wire \mem[1][2] ;
 wire \mem[1][3] ;
 wire \mem[1][4] ;
 wire \mem[1][5] ;
 wire \mem[1][6] ;
 wire \mem[1][7] ;
 wire \mem[1][8] ;
 wire \mem[1][9] ;
 wire \mem[20][0] ;
 wire \mem[20][10] ;
 wire \mem[20][11] ;
 wire \mem[20][12] ;
 wire \mem[20][13] ;
 wire \mem[20][14] ;
 wire \mem[20][15] ;
 wire \mem[20][1] ;
 wire \mem[20][2] ;
 wire \mem[20][3] ;
 wire \mem[20][4] ;
 wire \mem[20][5] ;
 wire \mem[20][6] ;
 wire \mem[20][7] ;
 wire \mem[20][8] ;
 wire \mem[20][9] ;
 wire \mem[21][0] ;
 wire \mem[21][10] ;
 wire \mem[21][11] ;
 wire \mem[21][12] ;
 wire \mem[21][13] ;
 wire \mem[21][14] ;
 wire \mem[21][15] ;
 wire \mem[21][1] ;
 wire \mem[21][2] ;
 wire \mem[21][3] ;
 wire \mem[21][4] ;
 wire \mem[21][5] ;
 wire \mem[21][6] ;
 wire \mem[21][7] ;
 wire \mem[21][8] ;
 wire \mem[21][9] ;
 wire \mem[22][0] ;
 wire \mem[22][10] ;
 wire \mem[22][11] ;
 wire \mem[22][12] ;
 wire \mem[22][13] ;
 wire \mem[22][14] ;
 wire \mem[22][15] ;
 wire \mem[22][1] ;
 wire \mem[22][2] ;
 wire \mem[22][3] ;
 wire \mem[22][4] ;
 wire \mem[22][5] ;
 wire \mem[22][6] ;
 wire \mem[22][7] ;
 wire \mem[22][8] ;
 wire \mem[22][9] ;
 wire \mem[23][0] ;
 wire \mem[23][10] ;
 wire \mem[23][11] ;
 wire \mem[23][12] ;
 wire \mem[23][13] ;
 wire \mem[23][14] ;
 wire \mem[23][15] ;
 wire \mem[23][1] ;
 wire \mem[23][2] ;
 wire \mem[23][3] ;
 wire \mem[23][4] ;
 wire \mem[23][5] ;
 wire \mem[23][6] ;
 wire \mem[23][7] ;
 wire \mem[23][8] ;
 wire \mem[23][9] ;
 wire \mem[24][0] ;
 wire \mem[24][10] ;
 wire \mem[24][11] ;
 wire \mem[24][12] ;
 wire \mem[24][13] ;
 wire \mem[24][14] ;
 wire \mem[24][15] ;
 wire \mem[24][1] ;
 wire \mem[24][2] ;
 wire \mem[24][3] ;
 wire \mem[24][4] ;
 wire \mem[24][5] ;
 wire \mem[24][6] ;
 wire \mem[24][7] ;
 wire \mem[24][8] ;
 wire \mem[24][9] ;
 wire \mem[25][0] ;
 wire \mem[25][10] ;
 wire \mem[25][11] ;
 wire \mem[25][12] ;
 wire \mem[25][13] ;
 wire \mem[25][14] ;
 wire \mem[25][15] ;
 wire \mem[25][1] ;
 wire \mem[25][2] ;
 wire \mem[25][3] ;
 wire \mem[25][4] ;
 wire \mem[25][5] ;
 wire \mem[25][6] ;
 wire \mem[25][7] ;
 wire \mem[25][8] ;
 wire \mem[25][9] ;
 wire \mem[26][0] ;
 wire \mem[26][10] ;
 wire \mem[26][11] ;
 wire \mem[26][12] ;
 wire \mem[26][13] ;
 wire \mem[26][14] ;
 wire \mem[26][15] ;
 wire \mem[26][1] ;
 wire \mem[26][2] ;
 wire \mem[26][3] ;
 wire \mem[26][4] ;
 wire \mem[26][5] ;
 wire \mem[26][6] ;
 wire \mem[26][7] ;
 wire \mem[26][8] ;
 wire \mem[26][9] ;
 wire \mem[27][0] ;
 wire \mem[27][10] ;
 wire \mem[27][11] ;
 wire \mem[27][12] ;
 wire \mem[27][13] ;
 wire \mem[27][14] ;
 wire \mem[27][15] ;
 wire \mem[27][1] ;
 wire \mem[27][2] ;
 wire \mem[27][3] ;
 wire \mem[27][4] ;
 wire \mem[27][5] ;
 wire \mem[27][6] ;
 wire \mem[27][7] ;
 wire \mem[27][8] ;
 wire \mem[27][9] ;
 wire \mem[28][0] ;
 wire \mem[28][10] ;
 wire \mem[28][11] ;
 wire \mem[28][12] ;
 wire \mem[28][13] ;
 wire \mem[28][14] ;
 wire \mem[28][15] ;
 wire \mem[28][1] ;
 wire \mem[28][2] ;
 wire \mem[28][3] ;
 wire \mem[28][4] ;
 wire \mem[28][5] ;
 wire \mem[28][6] ;
 wire \mem[28][7] ;
 wire \mem[28][8] ;
 wire \mem[28][9] ;
 wire \mem[29][0] ;
 wire \mem[29][10] ;
 wire \mem[29][11] ;
 wire \mem[29][12] ;
 wire \mem[29][13] ;
 wire \mem[29][14] ;
 wire \mem[29][15] ;
 wire \mem[29][1] ;
 wire \mem[29][2] ;
 wire \mem[29][3] ;
 wire \mem[29][4] ;
 wire \mem[29][5] ;
 wire \mem[29][6] ;
 wire \mem[29][7] ;
 wire \mem[29][8] ;
 wire \mem[29][9] ;
 wire \mem[2][0] ;
 wire \mem[2][10] ;
 wire \mem[2][11] ;
 wire \mem[2][12] ;
 wire \mem[2][13] ;
 wire \mem[2][14] ;
 wire \mem[2][15] ;
 wire \mem[2][1] ;
 wire \mem[2][2] ;
 wire \mem[2][3] ;
 wire \mem[2][4] ;
 wire \mem[2][5] ;
 wire \mem[2][6] ;
 wire \mem[2][7] ;
 wire \mem[2][8] ;
 wire \mem[2][9] ;
 wire \mem[30][0] ;
 wire \mem[30][10] ;
 wire \mem[30][11] ;
 wire \mem[30][12] ;
 wire \mem[30][13] ;
 wire \mem[30][14] ;
 wire \mem[30][15] ;
 wire \mem[30][1] ;
 wire \mem[30][2] ;
 wire \mem[30][3] ;
 wire \mem[30][4] ;
 wire \mem[30][5] ;
 wire \mem[30][6] ;
 wire \mem[30][7] ;
 wire \mem[30][8] ;
 wire \mem[30][9] ;
 wire \mem[31][0] ;
 wire \mem[31][10] ;
 wire \mem[31][11] ;
 wire \mem[31][12] ;
 wire \mem[31][13] ;
 wire \mem[31][14] ;
 wire \mem[31][15] ;
 wire \mem[31][1] ;
 wire \mem[31][2] ;
 wire \mem[31][3] ;
 wire \mem[31][4] ;
 wire \mem[31][5] ;
 wire \mem[31][6] ;
 wire \mem[31][7] ;
 wire \mem[31][8] ;
 wire \mem[31][9] ;
 wire \mem[32][0] ;
 wire \mem[32][10] ;
 wire \mem[32][11] ;
 wire \mem[32][12] ;
 wire \mem[32][13] ;
 wire \mem[32][14] ;
 wire \mem[32][15] ;
 wire \mem[32][1] ;
 wire \mem[32][2] ;
 wire \mem[32][3] ;
 wire \mem[32][4] ;
 wire \mem[32][5] ;
 wire \mem[32][6] ;
 wire \mem[32][7] ;
 wire \mem[32][8] ;
 wire \mem[32][9] ;
 wire \mem[33][0] ;
 wire \mem[33][10] ;
 wire \mem[33][11] ;
 wire \mem[33][12] ;
 wire \mem[33][13] ;
 wire \mem[33][14] ;
 wire \mem[33][15] ;
 wire \mem[33][1] ;
 wire \mem[33][2] ;
 wire \mem[33][3] ;
 wire \mem[33][4] ;
 wire \mem[33][5] ;
 wire \mem[33][6] ;
 wire \mem[33][7] ;
 wire \mem[33][8] ;
 wire \mem[33][9] ;
 wire \mem[34][0] ;
 wire \mem[34][10] ;
 wire \mem[34][11] ;
 wire \mem[34][12] ;
 wire \mem[34][13] ;
 wire \mem[34][14] ;
 wire \mem[34][15] ;
 wire \mem[34][1] ;
 wire \mem[34][2] ;
 wire \mem[34][3] ;
 wire \mem[34][4] ;
 wire \mem[34][5] ;
 wire \mem[34][6] ;
 wire \mem[34][7] ;
 wire \mem[34][8] ;
 wire \mem[34][9] ;
 wire \mem[35][0] ;
 wire \mem[35][10] ;
 wire \mem[35][11] ;
 wire \mem[35][12] ;
 wire \mem[35][13] ;
 wire \mem[35][14] ;
 wire \mem[35][15] ;
 wire \mem[35][1] ;
 wire \mem[35][2] ;
 wire \mem[35][3] ;
 wire \mem[35][4] ;
 wire \mem[35][5] ;
 wire \mem[35][6] ;
 wire \mem[35][7] ;
 wire \mem[35][8] ;
 wire \mem[35][9] ;
 wire \mem[36][0] ;
 wire \mem[36][10] ;
 wire \mem[36][11] ;
 wire \mem[36][12] ;
 wire \mem[36][13] ;
 wire \mem[36][14] ;
 wire \mem[36][15] ;
 wire \mem[36][1] ;
 wire \mem[36][2] ;
 wire \mem[36][3] ;
 wire \mem[36][4] ;
 wire \mem[36][5] ;
 wire \mem[36][6] ;
 wire \mem[36][7] ;
 wire \mem[36][8] ;
 wire \mem[36][9] ;
 wire \mem[37][0] ;
 wire \mem[37][10] ;
 wire \mem[37][11] ;
 wire \mem[37][12] ;
 wire \mem[37][13] ;
 wire \mem[37][14] ;
 wire \mem[37][15] ;
 wire \mem[37][1] ;
 wire \mem[37][2] ;
 wire \mem[37][3] ;
 wire \mem[37][4] ;
 wire \mem[37][5] ;
 wire \mem[37][6] ;
 wire \mem[37][7] ;
 wire \mem[37][8] ;
 wire \mem[37][9] ;
 wire \mem[38][0] ;
 wire \mem[38][10] ;
 wire \mem[38][11] ;
 wire \mem[38][12] ;
 wire \mem[38][13] ;
 wire \mem[38][14] ;
 wire \mem[38][15] ;
 wire \mem[38][1] ;
 wire \mem[38][2] ;
 wire \mem[38][3] ;
 wire \mem[38][4] ;
 wire \mem[38][5] ;
 wire \mem[38][6] ;
 wire \mem[38][7] ;
 wire \mem[38][8] ;
 wire \mem[38][9] ;
 wire \mem[39][0] ;
 wire \mem[39][10] ;
 wire \mem[39][11] ;
 wire \mem[39][12] ;
 wire \mem[39][13] ;
 wire \mem[39][14] ;
 wire \mem[39][15] ;
 wire \mem[39][1] ;
 wire \mem[39][2] ;
 wire \mem[39][3] ;
 wire \mem[39][4] ;
 wire \mem[39][5] ;
 wire \mem[39][6] ;
 wire \mem[39][7] ;
 wire \mem[39][8] ;
 wire \mem[39][9] ;
 wire \mem[3][0] ;
 wire \mem[3][10] ;
 wire \mem[3][11] ;
 wire \mem[3][12] ;
 wire \mem[3][13] ;
 wire \mem[3][14] ;
 wire \mem[3][15] ;
 wire \mem[3][1] ;
 wire \mem[3][2] ;
 wire \mem[3][3] ;
 wire \mem[3][4] ;
 wire \mem[3][5] ;
 wire \mem[3][6] ;
 wire \mem[3][7] ;
 wire \mem[3][8] ;
 wire \mem[3][9] ;
 wire \mem[40][0] ;
 wire \mem[40][10] ;
 wire \mem[40][11] ;
 wire \mem[40][12] ;
 wire \mem[40][13] ;
 wire \mem[40][14] ;
 wire \mem[40][15] ;
 wire \mem[40][1] ;
 wire \mem[40][2] ;
 wire \mem[40][3] ;
 wire \mem[40][4] ;
 wire \mem[40][5] ;
 wire \mem[40][6] ;
 wire \mem[40][7] ;
 wire \mem[40][8] ;
 wire \mem[40][9] ;
 wire \mem[41][0] ;
 wire \mem[41][10] ;
 wire \mem[41][11] ;
 wire \mem[41][12] ;
 wire \mem[41][13] ;
 wire \mem[41][14] ;
 wire \mem[41][15] ;
 wire \mem[41][1] ;
 wire \mem[41][2] ;
 wire \mem[41][3] ;
 wire \mem[41][4] ;
 wire \mem[41][5] ;
 wire \mem[41][6] ;
 wire \mem[41][7] ;
 wire \mem[41][8] ;
 wire \mem[41][9] ;
 wire \mem[42][0] ;
 wire \mem[42][10] ;
 wire \mem[42][11] ;
 wire \mem[42][12] ;
 wire \mem[42][13] ;
 wire \mem[42][14] ;
 wire \mem[42][15] ;
 wire \mem[42][1] ;
 wire \mem[42][2] ;
 wire \mem[42][3] ;
 wire \mem[42][4] ;
 wire \mem[42][5] ;
 wire \mem[42][6] ;
 wire \mem[42][7] ;
 wire \mem[42][8] ;
 wire \mem[42][9] ;
 wire \mem[43][0] ;
 wire \mem[43][10] ;
 wire \mem[43][11] ;
 wire \mem[43][12] ;
 wire \mem[43][13] ;
 wire \mem[43][14] ;
 wire \mem[43][15] ;
 wire \mem[43][1] ;
 wire \mem[43][2] ;
 wire \mem[43][3] ;
 wire \mem[43][4] ;
 wire \mem[43][5] ;
 wire \mem[43][6] ;
 wire \mem[43][7] ;
 wire \mem[43][8] ;
 wire \mem[43][9] ;
 wire \mem[44][0] ;
 wire \mem[44][10] ;
 wire \mem[44][11] ;
 wire \mem[44][12] ;
 wire \mem[44][13] ;
 wire \mem[44][14] ;
 wire \mem[44][15] ;
 wire \mem[44][1] ;
 wire \mem[44][2] ;
 wire \mem[44][3] ;
 wire \mem[44][4] ;
 wire \mem[44][5] ;
 wire \mem[44][6] ;
 wire \mem[44][7] ;
 wire \mem[44][8] ;
 wire \mem[44][9] ;
 wire \mem[45][0] ;
 wire \mem[45][10] ;
 wire \mem[45][11] ;
 wire \mem[45][12] ;
 wire \mem[45][13] ;
 wire \mem[45][14] ;
 wire \mem[45][15] ;
 wire \mem[45][1] ;
 wire \mem[45][2] ;
 wire \mem[45][3] ;
 wire \mem[45][4] ;
 wire \mem[45][5] ;
 wire \mem[45][6] ;
 wire \mem[45][7] ;
 wire \mem[45][8] ;
 wire \mem[45][9] ;
 wire \mem[46][0] ;
 wire \mem[46][10] ;
 wire \mem[46][11] ;
 wire \mem[46][12] ;
 wire \mem[46][13] ;
 wire \mem[46][14] ;
 wire \mem[46][15] ;
 wire \mem[46][1] ;
 wire \mem[46][2] ;
 wire \mem[46][3] ;
 wire \mem[46][4] ;
 wire \mem[46][5] ;
 wire \mem[46][6] ;
 wire \mem[46][7] ;
 wire \mem[46][8] ;
 wire \mem[46][9] ;
 wire \mem[47][0] ;
 wire \mem[47][10] ;
 wire \mem[47][11] ;
 wire \mem[47][12] ;
 wire \mem[47][13] ;
 wire \mem[47][14] ;
 wire \mem[47][15] ;
 wire \mem[47][1] ;
 wire \mem[47][2] ;
 wire \mem[47][3] ;
 wire \mem[47][4] ;
 wire \mem[47][5] ;
 wire \mem[47][6] ;
 wire \mem[47][7] ;
 wire \mem[47][8] ;
 wire \mem[47][9] ;
 wire \mem[48][0] ;
 wire \mem[48][10] ;
 wire \mem[48][11] ;
 wire \mem[48][12] ;
 wire \mem[48][13] ;
 wire \mem[48][14] ;
 wire \mem[48][15] ;
 wire \mem[48][1] ;
 wire \mem[48][2] ;
 wire \mem[48][3] ;
 wire \mem[48][4] ;
 wire \mem[48][5] ;
 wire \mem[48][6] ;
 wire \mem[48][7] ;
 wire \mem[48][8] ;
 wire \mem[48][9] ;
 wire \mem[49][0] ;
 wire \mem[49][10] ;
 wire \mem[49][11] ;
 wire \mem[49][12] ;
 wire \mem[49][13] ;
 wire \mem[49][14] ;
 wire \mem[49][15] ;
 wire \mem[49][1] ;
 wire \mem[49][2] ;
 wire \mem[49][3] ;
 wire \mem[49][4] ;
 wire \mem[49][5] ;
 wire \mem[49][6] ;
 wire \mem[49][7] ;
 wire \mem[49][8] ;
 wire \mem[49][9] ;
 wire \mem[4][0] ;
 wire \mem[4][10] ;
 wire \mem[4][11] ;
 wire \mem[4][12] ;
 wire \mem[4][13] ;
 wire \mem[4][14] ;
 wire \mem[4][15] ;
 wire \mem[4][1] ;
 wire \mem[4][2] ;
 wire \mem[4][3] ;
 wire \mem[4][4] ;
 wire \mem[4][5] ;
 wire \mem[4][6] ;
 wire \mem[4][7] ;
 wire \mem[4][8] ;
 wire \mem[4][9] ;
 wire \mem[50][0] ;
 wire \mem[50][10] ;
 wire \mem[50][11] ;
 wire \mem[50][12] ;
 wire \mem[50][13] ;
 wire \mem[50][14] ;
 wire \mem[50][15] ;
 wire \mem[50][1] ;
 wire \mem[50][2] ;
 wire \mem[50][3] ;
 wire \mem[50][4] ;
 wire \mem[50][5] ;
 wire \mem[50][6] ;
 wire \mem[50][7] ;
 wire \mem[50][8] ;
 wire \mem[50][9] ;
 wire \mem[51][0] ;
 wire \mem[51][10] ;
 wire \mem[51][11] ;
 wire \mem[51][12] ;
 wire \mem[51][13] ;
 wire \mem[51][14] ;
 wire \mem[51][15] ;
 wire \mem[51][1] ;
 wire \mem[51][2] ;
 wire \mem[51][3] ;
 wire \mem[51][4] ;
 wire \mem[51][5] ;
 wire \mem[51][6] ;
 wire \mem[51][7] ;
 wire \mem[51][8] ;
 wire \mem[51][9] ;
 wire \mem[52][0] ;
 wire \mem[52][10] ;
 wire \mem[52][11] ;
 wire \mem[52][12] ;
 wire \mem[52][13] ;
 wire \mem[52][14] ;
 wire \mem[52][15] ;
 wire \mem[52][1] ;
 wire \mem[52][2] ;
 wire \mem[52][3] ;
 wire \mem[52][4] ;
 wire \mem[52][5] ;
 wire \mem[52][6] ;
 wire \mem[52][7] ;
 wire \mem[52][8] ;
 wire \mem[52][9] ;
 wire \mem[53][0] ;
 wire \mem[53][10] ;
 wire \mem[53][11] ;
 wire \mem[53][12] ;
 wire \mem[53][13] ;
 wire \mem[53][14] ;
 wire \mem[53][15] ;
 wire \mem[53][1] ;
 wire \mem[53][2] ;
 wire \mem[53][3] ;
 wire \mem[53][4] ;
 wire \mem[53][5] ;
 wire \mem[53][6] ;
 wire \mem[53][7] ;
 wire \mem[53][8] ;
 wire \mem[53][9] ;
 wire \mem[54][0] ;
 wire \mem[54][10] ;
 wire \mem[54][11] ;
 wire \mem[54][12] ;
 wire \mem[54][13] ;
 wire \mem[54][14] ;
 wire \mem[54][15] ;
 wire \mem[54][1] ;
 wire \mem[54][2] ;
 wire \mem[54][3] ;
 wire \mem[54][4] ;
 wire \mem[54][5] ;
 wire \mem[54][6] ;
 wire \mem[54][7] ;
 wire \mem[54][8] ;
 wire \mem[54][9] ;
 wire \mem[55][0] ;
 wire \mem[55][10] ;
 wire \mem[55][11] ;
 wire \mem[55][12] ;
 wire \mem[55][13] ;
 wire \mem[55][14] ;
 wire \mem[55][15] ;
 wire \mem[55][1] ;
 wire \mem[55][2] ;
 wire \mem[55][3] ;
 wire \mem[55][4] ;
 wire \mem[55][5] ;
 wire \mem[55][6] ;
 wire \mem[55][7] ;
 wire \mem[55][8] ;
 wire \mem[55][9] ;
 wire \mem[56][0] ;
 wire \mem[56][10] ;
 wire \mem[56][11] ;
 wire \mem[56][12] ;
 wire \mem[56][13] ;
 wire \mem[56][14] ;
 wire \mem[56][15] ;
 wire \mem[56][1] ;
 wire \mem[56][2] ;
 wire \mem[56][3] ;
 wire \mem[56][4] ;
 wire \mem[56][5] ;
 wire \mem[56][6] ;
 wire \mem[56][7] ;
 wire \mem[56][8] ;
 wire \mem[56][9] ;
 wire \mem[57][0] ;
 wire \mem[57][10] ;
 wire \mem[57][11] ;
 wire \mem[57][12] ;
 wire \mem[57][13] ;
 wire \mem[57][14] ;
 wire \mem[57][15] ;
 wire \mem[57][1] ;
 wire \mem[57][2] ;
 wire \mem[57][3] ;
 wire \mem[57][4] ;
 wire \mem[57][5] ;
 wire \mem[57][6] ;
 wire \mem[57][7] ;
 wire \mem[57][8] ;
 wire \mem[57][9] ;
 wire \mem[58][0] ;
 wire \mem[58][10] ;
 wire \mem[58][11] ;
 wire \mem[58][12] ;
 wire \mem[58][13] ;
 wire \mem[58][14] ;
 wire \mem[58][15] ;
 wire \mem[58][1] ;
 wire \mem[58][2] ;
 wire \mem[58][3] ;
 wire \mem[58][4] ;
 wire \mem[58][5] ;
 wire \mem[58][6] ;
 wire \mem[58][7] ;
 wire \mem[58][8] ;
 wire \mem[58][9] ;
 wire \mem[59][0] ;
 wire \mem[59][10] ;
 wire \mem[59][11] ;
 wire \mem[59][12] ;
 wire \mem[59][13] ;
 wire \mem[59][14] ;
 wire \mem[59][15] ;
 wire \mem[59][1] ;
 wire \mem[59][2] ;
 wire \mem[59][3] ;
 wire \mem[59][4] ;
 wire \mem[59][5] ;
 wire \mem[59][6] ;
 wire \mem[59][7] ;
 wire \mem[59][8] ;
 wire \mem[59][9] ;
 wire \mem[5][0] ;
 wire \mem[5][10] ;
 wire \mem[5][11] ;
 wire \mem[5][12] ;
 wire \mem[5][13] ;
 wire \mem[5][14] ;
 wire \mem[5][15] ;
 wire \mem[5][1] ;
 wire \mem[5][2] ;
 wire \mem[5][3] ;
 wire \mem[5][4] ;
 wire \mem[5][5] ;
 wire \mem[5][6] ;
 wire \mem[5][7] ;
 wire \mem[5][8] ;
 wire \mem[5][9] ;
 wire \mem[60][0] ;
 wire \mem[60][10] ;
 wire \mem[60][11] ;
 wire \mem[60][12] ;
 wire \mem[60][13] ;
 wire \mem[60][14] ;
 wire \mem[60][15] ;
 wire \mem[60][1] ;
 wire \mem[60][2] ;
 wire \mem[60][3] ;
 wire \mem[60][4] ;
 wire \mem[60][5] ;
 wire \mem[60][6] ;
 wire \mem[60][7] ;
 wire \mem[60][8] ;
 wire \mem[60][9] ;
 wire \mem[61][0] ;
 wire \mem[61][10] ;
 wire \mem[61][11] ;
 wire \mem[61][12] ;
 wire \mem[61][13] ;
 wire \mem[61][14] ;
 wire \mem[61][15] ;
 wire \mem[61][1] ;
 wire \mem[61][2] ;
 wire \mem[61][3] ;
 wire \mem[61][4] ;
 wire \mem[61][5] ;
 wire \mem[61][6] ;
 wire \mem[61][7] ;
 wire \mem[61][8] ;
 wire \mem[61][9] ;
 wire \mem[62][0] ;
 wire \mem[62][10] ;
 wire \mem[62][11] ;
 wire \mem[62][12] ;
 wire \mem[62][13] ;
 wire \mem[62][14] ;
 wire \mem[62][15] ;
 wire \mem[62][1] ;
 wire \mem[62][2] ;
 wire \mem[62][3] ;
 wire \mem[62][4] ;
 wire \mem[62][5] ;
 wire \mem[62][6] ;
 wire \mem[62][7] ;
 wire \mem[62][8] ;
 wire \mem[62][9] ;
 wire \mem[63][0] ;
 wire \mem[63][10] ;
 wire \mem[63][11] ;
 wire \mem[63][12] ;
 wire \mem[63][13] ;
 wire \mem[63][14] ;
 wire \mem[63][15] ;
 wire \mem[63][1] ;
 wire \mem[63][2] ;
 wire \mem[63][3] ;
 wire \mem[63][4] ;
 wire \mem[63][5] ;
 wire \mem[63][6] ;
 wire \mem[63][7] ;
 wire \mem[63][8] ;
 wire \mem[63][9] ;
 wire \mem[64][0] ;
 wire \mem[64][10] ;
 wire \mem[64][11] ;
 wire \mem[64][12] ;
 wire \mem[64][13] ;
 wire \mem[64][14] ;
 wire \mem[64][15] ;
 wire \mem[64][1] ;
 wire \mem[64][2] ;
 wire \mem[64][3] ;
 wire \mem[64][4] ;
 wire \mem[64][5] ;
 wire \mem[64][6] ;
 wire \mem[64][7] ;
 wire \mem[64][8] ;
 wire \mem[64][9] ;
 wire \mem[65][0] ;
 wire \mem[65][10] ;
 wire \mem[65][11] ;
 wire \mem[65][12] ;
 wire \mem[65][13] ;
 wire \mem[65][14] ;
 wire \mem[65][15] ;
 wire \mem[65][1] ;
 wire \mem[65][2] ;
 wire \mem[65][3] ;
 wire \mem[65][4] ;
 wire \mem[65][5] ;
 wire \mem[65][6] ;
 wire \mem[65][7] ;
 wire \mem[65][8] ;
 wire \mem[65][9] ;
 wire \mem[66][0] ;
 wire \mem[66][10] ;
 wire \mem[66][11] ;
 wire \mem[66][12] ;
 wire \mem[66][13] ;
 wire \mem[66][14] ;
 wire \mem[66][15] ;
 wire \mem[66][1] ;
 wire \mem[66][2] ;
 wire \mem[66][3] ;
 wire \mem[66][4] ;
 wire \mem[66][5] ;
 wire \mem[66][6] ;
 wire \mem[66][7] ;
 wire \mem[66][8] ;
 wire \mem[66][9] ;
 wire \mem[67][0] ;
 wire \mem[67][10] ;
 wire \mem[67][11] ;
 wire \mem[67][12] ;
 wire \mem[67][13] ;
 wire \mem[67][14] ;
 wire \mem[67][15] ;
 wire \mem[67][1] ;
 wire \mem[67][2] ;
 wire \mem[67][3] ;
 wire \mem[67][4] ;
 wire \mem[67][5] ;
 wire \mem[67][6] ;
 wire \mem[67][7] ;
 wire \mem[67][8] ;
 wire \mem[67][9] ;
 wire \mem[68][0] ;
 wire \mem[68][10] ;
 wire \mem[68][11] ;
 wire \mem[68][12] ;
 wire \mem[68][13] ;
 wire \mem[68][14] ;
 wire \mem[68][15] ;
 wire \mem[68][1] ;
 wire \mem[68][2] ;
 wire \mem[68][3] ;
 wire \mem[68][4] ;
 wire \mem[68][5] ;
 wire \mem[68][6] ;
 wire \mem[68][7] ;
 wire \mem[68][8] ;
 wire \mem[68][9] ;
 wire \mem[69][0] ;
 wire \mem[69][10] ;
 wire \mem[69][11] ;
 wire \mem[69][12] ;
 wire \mem[69][13] ;
 wire \mem[69][14] ;
 wire \mem[69][15] ;
 wire \mem[69][1] ;
 wire \mem[69][2] ;
 wire \mem[69][3] ;
 wire \mem[69][4] ;
 wire \mem[69][5] ;
 wire \mem[69][6] ;
 wire \mem[69][7] ;
 wire \mem[69][8] ;
 wire \mem[69][9] ;
 wire \mem[6][0] ;
 wire \mem[6][10] ;
 wire \mem[6][11] ;
 wire \mem[6][12] ;
 wire \mem[6][13] ;
 wire \mem[6][14] ;
 wire \mem[6][15] ;
 wire \mem[6][1] ;
 wire \mem[6][2] ;
 wire \mem[6][3] ;
 wire \mem[6][4] ;
 wire \mem[6][5] ;
 wire \mem[6][6] ;
 wire \mem[6][7] ;
 wire \mem[6][8] ;
 wire \mem[6][9] ;
 wire \mem[70][0] ;
 wire \mem[70][10] ;
 wire \mem[70][11] ;
 wire \mem[70][12] ;
 wire \mem[70][13] ;
 wire \mem[70][14] ;
 wire \mem[70][15] ;
 wire \mem[70][1] ;
 wire \mem[70][2] ;
 wire \mem[70][3] ;
 wire \mem[70][4] ;
 wire \mem[70][5] ;
 wire \mem[70][6] ;
 wire \mem[70][7] ;
 wire \mem[70][8] ;
 wire \mem[70][9] ;
 wire \mem[71][0] ;
 wire \mem[71][10] ;
 wire \mem[71][11] ;
 wire \mem[71][12] ;
 wire \mem[71][13] ;
 wire \mem[71][14] ;
 wire \mem[71][15] ;
 wire \mem[71][1] ;
 wire \mem[71][2] ;
 wire \mem[71][3] ;
 wire \mem[71][4] ;
 wire \mem[71][5] ;
 wire \mem[71][6] ;
 wire \mem[71][7] ;
 wire \mem[71][8] ;
 wire \mem[71][9] ;
 wire \mem[72][0] ;
 wire \mem[72][10] ;
 wire \mem[72][11] ;
 wire \mem[72][12] ;
 wire \mem[72][13] ;
 wire \mem[72][14] ;
 wire \mem[72][15] ;
 wire \mem[72][1] ;
 wire \mem[72][2] ;
 wire \mem[72][3] ;
 wire \mem[72][4] ;
 wire \mem[72][5] ;
 wire \mem[72][6] ;
 wire \mem[72][7] ;
 wire \mem[72][8] ;
 wire \mem[72][9] ;
 wire \mem[73][0] ;
 wire \mem[73][10] ;
 wire \mem[73][11] ;
 wire \mem[73][12] ;
 wire \mem[73][13] ;
 wire \mem[73][14] ;
 wire \mem[73][15] ;
 wire \mem[73][1] ;
 wire \mem[73][2] ;
 wire \mem[73][3] ;
 wire \mem[73][4] ;
 wire \mem[73][5] ;
 wire \mem[73][6] ;
 wire \mem[73][7] ;
 wire \mem[73][8] ;
 wire \mem[73][9] ;
 wire \mem[74][0] ;
 wire \mem[74][10] ;
 wire \mem[74][11] ;
 wire \mem[74][12] ;
 wire \mem[74][13] ;
 wire \mem[74][14] ;
 wire \mem[74][15] ;
 wire \mem[74][1] ;
 wire \mem[74][2] ;
 wire \mem[74][3] ;
 wire \mem[74][4] ;
 wire \mem[74][5] ;
 wire \mem[74][6] ;
 wire \mem[74][7] ;
 wire \mem[74][8] ;
 wire \mem[74][9] ;
 wire \mem[75][0] ;
 wire \mem[75][10] ;
 wire \mem[75][11] ;
 wire \mem[75][12] ;
 wire \mem[75][13] ;
 wire \mem[75][14] ;
 wire \mem[75][15] ;
 wire \mem[75][1] ;
 wire \mem[75][2] ;
 wire \mem[75][3] ;
 wire \mem[75][4] ;
 wire \mem[75][5] ;
 wire \mem[75][6] ;
 wire \mem[75][7] ;
 wire \mem[75][8] ;
 wire \mem[75][9] ;
 wire \mem[76][0] ;
 wire \mem[76][10] ;
 wire \mem[76][11] ;
 wire \mem[76][12] ;
 wire \mem[76][13] ;
 wire \mem[76][14] ;
 wire \mem[76][15] ;
 wire \mem[76][1] ;
 wire \mem[76][2] ;
 wire \mem[76][3] ;
 wire \mem[76][4] ;
 wire \mem[76][5] ;
 wire \mem[76][6] ;
 wire \mem[76][7] ;
 wire \mem[76][8] ;
 wire \mem[76][9] ;
 wire \mem[77][0] ;
 wire \mem[77][10] ;
 wire \mem[77][11] ;
 wire \mem[77][12] ;
 wire \mem[77][13] ;
 wire \mem[77][14] ;
 wire \mem[77][15] ;
 wire \mem[77][1] ;
 wire \mem[77][2] ;
 wire \mem[77][3] ;
 wire \mem[77][4] ;
 wire \mem[77][5] ;
 wire \mem[77][6] ;
 wire \mem[77][7] ;
 wire \mem[77][8] ;
 wire \mem[77][9] ;
 wire \mem[78][0] ;
 wire \mem[78][10] ;
 wire \mem[78][11] ;
 wire \mem[78][12] ;
 wire \mem[78][13] ;
 wire \mem[78][14] ;
 wire \mem[78][15] ;
 wire \mem[78][1] ;
 wire \mem[78][2] ;
 wire \mem[78][3] ;
 wire \mem[78][4] ;
 wire \mem[78][5] ;
 wire \mem[78][6] ;
 wire \mem[78][7] ;
 wire \mem[78][8] ;
 wire \mem[78][9] ;
 wire \mem[79][0] ;
 wire \mem[79][10] ;
 wire \mem[79][11] ;
 wire \mem[79][12] ;
 wire \mem[79][13] ;
 wire \mem[79][14] ;
 wire \mem[79][15] ;
 wire \mem[79][1] ;
 wire \mem[79][2] ;
 wire \mem[79][3] ;
 wire \mem[79][4] ;
 wire \mem[79][5] ;
 wire \mem[79][6] ;
 wire \mem[79][7] ;
 wire \mem[79][8] ;
 wire \mem[79][9] ;
 wire \mem[7][0] ;
 wire \mem[7][10] ;
 wire \mem[7][11] ;
 wire \mem[7][12] ;
 wire \mem[7][13] ;
 wire \mem[7][14] ;
 wire \mem[7][15] ;
 wire \mem[7][1] ;
 wire \mem[7][2] ;
 wire \mem[7][3] ;
 wire \mem[7][4] ;
 wire \mem[7][5] ;
 wire \mem[7][6] ;
 wire \mem[7][7] ;
 wire \mem[7][8] ;
 wire \mem[7][9] ;
 wire \mem[80][0] ;
 wire \mem[80][10] ;
 wire \mem[80][11] ;
 wire \mem[80][12] ;
 wire \mem[80][13] ;
 wire \mem[80][14] ;
 wire \mem[80][15] ;
 wire \mem[80][1] ;
 wire \mem[80][2] ;
 wire \mem[80][3] ;
 wire \mem[80][4] ;
 wire \mem[80][5] ;
 wire \mem[80][6] ;
 wire \mem[80][7] ;
 wire \mem[80][8] ;
 wire \mem[80][9] ;
 wire \mem[81][0] ;
 wire \mem[81][10] ;
 wire \mem[81][11] ;
 wire \mem[81][12] ;
 wire \mem[81][13] ;
 wire \mem[81][14] ;
 wire \mem[81][15] ;
 wire \mem[81][1] ;
 wire \mem[81][2] ;
 wire \mem[81][3] ;
 wire \mem[81][4] ;
 wire \mem[81][5] ;
 wire \mem[81][6] ;
 wire \mem[81][7] ;
 wire \mem[81][8] ;
 wire \mem[81][9] ;
 wire \mem[82][0] ;
 wire \mem[82][10] ;
 wire \mem[82][11] ;
 wire \mem[82][12] ;
 wire \mem[82][13] ;
 wire \mem[82][14] ;
 wire \mem[82][15] ;
 wire \mem[82][1] ;
 wire \mem[82][2] ;
 wire \mem[82][3] ;
 wire \mem[82][4] ;
 wire \mem[82][5] ;
 wire \mem[82][6] ;
 wire \mem[82][7] ;
 wire \mem[82][8] ;
 wire \mem[82][9] ;
 wire \mem[83][0] ;
 wire \mem[83][10] ;
 wire \mem[83][11] ;
 wire \mem[83][12] ;
 wire \mem[83][13] ;
 wire \mem[83][14] ;
 wire \mem[83][15] ;
 wire \mem[83][1] ;
 wire \mem[83][2] ;
 wire \mem[83][3] ;
 wire \mem[83][4] ;
 wire \mem[83][5] ;
 wire \mem[83][6] ;
 wire \mem[83][7] ;
 wire \mem[83][8] ;
 wire \mem[83][9] ;
 wire \mem[84][0] ;
 wire \mem[84][10] ;
 wire \mem[84][11] ;
 wire \mem[84][12] ;
 wire \mem[84][13] ;
 wire \mem[84][14] ;
 wire \mem[84][15] ;
 wire \mem[84][1] ;
 wire \mem[84][2] ;
 wire \mem[84][3] ;
 wire \mem[84][4] ;
 wire \mem[84][5] ;
 wire \mem[84][6] ;
 wire \mem[84][7] ;
 wire \mem[84][8] ;
 wire \mem[84][9] ;
 wire \mem[85][0] ;
 wire \mem[85][10] ;
 wire \mem[85][11] ;
 wire \mem[85][12] ;
 wire \mem[85][13] ;
 wire \mem[85][14] ;
 wire \mem[85][15] ;
 wire \mem[85][1] ;
 wire \mem[85][2] ;
 wire \mem[85][3] ;
 wire \mem[85][4] ;
 wire \mem[85][5] ;
 wire \mem[85][6] ;
 wire \mem[85][7] ;
 wire \mem[85][8] ;
 wire \mem[85][9] ;
 wire \mem[86][0] ;
 wire \mem[86][10] ;
 wire \mem[86][11] ;
 wire \mem[86][12] ;
 wire \mem[86][13] ;
 wire \mem[86][14] ;
 wire \mem[86][15] ;
 wire \mem[86][1] ;
 wire \mem[86][2] ;
 wire \mem[86][3] ;
 wire \mem[86][4] ;
 wire \mem[86][5] ;
 wire \mem[86][6] ;
 wire \mem[86][7] ;
 wire \mem[86][8] ;
 wire \mem[86][9] ;
 wire \mem[87][0] ;
 wire \mem[87][10] ;
 wire \mem[87][11] ;
 wire \mem[87][12] ;
 wire \mem[87][13] ;
 wire \mem[87][14] ;
 wire \mem[87][15] ;
 wire \mem[87][1] ;
 wire \mem[87][2] ;
 wire \mem[87][3] ;
 wire \mem[87][4] ;
 wire \mem[87][5] ;
 wire \mem[87][6] ;
 wire \mem[87][7] ;
 wire \mem[87][8] ;
 wire \mem[87][9] ;
 wire \mem[88][0] ;
 wire \mem[88][10] ;
 wire \mem[88][11] ;
 wire \mem[88][12] ;
 wire \mem[88][13] ;
 wire \mem[88][14] ;
 wire \mem[88][15] ;
 wire \mem[88][1] ;
 wire \mem[88][2] ;
 wire \mem[88][3] ;
 wire \mem[88][4] ;
 wire \mem[88][5] ;
 wire \mem[88][6] ;
 wire \mem[88][7] ;
 wire \mem[88][8] ;
 wire \mem[88][9] ;
 wire \mem[89][0] ;
 wire \mem[89][10] ;
 wire \mem[89][11] ;
 wire \mem[89][12] ;
 wire \mem[89][13] ;
 wire \mem[89][14] ;
 wire \mem[89][15] ;
 wire \mem[89][1] ;
 wire \mem[89][2] ;
 wire \mem[89][3] ;
 wire \mem[89][4] ;
 wire \mem[89][5] ;
 wire \mem[89][6] ;
 wire \mem[89][7] ;
 wire \mem[89][8] ;
 wire \mem[89][9] ;
 wire \mem[8][0] ;
 wire \mem[8][10] ;
 wire \mem[8][11] ;
 wire \mem[8][12] ;
 wire \mem[8][13] ;
 wire \mem[8][14] ;
 wire \mem[8][15] ;
 wire \mem[8][1] ;
 wire \mem[8][2] ;
 wire \mem[8][3] ;
 wire \mem[8][4] ;
 wire \mem[8][5] ;
 wire \mem[8][6] ;
 wire \mem[8][7] ;
 wire \mem[8][8] ;
 wire \mem[8][9] ;
 wire \mem[90][0] ;
 wire \mem[90][10] ;
 wire \mem[90][11] ;
 wire \mem[90][12] ;
 wire \mem[90][13] ;
 wire \mem[90][14] ;
 wire \mem[90][15] ;
 wire \mem[90][1] ;
 wire \mem[90][2] ;
 wire \mem[90][3] ;
 wire \mem[90][4] ;
 wire \mem[90][5] ;
 wire \mem[90][6] ;
 wire \mem[90][7] ;
 wire \mem[90][8] ;
 wire \mem[90][9] ;
 wire \mem[91][0] ;
 wire \mem[91][10] ;
 wire \mem[91][11] ;
 wire \mem[91][12] ;
 wire \mem[91][13] ;
 wire \mem[91][14] ;
 wire \mem[91][15] ;
 wire \mem[91][1] ;
 wire \mem[91][2] ;
 wire \mem[91][3] ;
 wire \mem[91][4] ;
 wire \mem[91][5] ;
 wire \mem[91][6] ;
 wire \mem[91][7] ;
 wire \mem[91][8] ;
 wire \mem[91][9] ;
 wire \mem[92][0] ;
 wire \mem[92][10] ;
 wire \mem[92][11] ;
 wire \mem[92][12] ;
 wire \mem[92][13] ;
 wire \mem[92][14] ;
 wire \mem[92][15] ;
 wire \mem[92][1] ;
 wire \mem[92][2] ;
 wire \mem[92][3] ;
 wire \mem[92][4] ;
 wire \mem[92][5] ;
 wire \mem[92][6] ;
 wire \mem[92][7] ;
 wire \mem[92][8] ;
 wire \mem[92][9] ;
 wire \mem[93][0] ;
 wire \mem[93][10] ;
 wire \mem[93][11] ;
 wire \mem[93][12] ;
 wire \mem[93][13] ;
 wire \mem[93][14] ;
 wire \mem[93][15] ;
 wire \mem[93][1] ;
 wire \mem[93][2] ;
 wire \mem[93][3] ;
 wire \mem[93][4] ;
 wire \mem[93][5] ;
 wire \mem[93][6] ;
 wire \mem[93][7] ;
 wire \mem[93][8] ;
 wire \mem[93][9] ;
 wire \mem[94][0] ;
 wire \mem[94][10] ;
 wire \mem[94][11] ;
 wire \mem[94][12] ;
 wire \mem[94][13] ;
 wire \mem[94][14] ;
 wire \mem[94][15] ;
 wire \mem[94][1] ;
 wire \mem[94][2] ;
 wire \mem[94][3] ;
 wire \mem[94][4] ;
 wire \mem[94][5] ;
 wire \mem[94][6] ;
 wire \mem[94][7] ;
 wire \mem[94][8] ;
 wire \mem[94][9] ;
 wire \mem[95][0] ;
 wire \mem[95][10] ;
 wire \mem[95][11] ;
 wire \mem[95][12] ;
 wire \mem[95][13] ;
 wire \mem[95][14] ;
 wire \mem[95][15] ;
 wire \mem[95][1] ;
 wire \mem[95][2] ;
 wire \mem[95][3] ;
 wire \mem[95][4] ;
 wire \mem[95][5] ;
 wire \mem[95][6] ;
 wire \mem[95][7] ;
 wire \mem[95][8] ;
 wire \mem[95][9] ;
 wire \mem[96][0] ;
 wire \mem[96][10] ;
 wire \mem[96][11] ;
 wire \mem[96][12] ;
 wire \mem[96][13] ;
 wire \mem[96][14] ;
 wire \mem[96][15] ;
 wire \mem[96][1] ;
 wire \mem[96][2] ;
 wire \mem[96][3] ;
 wire \mem[96][4] ;
 wire \mem[96][5] ;
 wire \mem[96][6] ;
 wire \mem[96][7] ;
 wire \mem[96][8] ;
 wire \mem[96][9] ;
 wire \mem[97][0] ;
 wire \mem[97][10] ;
 wire \mem[97][11] ;
 wire \mem[97][12] ;
 wire \mem[97][13] ;
 wire \mem[97][14] ;
 wire \mem[97][15] ;
 wire \mem[97][1] ;
 wire \mem[97][2] ;
 wire \mem[97][3] ;
 wire \mem[97][4] ;
 wire \mem[97][5] ;
 wire \mem[97][6] ;
 wire \mem[97][7] ;
 wire \mem[97][8] ;
 wire \mem[97][9] ;
 wire \mem[98][0] ;
 wire \mem[98][10] ;
 wire \mem[98][11] ;
 wire \mem[98][12] ;
 wire \mem[98][13] ;
 wire \mem[98][14] ;
 wire \mem[98][15] ;
 wire \mem[98][1] ;
 wire \mem[98][2] ;
 wire \mem[98][3] ;
 wire \mem[98][4] ;
 wire \mem[98][5] ;
 wire \mem[98][6] ;
 wire \mem[98][7] ;
 wire \mem[98][8] ;
 wire \mem[98][9] ;
 wire \mem[99][0] ;
 wire \mem[99][10] ;
 wire \mem[99][11] ;
 wire \mem[99][12] ;
 wire \mem[99][13] ;
 wire \mem[99][14] ;
 wire \mem[99][15] ;
 wire \mem[99][1] ;
 wire \mem[99][2] ;
 wire \mem[99][3] ;
 wire \mem[99][4] ;
 wire \mem[99][5] ;
 wire \mem[99][6] ;
 wire \mem[99][7] ;
 wire \mem[99][8] ;
 wire \mem[99][9] ;
 wire \mem[9][0] ;
 wire \mem[9][10] ;
 wire \mem[9][11] ;
 wire \mem[9][12] ;
 wire \mem[9][13] ;
 wire \mem[9][14] ;
 wire \mem[9][15] ;
 wire \mem[9][1] ;
 wire \mem[9][2] ;
 wire \mem[9][3] ;
 wire \mem[9][4] ;
 wire \mem[9][5] ;
 wire \mem[9][6] ;
 wire \mem[9][7] ;
 wire \mem[9][8] ;
 wire \mem[9][9] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire clknet_leaf_0_i_clk;
 wire clknet_leaf_1_i_clk;
 wire clknet_leaf_2_i_clk;
 wire clknet_leaf_3_i_clk;
 wire clknet_leaf_4_i_clk;
 wire clknet_leaf_5_i_clk;
 wire clknet_leaf_6_i_clk;
 wire clknet_leaf_7_i_clk;
 wire clknet_leaf_8_i_clk;
 wire clknet_leaf_9_i_clk;
 wire clknet_leaf_10_i_clk;
 wire clknet_leaf_11_i_clk;
 wire clknet_leaf_12_i_clk;
 wire clknet_leaf_13_i_clk;
 wire clknet_leaf_14_i_clk;
 wire clknet_leaf_15_i_clk;
 wire clknet_leaf_16_i_clk;
 wire clknet_leaf_17_i_clk;
 wire clknet_leaf_18_i_clk;
 wire clknet_leaf_19_i_clk;
 wire clknet_leaf_20_i_clk;
 wire clknet_leaf_21_i_clk;
 wire clknet_leaf_22_i_clk;
 wire clknet_leaf_23_i_clk;
 wire clknet_leaf_24_i_clk;
 wire clknet_leaf_25_i_clk;
 wire clknet_leaf_26_i_clk;
 wire clknet_leaf_27_i_clk;
 wire clknet_leaf_28_i_clk;
 wire clknet_leaf_29_i_clk;
 wire clknet_leaf_30_i_clk;
 wire clknet_leaf_31_i_clk;
 wire clknet_leaf_32_i_clk;
 wire clknet_leaf_33_i_clk;
 wire clknet_leaf_34_i_clk;
 wire clknet_leaf_35_i_clk;
 wire clknet_leaf_36_i_clk;
 wire clknet_leaf_37_i_clk;
 wire clknet_leaf_38_i_clk;
 wire clknet_leaf_39_i_clk;
 wire clknet_leaf_40_i_clk;
 wire clknet_leaf_41_i_clk;
 wire clknet_leaf_42_i_clk;
 wire clknet_leaf_43_i_clk;
 wire clknet_leaf_44_i_clk;
 wire clknet_leaf_45_i_clk;
 wire clknet_leaf_46_i_clk;
 wire clknet_leaf_47_i_clk;
 wire clknet_leaf_48_i_clk;
 wire clknet_leaf_49_i_clk;
 wire clknet_leaf_50_i_clk;
 wire clknet_leaf_51_i_clk;
 wire clknet_leaf_52_i_clk;
 wire clknet_leaf_53_i_clk;
 wire clknet_leaf_54_i_clk;
 wire clknet_leaf_55_i_clk;
 wire clknet_leaf_56_i_clk;
 wire clknet_leaf_57_i_clk;
 wire clknet_leaf_58_i_clk;
 wire clknet_leaf_59_i_clk;
 wire clknet_leaf_60_i_clk;
 wire clknet_leaf_61_i_clk;
 wire clknet_leaf_62_i_clk;
 wire clknet_leaf_63_i_clk;
 wire clknet_leaf_64_i_clk;
 wire clknet_leaf_65_i_clk;
 wire clknet_leaf_66_i_clk;
 wire clknet_leaf_67_i_clk;
 wire clknet_leaf_68_i_clk;
 wire clknet_leaf_69_i_clk;
 wire clknet_leaf_70_i_clk;
 wire clknet_leaf_71_i_clk;
 wire clknet_leaf_72_i_clk;
 wire clknet_leaf_73_i_clk;
 wire clknet_leaf_74_i_clk;
 wire clknet_leaf_75_i_clk;
 wire clknet_leaf_76_i_clk;
 wire clknet_leaf_77_i_clk;
 wire clknet_leaf_78_i_clk;
 wire clknet_leaf_79_i_clk;
 wire clknet_leaf_80_i_clk;
 wire clknet_leaf_81_i_clk;
 wire clknet_leaf_82_i_clk;
 wire clknet_leaf_83_i_clk;
 wire clknet_leaf_84_i_clk;
 wire clknet_leaf_85_i_clk;
 wire clknet_leaf_86_i_clk;
 wire clknet_leaf_87_i_clk;
 wire clknet_leaf_88_i_clk;
 wire clknet_leaf_89_i_clk;
 wire clknet_leaf_90_i_clk;
 wire clknet_leaf_91_i_clk;
 wire clknet_leaf_92_i_clk;
 wire clknet_leaf_93_i_clk;
 wire clknet_leaf_94_i_clk;
 wire clknet_leaf_95_i_clk;
 wire clknet_leaf_96_i_clk;
 wire clknet_leaf_97_i_clk;
 wire clknet_leaf_98_i_clk;
 wire clknet_leaf_99_i_clk;
 wire clknet_leaf_100_i_clk;
 wire clknet_leaf_101_i_clk;
 wire clknet_leaf_102_i_clk;
 wire clknet_leaf_103_i_clk;
 wire clknet_leaf_104_i_clk;
 wire clknet_leaf_105_i_clk;
 wire clknet_leaf_106_i_clk;
 wire clknet_leaf_107_i_clk;
 wire clknet_leaf_108_i_clk;
 wire clknet_leaf_109_i_clk;
 wire clknet_leaf_110_i_clk;
 wire clknet_leaf_111_i_clk;
 wire clknet_leaf_112_i_clk;
 wire clknet_leaf_113_i_clk;
 wire clknet_leaf_114_i_clk;
 wire clknet_leaf_115_i_clk;
 wire clknet_leaf_116_i_clk;
 wire clknet_leaf_117_i_clk;
 wire clknet_leaf_118_i_clk;
 wire clknet_leaf_119_i_clk;
 wire clknet_leaf_120_i_clk;
 wire clknet_leaf_121_i_clk;
 wire clknet_leaf_122_i_clk;
 wire clknet_leaf_123_i_clk;
 wire clknet_leaf_124_i_clk;
 wire clknet_leaf_125_i_clk;
 wire clknet_leaf_126_i_clk;
 wire clknet_leaf_127_i_clk;
 wire clknet_leaf_128_i_clk;
 wire clknet_leaf_129_i_clk;
 wire clknet_leaf_130_i_clk;
 wire clknet_leaf_131_i_clk;
 wire clknet_leaf_132_i_clk;
 wire clknet_leaf_133_i_clk;
 wire clknet_leaf_134_i_clk;
 wire clknet_leaf_135_i_clk;
 wire clknet_leaf_136_i_clk;
 wire clknet_leaf_137_i_clk;
 wire clknet_leaf_138_i_clk;
 wire clknet_leaf_139_i_clk;
 wire clknet_leaf_140_i_clk;
 wire clknet_leaf_141_i_clk;
 wire clknet_leaf_142_i_clk;
 wire clknet_leaf_143_i_clk;
 wire clknet_leaf_144_i_clk;
 wire clknet_leaf_145_i_clk;
 wire clknet_leaf_146_i_clk;
 wire clknet_leaf_147_i_clk;
 wire clknet_leaf_148_i_clk;
 wire clknet_leaf_149_i_clk;
 wire clknet_leaf_150_i_clk;
 wire clknet_leaf_151_i_clk;
 wire clknet_leaf_152_i_clk;
 wire clknet_leaf_153_i_clk;
 wire clknet_leaf_154_i_clk;
 wire clknet_leaf_155_i_clk;
 wire clknet_leaf_156_i_clk;
 wire clknet_leaf_157_i_clk;
 wire clknet_leaf_158_i_clk;
 wire clknet_leaf_159_i_clk;
 wire clknet_leaf_160_i_clk;
 wire clknet_leaf_161_i_clk;
 wire clknet_leaf_162_i_clk;
 wire clknet_leaf_163_i_clk;
 wire clknet_leaf_164_i_clk;
 wire clknet_leaf_165_i_clk;
 wire clknet_leaf_166_i_clk;
 wire clknet_leaf_167_i_clk;
 wire clknet_leaf_168_i_clk;
 wire clknet_leaf_169_i_clk;
 wire clknet_leaf_170_i_clk;
 wire clknet_leaf_171_i_clk;
 wire clknet_leaf_172_i_clk;
 wire clknet_leaf_173_i_clk;
 wire clknet_leaf_174_i_clk;
 wire clknet_leaf_175_i_clk;
 wire clknet_leaf_176_i_clk;
 wire clknet_leaf_177_i_clk;
 wire clknet_leaf_178_i_clk;
 wire clknet_leaf_179_i_clk;
 wire clknet_leaf_180_i_clk;
 wire clknet_leaf_181_i_clk;
 wire clknet_leaf_182_i_clk;
 wire clknet_leaf_183_i_clk;
 wire clknet_leaf_184_i_clk;
 wire clknet_leaf_185_i_clk;
 wire clknet_leaf_186_i_clk;
 wire clknet_leaf_187_i_clk;
 wire clknet_leaf_188_i_clk;
 wire clknet_leaf_189_i_clk;
 wire clknet_leaf_190_i_clk;
 wire clknet_leaf_191_i_clk;
 wire clknet_leaf_192_i_clk;
 wire clknet_leaf_193_i_clk;
 wire clknet_leaf_194_i_clk;
 wire clknet_leaf_195_i_clk;
 wire clknet_leaf_196_i_clk;
 wire clknet_leaf_197_i_clk;
 wire clknet_leaf_198_i_clk;
 wire clknet_leaf_199_i_clk;
 wire clknet_leaf_200_i_clk;
 wire clknet_leaf_201_i_clk;
 wire clknet_leaf_202_i_clk;
 wire clknet_leaf_203_i_clk;
 wire clknet_leaf_204_i_clk;
 wire clknet_leaf_205_i_clk;
 wire clknet_leaf_206_i_clk;
 wire clknet_leaf_207_i_clk;
 wire clknet_leaf_208_i_clk;
 wire clknet_leaf_209_i_clk;
 wire clknet_leaf_210_i_clk;
 wire clknet_leaf_211_i_clk;
 wire clknet_leaf_212_i_clk;
 wire clknet_leaf_213_i_clk;
 wire clknet_leaf_214_i_clk;
 wire clknet_leaf_215_i_clk;
 wire clknet_leaf_216_i_clk;
 wire clknet_leaf_217_i_clk;
 wire clknet_leaf_218_i_clk;
 wire clknet_leaf_219_i_clk;
 wire clknet_leaf_220_i_clk;
 wire clknet_leaf_221_i_clk;
 wire clknet_leaf_222_i_clk;
 wire clknet_leaf_223_i_clk;
 wire clknet_leaf_224_i_clk;
 wire clknet_leaf_225_i_clk;
 wire clknet_leaf_226_i_clk;
 wire clknet_leaf_227_i_clk;
 wire clknet_leaf_228_i_clk;
 wire clknet_leaf_229_i_clk;
 wire clknet_leaf_230_i_clk;
 wire clknet_leaf_231_i_clk;
 wire clknet_leaf_232_i_clk;
 wire clknet_leaf_233_i_clk;
 wire clknet_leaf_234_i_clk;
 wire clknet_leaf_235_i_clk;
 wire clknet_leaf_236_i_clk;
 wire clknet_leaf_237_i_clk;
 wire clknet_leaf_238_i_clk;
 wire clknet_leaf_239_i_clk;
 wire clknet_leaf_240_i_clk;
 wire clknet_leaf_241_i_clk;
 wire clknet_leaf_242_i_clk;
 wire clknet_leaf_243_i_clk;
 wire clknet_leaf_244_i_clk;
 wire clknet_leaf_245_i_clk;
 wire clknet_leaf_246_i_clk;
 wire clknet_leaf_247_i_clk;
 wire clknet_leaf_248_i_clk;
 wire clknet_leaf_249_i_clk;
 wire clknet_leaf_250_i_clk;
 wire clknet_leaf_251_i_clk;
 wire clknet_leaf_252_i_clk;
 wire clknet_leaf_253_i_clk;
 wire clknet_leaf_254_i_clk;
 wire clknet_leaf_255_i_clk;
 wire clknet_leaf_256_i_clk;
 wire clknet_leaf_257_i_clk;
 wire clknet_leaf_258_i_clk;
 wire clknet_leaf_259_i_clk;
 wire clknet_leaf_260_i_clk;
 wire clknet_leaf_261_i_clk;
 wire clknet_leaf_262_i_clk;
 wire clknet_leaf_263_i_clk;
 wire clknet_leaf_264_i_clk;
 wire clknet_leaf_265_i_clk;
 wire clknet_leaf_266_i_clk;
 wire clknet_leaf_267_i_clk;
 wire clknet_leaf_268_i_clk;
 wire clknet_leaf_269_i_clk;
 wire clknet_leaf_270_i_clk;
 wire clknet_leaf_271_i_clk;
 wire clknet_leaf_272_i_clk;
 wire clknet_leaf_273_i_clk;
 wire clknet_leaf_274_i_clk;
 wire clknet_leaf_275_i_clk;
 wire clknet_leaf_276_i_clk;
 wire clknet_leaf_277_i_clk;
 wire clknet_leaf_278_i_clk;
 wire clknet_leaf_279_i_clk;
 wire clknet_leaf_280_i_clk;
 wire clknet_leaf_281_i_clk;
 wire clknet_leaf_282_i_clk;
 wire clknet_leaf_283_i_clk;
 wire clknet_leaf_284_i_clk;
 wire clknet_leaf_285_i_clk;
 wire clknet_leaf_286_i_clk;
 wire clknet_leaf_287_i_clk;
 wire clknet_leaf_288_i_clk;
 wire clknet_0_i_clk;
 wire clknet_1_0_0_i_clk;
 wire clknet_1_0_1_i_clk;
 wire clknet_1_1_0_i_clk;
 wire clknet_1_1_1_i_clk;
 wire clknet_2_0_0_i_clk;
 wire clknet_2_0_1_i_clk;
 wire clknet_2_1_0_i_clk;
 wire clknet_2_1_1_i_clk;
 wire clknet_2_2_0_i_clk;
 wire clknet_2_2_1_i_clk;
 wire clknet_2_3_0_i_clk;
 wire clknet_2_3_1_i_clk;
 wire clknet_3_0_0_i_clk;
 wire clknet_3_1_0_i_clk;
 wire clknet_3_2_0_i_clk;
 wire clknet_3_3_0_i_clk;
 wire clknet_3_4_0_i_clk;
 wire clknet_3_5_0_i_clk;
 wire clknet_3_6_0_i_clk;
 wire clknet_3_7_0_i_clk;
 wire clknet_4_0_0_i_clk;
 wire clknet_4_1_0_i_clk;
 wire clknet_4_2_0_i_clk;
 wire clknet_4_3_0_i_clk;
 wire clknet_4_4_0_i_clk;
 wire clknet_4_5_0_i_clk;
 wire clknet_4_6_0_i_clk;
 wire clknet_4_7_0_i_clk;
 wire clknet_4_8_0_i_clk;
 wire clknet_4_9_0_i_clk;
 wire clknet_4_10_0_i_clk;
 wire clknet_4_11_0_i_clk;
 wire clknet_4_12_0_i_clk;
 wire clknet_4_13_0_i_clk;
 wire clknet_4_14_0_i_clk;
 wire clknet_4_15_0_i_clk;
 wire clknet_5_0_0_i_clk;
 wire clknet_5_1_0_i_clk;
 wire clknet_5_2_0_i_clk;
 wire clknet_5_3_0_i_clk;
 wire clknet_5_4_0_i_clk;
 wire clknet_5_5_0_i_clk;
 wire clknet_5_6_0_i_clk;
 wire clknet_5_7_0_i_clk;
 wire clknet_5_8_0_i_clk;
 wire clknet_5_9_0_i_clk;
 wire clknet_5_10_0_i_clk;
 wire clknet_5_11_0_i_clk;
 wire clknet_5_12_0_i_clk;
 wire clknet_5_13_0_i_clk;
 wire clknet_5_14_0_i_clk;
 wire clknet_5_15_0_i_clk;
 wire clknet_5_16_0_i_clk;
 wire clknet_5_17_0_i_clk;
 wire clknet_5_18_0_i_clk;
 wire clknet_5_19_0_i_clk;
 wire clknet_5_20_0_i_clk;
 wire clknet_5_21_0_i_clk;
 wire clknet_5_22_0_i_clk;
 wire clknet_5_23_0_i_clk;
 wire clknet_5_24_0_i_clk;
 wire clknet_5_25_0_i_clk;
 wire clknet_5_26_0_i_clk;
 wire clknet_5_27_0_i_clk;
 wire clknet_5_28_0_i_clk;
 wire clknet_5_29_0_i_clk;
 wire clknet_5_30_0_i_clk;
 wire clknet_5_31_0_i_clk;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net1657;
 wire net1658;
 wire net1659;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1687;
 wire net1688;
 wire net1689;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;

 sky130_fd_sc_hd__inv_2 _06406_ (.A(net6),
    .Y(_02355_));
 sky130_fd_sc_hd__clkbuf_4 _06407_ (.A(_02355_),
    .X(_02356_));
 sky130_fd_sc_hd__inv_6 _06408_ (.A(net5),
    .Y(_02357_));
 sky130_fd_sc_hd__clkbuf_8 _06409_ (.A(_02357_),
    .X(_02358_));
 sky130_fd_sc_hd__buf_4 _06410_ (.A(net2),
    .X(_02359_));
 sky130_fd_sc_hd__buf_6 _06411_ (.A(net1),
    .X(_02360_));
 sky130_fd_sc_hd__nand2b_1 _06412_ (.A_N(_02359_),
    .B(_02360_),
    .Y(_02361_));
 sky130_fd_sc_hd__clkbuf_4 _06413_ (.A(_02361_),
    .X(_02362_));
 sky130_fd_sc_hd__buf_4 _06414_ (.A(_02362_),
    .X(_02363_));
 sky130_fd_sc_hd__and2_1 _06415_ (.A(net3),
    .B(net4),
    .X(_02364_));
 sky130_fd_sc_hd__buf_2 _06416_ (.A(_02364_),
    .X(_02365_));
 sky130_fd_sc_hd__buf_4 _06417_ (.A(_02365_),
    .X(_02366_));
 sky130_fd_sc_hd__o21a_1 _06418_ (.A1(\mem[29][0] ),
    .A2(_02363_),
    .B1(_02366_),
    .X(_02367_));
 sky130_fd_sc_hd__nand2b_1 _06419_ (.A_N(net1),
    .B(_02359_),
    .Y(_02368_));
 sky130_fd_sc_hd__buf_8 _06420_ (.A(_02368_),
    .X(_02369_));
 sky130_fd_sc_hd__buf_6 _06421_ (.A(_02369_),
    .X(_02370_));
 sky130_fd_sc_hd__nand2_2 _06422_ (.A(_02360_),
    .B(_02359_),
    .Y(_02371_));
 sky130_fd_sc_hd__buf_4 _06423_ (.A(_02371_),
    .X(_02372_));
 sky130_fd_sc_hd__buf_6 _06424_ (.A(_02360_),
    .X(_02373_));
 sky130_fd_sc_hd__buf_8 _06425_ (.A(_02373_),
    .X(_02374_));
 sky130_fd_sc_hd__clkbuf_16 _06426_ (.A(_02359_),
    .X(_02375_));
 sky130_fd_sc_hd__or3_1 _06427_ (.A(_02374_),
    .B(_02375_),
    .C(\mem[28][0] ),
    .X(_02376_));
 sky130_fd_sc_hd__o221a_1 _06428_ (.A1(\mem[30][0] ),
    .A2(_02370_),
    .B1(_02372_),
    .B2(\mem[31][0] ),
    .C1(_02376_),
    .X(_02377_));
 sky130_fd_sc_hd__or2_2 _06429_ (.A(_02360_),
    .B(_02359_),
    .X(_02378_));
 sky130_fd_sc_hd__buf_4 _06430_ (.A(_02378_),
    .X(_02379_));
 sky130_fd_sc_hd__buf_4 _06431_ (.A(_02379_),
    .X(_02380_));
 sky130_fd_sc_hd__buf_8 _06432_ (.A(net3),
    .X(_02381_));
 sky130_fd_sc_hd__nor2_1 _06433_ (.A(_02381_),
    .B(net4),
    .Y(_02382_));
 sky130_fd_sc_hd__clkbuf_8 _06434_ (.A(_02382_),
    .X(_02383_));
 sky130_fd_sc_hd__o21a_1 _06435_ (.A1(\mem[16][0] ),
    .A2(_02380_),
    .B1(_02383_),
    .X(_02384_));
 sky130_fd_sc_hd__buf_6 _06436_ (.A(_02362_),
    .X(_02385_));
 sky130_fd_sc_hd__buf_6 _06437_ (.A(_02371_),
    .X(_02386_));
 sky130_fd_sc_hd__buf_4 _06438_ (.A(_02373_),
    .X(_02387_));
 sky130_fd_sc_hd__buf_6 _06439_ (.A(net2),
    .X(_02388_));
 sky130_fd_sc_hd__buf_4 _06440_ (.A(_02388_),
    .X(_02389_));
 sky130_fd_sc_hd__or3b_1 _06441_ (.A(_02387_),
    .B(\mem[18][0] ),
    .C_N(_02389_),
    .X(_02390_));
 sky130_fd_sc_hd__o221a_1 _06442_ (.A1(\mem[17][0] ),
    .A2(_02385_),
    .B1(_02386_),
    .B2(\mem[19][0] ),
    .C1(_02390_),
    .X(_02391_));
 sky130_fd_sc_hd__a22o_1 _06443_ (.A1(_02367_),
    .A2(_02377_),
    .B1(_02384_),
    .B2(_02391_),
    .X(_02392_));
 sky130_fd_sc_hd__buf_6 _06444_ (.A(_02369_),
    .X(_02393_));
 sky130_fd_sc_hd__buf_4 _06445_ (.A(_02393_),
    .X(_02394_));
 sky130_fd_sc_hd__buf_4 _06446_ (.A(_02379_),
    .X(_02395_));
 sky130_fd_sc_hd__nor2b_4 _06447_ (.A(_02381_),
    .B_N(net4),
    .Y(_02396_));
 sky130_fd_sc_hd__buf_4 _06448_ (.A(_02396_),
    .X(_02397_));
 sky130_fd_sc_hd__o21a_1 _06449_ (.A1(\mem[24][0] ),
    .A2(_02395_),
    .B1(_02397_),
    .X(_02398_));
 sky130_fd_sc_hd__buf_4 _06450_ (.A(_02362_),
    .X(_02399_));
 sky130_fd_sc_hd__buf_4 _06451_ (.A(_02371_),
    .X(_02400_));
 sky130_fd_sc_hd__buf_6 _06452_ (.A(_02400_),
    .X(_02401_));
 sky130_fd_sc_hd__o22a_1 _06453_ (.A1(\mem[25][0] ),
    .A2(_02399_),
    .B1(_02401_),
    .B2(\mem[27][0] ),
    .X(_02402_));
 sky130_fd_sc_hd__o211a_1 _06454_ (.A1(\mem[26][0] ),
    .A2(_02394_),
    .B1(_02398_),
    .C1(_02402_),
    .X(_02403_));
 sky130_fd_sc_hd__buf_8 _06455_ (.A(_02361_),
    .X(_02404_));
 sky130_fd_sc_hd__buf_6 _06456_ (.A(_02404_),
    .X(_02405_));
 sky130_fd_sc_hd__buf_6 _06457_ (.A(_02405_),
    .X(_02406_));
 sky130_fd_sc_hd__buf_8 _06458_ (.A(_02369_),
    .X(_02407_));
 sky130_fd_sc_hd__buf_4 _06459_ (.A(_02371_),
    .X(_02408_));
 sky130_fd_sc_hd__buf_6 _06460_ (.A(_02408_),
    .X(_02409_));
 sky130_fd_sc_hd__buf_8 _06461_ (.A(_02360_),
    .X(_02410_));
 sky130_fd_sc_hd__buf_8 _06462_ (.A(_02410_),
    .X(_02411_));
 sky130_fd_sc_hd__buf_4 _06463_ (.A(_02388_),
    .X(_02412_));
 sky130_fd_sc_hd__or3_1 _06464_ (.A(_02411_),
    .B(_02412_),
    .C(\mem[20][0] ),
    .X(_02413_));
 sky130_fd_sc_hd__o221a_1 _06465_ (.A1(\mem[22][0] ),
    .A2(_02407_),
    .B1(_02409_),
    .B2(\mem[23][0] ),
    .C1(_02413_),
    .X(_02414_));
 sky130_fd_sc_hd__and2b_1 _06466_ (.A_N(net4),
    .B(_02381_),
    .X(_02415_));
 sky130_fd_sc_hd__buf_6 _06467_ (.A(_02415_),
    .X(_02416_));
 sky130_fd_sc_hd__buf_4 _06468_ (.A(_02416_),
    .X(_02417_));
 sky130_fd_sc_hd__o211a_1 _06469_ (.A1(\mem[21][0] ),
    .A2(_02406_),
    .B1(_02414_),
    .C1(_02417_),
    .X(_02418_));
 sky130_fd_sc_hd__or4_2 _06470_ (.A(_02358_),
    .B(_02392_),
    .C(_02403_),
    .D(_02418_),
    .X(_02419_));
 sky130_fd_sc_hd__clkbuf_4 _06471_ (.A(net5),
    .X(_02420_));
 sky130_fd_sc_hd__clkbuf_4 _06472_ (.A(_02420_),
    .X(_02421_));
 sky130_fd_sc_hd__buf_4 _06473_ (.A(_02365_),
    .X(_02422_));
 sky130_fd_sc_hd__or2_1 _06474_ (.A(\mem[13][0] ),
    .B(_02385_),
    .X(_02423_));
 sky130_fd_sc_hd__buf_4 _06475_ (.A(_02371_),
    .X(_02424_));
 sky130_fd_sc_hd__or3_1 _06476_ (.A(_02374_),
    .B(_02375_),
    .C(\mem[12][0] ),
    .X(_02425_));
 sky130_fd_sc_hd__o221a_1 _06477_ (.A1(\mem[14][0] ),
    .A2(_02370_),
    .B1(_02424_),
    .B2(\mem[15][0] ),
    .C1(_02425_),
    .X(_02426_));
 sky130_fd_sc_hd__buf_12 _06478_ (.A(_02410_),
    .X(_02427_));
 sky130_fd_sc_hd__buf_6 _06479_ (.A(_02427_),
    .X(_02428_));
 sky130_fd_sc_hd__buf_6 _06480_ (.A(_02359_),
    .X(_02429_));
 sky130_fd_sc_hd__buf_6 _06481_ (.A(_02429_),
    .X(_02430_));
 sky130_fd_sc_hd__o31a_1 _06482_ (.A1(\mem[0][0] ),
    .A2(_02428_),
    .A3(_02430_),
    .B1(_02383_),
    .X(_02431_));
 sky130_fd_sc_hd__buf_4 _06483_ (.A(_02360_),
    .X(_02432_));
 sky130_fd_sc_hd__buf_4 _06484_ (.A(_02388_),
    .X(_02433_));
 sky130_fd_sc_hd__or3b_1 _06485_ (.A(_02432_),
    .B(\mem[2][0] ),
    .C_N(_02433_),
    .X(_02434_));
 sky130_fd_sc_hd__o221a_1 _06486_ (.A1(\mem[1][0] ),
    .A2(_02385_),
    .B1(_02386_),
    .B2(\mem[3][0] ),
    .C1(_02434_),
    .X(_02435_));
 sky130_fd_sc_hd__a32o_1 _06487_ (.A1(_02422_),
    .A2(_02423_),
    .A3(_02426_),
    .B1(_02431_),
    .B2(_02435_),
    .X(_02436_));
 sky130_fd_sc_hd__buf_6 _06488_ (.A(_02393_),
    .X(_02437_));
 sky130_fd_sc_hd__buf_4 _06489_ (.A(_02379_),
    .X(_02438_));
 sky130_fd_sc_hd__clkbuf_8 _06490_ (.A(_02396_),
    .X(_02439_));
 sky130_fd_sc_hd__o21a_1 _06491_ (.A1(\mem[8][0] ),
    .A2(_02438_),
    .B1(_02439_),
    .X(_02440_));
 sky130_fd_sc_hd__clkbuf_8 _06492_ (.A(_02404_),
    .X(_02441_));
 sky130_fd_sc_hd__buf_6 _06493_ (.A(_02400_),
    .X(_02442_));
 sky130_fd_sc_hd__o22a_1 _06494_ (.A1(\mem[9][0] ),
    .A2(_02441_),
    .B1(_02442_),
    .B2(\mem[11][0] ),
    .X(_02443_));
 sky130_fd_sc_hd__o211a_1 _06495_ (.A1(\mem[10][0] ),
    .A2(_02437_),
    .B1(_02440_),
    .C1(_02443_),
    .X(_02444_));
 sky130_fd_sc_hd__buf_4 _06496_ (.A(_02369_),
    .X(_02445_));
 sky130_fd_sc_hd__clkbuf_4 _06497_ (.A(_02408_),
    .X(_02446_));
 sky130_fd_sc_hd__clkbuf_4 _06498_ (.A(_02410_),
    .X(_02447_));
 sky130_fd_sc_hd__or3_1 _06499_ (.A(_02447_),
    .B(_02429_),
    .C(\mem[4][0] ),
    .X(_02448_));
 sky130_fd_sc_hd__o221a_2 _06500_ (.A1(\mem[6][0] ),
    .A2(_02445_),
    .B1(_02446_),
    .B2(\mem[7][0] ),
    .C1(_02448_),
    .X(_02449_));
 sky130_fd_sc_hd__clkbuf_16 _06501_ (.A(_02416_),
    .X(_02450_));
 sky130_fd_sc_hd__o211a_1 _06502_ (.A1(\mem[5][0] ),
    .A2(_02406_),
    .B1(_02449_),
    .C1(_02450_),
    .X(_02451_));
 sky130_fd_sc_hd__or4_1 _06503_ (.A(_02421_),
    .B(_02436_),
    .C(_02444_),
    .D(_02451_),
    .X(_02452_));
 sky130_fd_sc_hd__buf_6 _06504_ (.A(_02420_),
    .X(_02453_));
 sky130_fd_sc_hd__buf_6 _06505_ (.A(_02382_),
    .X(_02454_));
 sky130_fd_sc_hd__buf_6 _06506_ (.A(_02454_),
    .X(_02455_));
 sky130_fd_sc_hd__buf_4 _06507_ (.A(_02455_),
    .X(_02456_));
 sky130_fd_sc_hd__buf_6 _06508_ (.A(_02360_),
    .X(_02457_));
 sky130_fd_sc_hd__buf_6 _06509_ (.A(_02457_),
    .X(_02458_));
 sky130_fd_sc_hd__buf_6 _06510_ (.A(_02359_),
    .X(_02459_));
 sky130_fd_sc_hd__buf_6 _06511_ (.A(_02459_),
    .X(_02460_));
 sky130_fd_sc_hd__buf_6 _06512_ (.A(_02460_),
    .X(_02461_));
 sky130_fd_sc_hd__mux4_1 _06513_ (.A0(\mem[32][0] ),
    .A1(\mem[33][0] ),
    .A2(\mem[34][0] ),
    .A3(\mem[35][0] ),
    .S0(_02458_),
    .S1(_02461_),
    .X(_02462_));
 sky130_fd_sc_hd__buf_4 _06514_ (.A(_02415_),
    .X(_02463_));
 sky130_fd_sc_hd__buf_6 _06515_ (.A(_02463_),
    .X(_02464_));
 sky130_fd_sc_hd__buf_8 _06516_ (.A(_02464_),
    .X(_02465_));
 sky130_fd_sc_hd__clkbuf_4 _06517_ (.A(_02373_),
    .X(_02466_));
 sky130_fd_sc_hd__buf_8 _06518_ (.A(_02466_),
    .X(_02467_));
 sky130_fd_sc_hd__buf_6 _06519_ (.A(_02460_),
    .X(_02468_));
 sky130_fd_sc_hd__mux4_1 _06520_ (.A0(\mem[36][0] ),
    .A1(\mem[37][0] ),
    .A2(\mem[38][0] ),
    .A3(\mem[39][0] ),
    .S0(_02467_),
    .S1(_02468_),
    .X(_02469_));
 sky130_fd_sc_hd__a22o_1 _06521_ (.A1(_02456_),
    .A2(_02462_),
    .B1(_02465_),
    .B2(_02469_),
    .X(_02470_));
 sky130_fd_sc_hd__inv_2 _06522_ (.A(_02381_),
    .Y(_02471_));
 sky130_fd_sc_hd__buf_4 _06523_ (.A(_02471_),
    .X(_02472_));
 sky130_fd_sc_hd__mux4_1 _06524_ (.A0(\mem[44][0] ),
    .A1(\mem[45][0] ),
    .A2(\mem[46][0] ),
    .A3(\mem[47][0] ),
    .S0(_02467_),
    .S1(_02468_),
    .X(_02473_));
 sky130_fd_sc_hd__clkbuf_2 _06525_ (.A(_02381_),
    .X(_02474_));
 sky130_fd_sc_hd__buf_4 _06526_ (.A(_02474_),
    .X(_02475_));
 sky130_fd_sc_hd__mux4_1 _06527_ (.A0(\mem[40][0] ),
    .A1(\mem[41][0] ),
    .A2(\mem[42][0] ),
    .A3(\mem[43][0] ),
    .S0(_02457_),
    .S1(_02460_),
    .X(_02476_));
 sky130_fd_sc_hd__or2_1 _06528_ (.A(_02475_),
    .B(_02476_),
    .X(_02477_));
 sky130_fd_sc_hd__buf_2 _06529_ (.A(net4),
    .X(_02478_));
 sky130_fd_sc_hd__buf_4 _06530_ (.A(_02478_),
    .X(_02479_));
 sky130_fd_sc_hd__o211a_1 _06531_ (.A1(_02472_),
    .A2(_02473_),
    .B1(_02477_),
    .C1(_02479_),
    .X(_02480_));
 sky130_fd_sc_hd__or3_4 _06532_ (.A(_02453_),
    .B(_02470_),
    .C(_02480_),
    .X(_02481_));
 sky130_fd_sc_hd__clkbuf_4 _06533_ (.A(_02357_),
    .X(_02482_));
 sky130_fd_sc_hd__nand2_2 _06534_ (.A(_02381_),
    .B(net4),
    .Y(_02483_));
 sky130_fd_sc_hd__buf_6 _06535_ (.A(_02483_),
    .X(_02484_));
 sky130_fd_sc_hd__buf_6 _06536_ (.A(_02484_),
    .X(_02485_));
 sky130_fd_sc_hd__buf_6 _06537_ (.A(_02373_),
    .X(_02486_));
 sky130_fd_sc_hd__buf_6 _06538_ (.A(_02486_),
    .X(_02487_));
 sky130_fd_sc_hd__buf_6 _06539_ (.A(_02459_),
    .X(_02488_));
 sky130_fd_sc_hd__clkbuf_16 _06540_ (.A(_02488_),
    .X(_02489_));
 sky130_fd_sc_hd__mux4_1 _06541_ (.A0(\mem[60][0] ),
    .A1(\mem[61][0] ),
    .A2(\mem[62][0] ),
    .A3(\mem[63][0] ),
    .S0(_02487_),
    .S1(_02489_),
    .X(_02490_));
 sky130_fd_sc_hd__buf_6 _06542_ (.A(_02447_),
    .X(_02491_));
 sky130_fd_sc_hd__buf_6 _06543_ (.A(_02429_),
    .X(_02492_));
 sky130_fd_sc_hd__mux4_1 _06544_ (.A0(\mem[48][0] ),
    .A1(\mem[49][0] ),
    .A2(\mem[50][0] ),
    .A3(\mem[51][0] ),
    .S0(_02491_),
    .S1(_02492_),
    .X(_02493_));
 sky130_fd_sc_hd__or2_1 _06545_ (.A(_02381_),
    .B(net4),
    .X(_02494_));
 sky130_fd_sc_hd__buf_4 _06546_ (.A(_02494_),
    .X(_02495_));
 sky130_fd_sc_hd__clkbuf_8 _06547_ (.A(_02495_),
    .X(_02496_));
 sky130_fd_sc_hd__nand2b_4 _06548_ (.A_N(net4),
    .B(_02381_),
    .Y(_02497_));
 sky130_fd_sc_hd__buf_8 _06549_ (.A(_02497_),
    .X(_02498_));
 sky130_fd_sc_hd__buf_8 _06550_ (.A(_02375_),
    .X(_02499_));
 sky130_fd_sc_hd__mux4_1 _06551_ (.A0(\mem[52][0] ),
    .A1(\mem[53][0] ),
    .A2(\mem[54][0] ),
    .A3(\mem[55][0] ),
    .S0(_02427_),
    .S1(_02499_),
    .X(_02500_));
 sky130_fd_sc_hd__buf_4 _06552_ (.A(_02360_),
    .X(_02501_));
 sky130_fd_sc_hd__buf_8 _06553_ (.A(_02501_),
    .X(_02502_));
 sky130_fd_sc_hd__buf_6 _06554_ (.A(_02375_),
    .X(_02503_));
 sky130_fd_sc_hd__mux4_1 _06555_ (.A0(\mem[56][0] ),
    .A1(\mem[57][0] ),
    .A2(\mem[58][0] ),
    .A3(\mem[59][0] ),
    .S0(_02502_),
    .S1(_02503_),
    .X(_02504_));
 sky130_fd_sc_hd__nand2b_4 _06556_ (.A_N(_02381_),
    .B(net4),
    .Y(_02505_));
 sky130_fd_sc_hd__buf_6 _06557_ (.A(_02505_),
    .X(_02506_));
 sky130_fd_sc_hd__o22a_1 _06558_ (.A1(_02498_),
    .A2(_02500_),
    .B1(_02504_),
    .B2(_02506_),
    .X(_02507_));
 sky130_fd_sc_hd__o221a_2 _06559_ (.A1(_02485_),
    .A2(_02490_),
    .B1(_02493_),
    .B2(_02496_),
    .C1(_02507_),
    .X(_02508_));
 sky130_fd_sc_hd__buf_4 _06560_ (.A(net6),
    .X(_02509_));
 sky130_fd_sc_hd__clkbuf_4 _06561_ (.A(_02509_),
    .X(_02510_));
 sky130_fd_sc_hd__o21a_1 _06562_ (.A1(_02482_),
    .A2(_02508_),
    .B1(_02510_),
    .X(_02511_));
 sky130_fd_sc_hd__a32o_1 _06563_ (.A1(_02356_),
    .A2(_02419_),
    .A3(_02452_),
    .B1(_02481_),
    .B2(_02511_),
    .X(_02512_));
 sky130_fd_sc_hd__buf_2 _06564_ (.A(_02355_),
    .X(_02513_));
 sky130_fd_sc_hd__clkbuf_4 _06565_ (.A(_02357_),
    .X(_02514_));
 sky130_fd_sc_hd__buf_4 _06566_ (.A(_02362_),
    .X(_02515_));
 sky130_fd_sc_hd__clkbuf_4 _06567_ (.A(_02365_),
    .X(_02516_));
 sky130_fd_sc_hd__o21a_1 _06568_ (.A1(\mem[93][0] ),
    .A2(_02515_),
    .B1(_02516_),
    .X(_02517_));
 sky130_fd_sc_hd__buf_4 _06569_ (.A(_02368_),
    .X(_02518_));
 sky130_fd_sc_hd__clkbuf_4 _06570_ (.A(_02371_),
    .X(_02519_));
 sky130_fd_sc_hd__buf_2 _06571_ (.A(_02360_),
    .X(_02520_));
 sky130_fd_sc_hd__buf_2 _06572_ (.A(_02359_),
    .X(_02521_));
 sky130_fd_sc_hd__or3_1 _06573_ (.A(_02520_),
    .B(_02521_),
    .C(\mem[92][0] ),
    .X(_02522_));
 sky130_fd_sc_hd__o221a_1 _06574_ (.A1(\mem[94][0] ),
    .A2(_02518_),
    .B1(_02519_),
    .B2(\mem[95][0] ),
    .C1(_02522_),
    .X(_02523_));
 sky130_fd_sc_hd__buf_4 _06575_ (.A(_02379_),
    .X(_02524_));
 sky130_fd_sc_hd__clkbuf_4 _06576_ (.A(_02382_),
    .X(_02525_));
 sky130_fd_sc_hd__o21a_1 _06577_ (.A1(\mem[80][0] ),
    .A2(_02524_),
    .B1(_02525_),
    .X(_02526_));
 sky130_fd_sc_hd__clkbuf_4 _06578_ (.A(_02361_),
    .X(_02527_));
 sky130_fd_sc_hd__buf_4 _06579_ (.A(_02371_),
    .X(_02528_));
 sky130_fd_sc_hd__clkbuf_4 _06580_ (.A(_02373_),
    .X(_02529_));
 sky130_fd_sc_hd__buf_2 _06581_ (.A(_02359_),
    .X(_02530_));
 sky130_fd_sc_hd__or3b_1 _06582_ (.A(_02529_),
    .B(\mem[82][0] ),
    .C_N(_02530_),
    .X(_02531_));
 sky130_fd_sc_hd__o221a_1 _06583_ (.A1(\mem[81][0] ),
    .A2(_02527_),
    .B1(_02528_),
    .B2(\mem[83][0] ),
    .C1(_02531_),
    .X(_02532_));
 sky130_fd_sc_hd__a22o_1 _06584_ (.A1(_02517_),
    .A2(_02523_),
    .B1(_02526_),
    .B2(_02532_),
    .X(_02533_));
 sky130_fd_sc_hd__buf_4 _06585_ (.A(_02393_),
    .X(_02534_));
 sky130_fd_sc_hd__buf_4 _06586_ (.A(_02379_),
    .X(_02535_));
 sky130_fd_sc_hd__buf_4 _06587_ (.A(_02396_),
    .X(_02536_));
 sky130_fd_sc_hd__o21a_1 _06588_ (.A1(\mem[88][0] ),
    .A2(_02535_),
    .B1(_02536_),
    .X(_02537_));
 sky130_fd_sc_hd__clkbuf_8 _06589_ (.A(_02362_),
    .X(_02538_));
 sky130_fd_sc_hd__buf_4 _06590_ (.A(_02400_),
    .X(_02539_));
 sky130_fd_sc_hd__o22a_1 _06591_ (.A1(\mem[89][0] ),
    .A2(_02538_),
    .B1(_02539_),
    .B2(\mem[91][0] ),
    .X(_02540_));
 sky130_fd_sc_hd__o211a_1 _06592_ (.A1(\mem[90][0] ),
    .A2(_02534_),
    .B1(_02537_),
    .C1(_02540_),
    .X(_02541_));
 sky130_fd_sc_hd__buf_4 _06593_ (.A(_02405_),
    .X(_02542_));
 sky130_fd_sc_hd__buf_4 _06594_ (.A(_02369_),
    .X(_02543_));
 sky130_fd_sc_hd__clkbuf_8 _06595_ (.A(_02408_),
    .X(_02544_));
 sky130_fd_sc_hd__buf_6 _06596_ (.A(_02410_),
    .X(_02545_));
 sky130_fd_sc_hd__buf_4 _06597_ (.A(_02388_),
    .X(_02546_));
 sky130_fd_sc_hd__or3_1 _06598_ (.A(_02545_),
    .B(_02546_),
    .C(\mem[84][0] ),
    .X(_02547_));
 sky130_fd_sc_hd__o221a_1 _06599_ (.A1(\mem[86][0] ),
    .A2(_02543_),
    .B1(_02544_),
    .B2(\mem[87][0] ),
    .C1(_02547_),
    .X(_02548_));
 sky130_fd_sc_hd__buf_4 _06600_ (.A(_02416_),
    .X(_02549_));
 sky130_fd_sc_hd__o211a_1 _06601_ (.A1(\mem[85][0] ),
    .A2(_02542_),
    .B1(_02548_),
    .C1(_02549_),
    .X(_02550_));
 sky130_fd_sc_hd__or4_4 _06602_ (.A(_02514_),
    .B(_02533_),
    .C(_02541_),
    .D(_02550_),
    .X(_02551_));
 sky130_fd_sc_hd__clkbuf_4 _06603_ (.A(_02420_),
    .X(_02552_));
 sky130_fd_sc_hd__clkbuf_4 _06604_ (.A(_02538_),
    .X(_02553_));
 sky130_fd_sc_hd__buf_4 _06605_ (.A(_02369_),
    .X(_02554_));
 sky130_fd_sc_hd__buf_4 _06606_ (.A(_02371_),
    .X(_02555_));
 sky130_fd_sc_hd__buf_2 _06607_ (.A(_02373_),
    .X(_02556_));
 sky130_fd_sc_hd__or3_1 _06608_ (.A(_02556_),
    .B(_02433_),
    .C(\mem[76][0] ),
    .X(_02557_));
 sky130_fd_sc_hd__o221a_1 _06609_ (.A1(\mem[78][0] ),
    .A2(_02554_),
    .B1(_02555_),
    .B2(\mem[79][0] ),
    .C1(_02557_),
    .X(_02558_));
 sky130_fd_sc_hd__clkbuf_4 _06610_ (.A(_02422_),
    .X(_02559_));
 sky130_fd_sc_hd__o211a_1 _06611_ (.A1(\mem[77][0] ),
    .A2(_02553_),
    .B1(_02558_),
    .C1(_02559_),
    .X(_02560_));
 sky130_fd_sc_hd__buf_4 _06612_ (.A(_02393_),
    .X(_02561_));
 sky130_fd_sc_hd__buf_4 _06613_ (.A(_02379_),
    .X(_02562_));
 sky130_fd_sc_hd__clkbuf_4 _06614_ (.A(_02454_),
    .X(_02563_));
 sky130_fd_sc_hd__o21a_1 _06615_ (.A1(\mem[64][0] ),
    .A2(_02562_),
    .B1(_02563_),
    .X(_02564_));
 sky130_fd_sc_hd__buf_4 _06616_ (.A(_02404_),
    .X(_02565_));
 sky130_fd_sc_hd__buf_4 _06617_ (.A(_02400_),
    .X(_02566_));
 sky130_fd_sc_hd__o22a_1 _06618_ (.A1(\mem[65][0] ),
    .A2(_02565_),
    .B1(_02566_),
    .B2(\mem[67][0] ),
    .X(_02567_));
 sky130_fd_sc_hd__o211a_1 _06619_ (.A1(\mem[66][0] ),
    .A2(_02561_),
    .B1(_02564_),
    .C1(_02567_),
    .X(_02568_));
 sky130_fd_sc_hd__clkbuf_4 _06620_ (.A(_02439_),
    .X(_02569_));
 sky130_fd_sc_hd__clkbuf_4 _06621_ (.A(_02378_),
    .X(_02570_));
 sky130_fd_sc_hd__or2_1 _06622_ (.A(\mem[72][0] ),
    .B(_02570_),
    .X(_02571_));
 sky130_fd_sc_hd__buf_6 _06623_ (.A(_02362_),
    .X(_02572_));
 sky130_fd_sc_hd__buf_4 _06624_ (.A(_02408_),
    .X(_02573_));
 sky130_fd_sc_hd__clkbuf_4 _06625_ (.A(_02373_),
    .X(_02574_));
 sky130_fd_sc_hd__buf_2 _06626_ (.A(_02388_),
    .X(_02575_));
 sky130_fd_sc_hd__or3b_1 _06627_ (.A(_02574_),
    .B(\mem[74][0] ),
    .C_N(_02575_),
    .X(_02576_));
 sky130_fd_sc_hd__o221a_1 _06628_ (.A1(\mem[73][0] ),
    .A2(_02572_),
    .B1(_02573_),
    .B2(\mem[75][0] ),
    .C1(_02576_),
    .X(_02577_));
 sky130_fd_sc_hd__buf_2 _06629_ (.A(_02404_),
    .X(_02578_));
 sky130_fd_sc_hd__clkbuf_4 _06630_ (.A(_02415_),
    .X(_02579_));
 sky130_fd_sc_hd__o21a_1 _06631_ (.A1(\mem[69][0] ),
    .A2(_02578_),
    .B1(_02579_),
    .X(_02580_));
 sky130_fd_sc_hd__buf_4 _06632_ (.A(_02369_),
    .X(_02581_));
 sky130_fd_sc_hd__clkbuf_4 _06633_ (.A(_02408_),
    .X(_02582_));
 sky130_fd_sc_hd__clkbuf_4 _06634_ (.A(_02410_),
    .X(_02583_));
 sky130_fd_sc_hd__buf_4 _06635_ (.A(_02459_),
    .X(_02584_));
 sky130_fd_sc_hd__or3_1 _06636_ (.A(_02583_),
    .B(_02584_),
    .C(\mem[68][0] ),
    .X(_02585_));
 sky130_fd_sc_hd__o221a_1 _06637_ (.A1(\mem[70][0] ),
    .A2(_02581_),
    .B1(_02582_),
    .B2(\mem[71][0] ),
    .C1(_02585_),
    .X(_02586_));
 sky130_fd_sc_hd__a32o_1 _06638_ (.A1(_02569_),
    .A2(_02571_),
    .A3(_02577_),
    .B1(_02580_),
    .B2(_02586_),
    .X(_02587_));
 sky130_fd_sc_hd__or4_4 _06639_ (.A(_02552_),
    .B(_02560_),
    .C(_02568_),
    .D(_02587_),
    .X(_02588_));
 sky130_fd_sc_hd__clkbuf_4 _06640_ (.A(_02420_),
    .X(_02589_));
 sky130_fd_sc_hd__buf_6 _06641_ (.A(_02457_),
    .X(_02590_));
 sky130_fd_sc_hd__buf_4 _06642_ (.A(_02460_),
    .X(_02591_));
 sky130_fd_sc_hd__mux4_1 _06643_ (.A0(\mem[100][0] ),
    .A1(\mem[101][0] ),
    .A2(\mem[102][0] ),
    .A3(\mem[103][0] ),
    .S0(_02590_),
    .S1(_02591_),
    .X(_02592_));
 sky130_fd_sc_hd__buf_6 _06644_ (.A(_02374_),
    .X(_02593_));
 sky130_fd_sc_hd__buf_4 _06645_ (.A(_02488_),
    .X(_02594_));
 sky130_fd_sc_hd__mux4_1 _06646_ (.A0(\mem[96][0] ),
    .A1(\mem[97][0] ),
    .A2(\mem[98][0] ),
    .A3(\mem[99][0] ),
    .S0(_02593_),
    .S1(_02594_),
    .X(_02595_));
 sky130_fd_sc_hd__buf_8 _06647_ (.A(_02455_),
    .X(_02596_));
 sky130_fd_sc_hd__a22o_1 _06648_ (.A1(_02450_),
    .A2(_02592_),
    .B1(_02595_),
    .B2(_02596_),
    .X(_02597_));
 sky130_fd_sc_hd__buf_2 _06649_ (.A(_02471_),
    .X(_02598_));
 sky130_fd_sc_hd__clkbuf_4 _06650_ (.A(_02598_),
    .X(_02599_));
 sky130_fd_sc_hd__buf_6 _06651_ (.A(_02457_),
    .X(_02600_));
 sky130_fd_sc_hd__buf_4 _06652_ (.A(_02460_),
    .X(_02601_));
 sky130_fd_sc_hd__mux4_2 _06653_ (.A0(\mem[108][0] ),
    .A1(\mem[109][0] ),
    .A2(\mem[110][0] ),
    .A3(\mem[111][0] ),
    .S0(_02600_),
    .S1(_02601_),
    .X(_02602_));
 sky130_fd_sc_hd__clkbuf_4 _06654_ (.A(_02381_),
    .X(_02603_));
 sky130_fd_sc_hd__buf_4 _06655_ (.A(_02360_),
    .X(_02604_));
 sky130_fd_sc_hd__buf_6 _06656_ (.A(_02459_),
    .X(_02605_));
 sky130_fd_sc_hd__mux4_1 _06657_ (.A0(\mem[104][0] ),
    .A1(\mem[105][0] ),
    .A2(\mem[106][0] ),
    .A3(\mem[107][0] ),
    .S0(_02604_),
    .S1(_02605_),
    .X(_02606_));
 sky130_fd_sc_hd__or2_1 _06658_ (.A(_02603_),
    .B(_02606_),
    .X(_02607_));
 sky130_fd_sc_hd__clkbuf_4 _06659_ (.A(net4),
    .X(_02608_));
 sky130_fd_sc_hd__o211a_1 _06660_ (.A1(_02599_),
    .A2(_02602_),
    .B1(_02607_),
    .C1(_02608_),
    .X(_02609_));
 sky130_fd_sc_hd__or3_2 _06661_ (.A(_02589_),
    .B(_02597_),
    .C(_02609_),
    .X(_02610_));
 sky130_fd_sc_hd__buf_2 _06662_ (.A(_02357_),
    .X(_02611_));
 sky130_fd_sc_hd__buf_4 _06663_ (.A(_02483_),
    .X(_02612_));
 sky130_fd_sc_hd__buf_6 _06664_ (.A(_02486_),
    .X(_02613_));
 sky130_fd_sc_hd__clkbuf_8 _06665_ (.A(_02488_),
    .X(_02614_));
 sky130_fd_sc_hd__mux4_1 _06666_ (.A0(\mem[124][0] ),
    .A1(\mem[125][0] ),
    .A2(\mem[126][0] ),
    .A3(\mem[127][0] ),
    .S0(_02613_),
    .S1(_02614_),
    .X(_02615_));
 sky130_fd_sc_hd__buf_6 _06667_ (.A(_02545_),
    .X(_02616_));
 sky130_fd_sc_hd__buf_6 _06668_ (.A(_02459_),
    .X(_02617_));
 sky130_fd_sc_hd__buf_4 _06669_ (.A(_02617_),
    .X(_02618_));
 sky130_fd_sc_hd__mux4_2 _06670_ (.A0(\mem[112][0] ),
    .A1(\mem[113][0] ),
    .A2(\mem[114][0] ),
    .A3(\mem[115][0] ),
    .S0(_02616_),
    .S1(_02618_),
    .X(_02619_));
 sky130_fd_sc_hd__buf_4 _06671_ (.A(_02495_),
    .X(_02620_));
 sky130_fd_sc_hd__clkbuf_4 _06672_ (.A(_02497_),
    .X(_02621_));
 sky130_fd_sc_hd__clkbuf_8 _06673_ (.A(_02410_),
    .X(_02622_));
 sky130_fd_sc_hd__buf_8 _06674_ (.A(_02521_),
    .X(_02623_));
 sky130_fd_sc_hd__mux4_1 _06675_ (.A0(\mem[116][0] ),
    .A1(\mem[117][0] ),
    .A2(\mem[118][0] ),
    .A3(\mem[119][0] ),
    .S0(_02622_),
    .S1(_02623_),
    .X(_02624_));
 sky130_fd_sc_hd__buf_6 _06676_ (.A(_02410_),
    .X(_02625_));
 sky130_fd_sc_hd__buf_4 _06677_ (.A(_02375_),
    .X(_02626_));
 sky130_fd_sc_hd__mux4_1 _06678_ (.A0(\mem[120][0] ),
    .A1(\mem[121][0] ),
    .A2(\mem[122][0] ),
    .A3(\mem[123][0] ),
    .S0(_02625_),
    .S1(_02626_),
    .X(_02627_));
 sky130_fd_sc_hd__clkbuf_4 _06679_ (.A(_02505_),
    .X(_02628_));
 sky130_fd_sc_hd__o22a_1 _06680_ (.A1(_02621_),
    .A2(_02624_),
    .B1(_02627_),
    .B2(_02628_),
    .X(_02629_));
 sky130_fd_sc_hd__o221a_1 _06681_ (.A1(_02612_),
    .A2(_02615_),
    .B1(_02619_),
    .B2(_02620_),
    .C1(_02629_),
    .X(_02630_));
 sky130_fd_sc_hd__buf_2 _06682_ (.A(_02509_),
    .X(_02631_));
 sky130_fd_sc_hd__o21a_1 _06683_ (.A1(_02611_),
    .A2(_02630_),
    .B1(_02631_),
    .X(_02632_));
 sky130_fd_sc_hd__a32o_1 _06684_ (.A1(_02513_),
    .A2(_02551_),
    .A3(_02588_),
    .B1(_02610_),
    .B2(_02632_),
    .X(_02633_));
 sky130_fd_sc_hd__clkbuf_4 _06685_ (.A(net7),
    .X(_02634_));
 sky130_fd_sc_hd__clkbuf_4 _06686_ (.A(_02634_),
    .X(_02635_));
 sky130_fd_sc_hd__mux2_1 _06687_ (.A0(_02512_),
    .A1(_02633_),
    .S(_02635_),
    .X(_02636_));
 sky130_fd_sc_hd__clkbuf_1 _06688_ (.A(_02636_),
    .X(_00000_));
 sky130_fd_sc_hd__clkbuf_4 _06689_ (.A(_02510_),
    .X(_02637_));
 sky130_fd_sc_hd__buf_8 _06690_ (.A(_02482_),
    .X(_02638_));
 sky130_fd_sc_hd__buf_4 _06691_ (.A(_02404_),
    .X(_02639_));
 sky130_fd_sc_hd__clkbuf_8 _06692_ (.A(_02639_),
    .X(_02640_));
 sky130_fd_sc_hd__clkbuf_8 _06693_ (.A(_02422_),
    .X(_02641_));
 sky130_fd_sc_hd__o21a_1 _06694_ (.A1(\mem[93][1] ),
    .A2(_02640_),
    .B1(_02641_),
    .X(_02642_));
 sky130_fd_sc_hd__buf_4 _06695_ (.A(_02393_),
    .X(_02643_));
 sky130_fd_sc_hd__buf_6 _06696_ (.A(_02386_),
    .X(_02644_));
 sky130_fd_sc_hd__buf_6 _06697_ (.A(_02501_),
    .X(_02645_));
 sky130_fd_sc_hd__buf_6 _06698_ (.A(_02645_),
    .X(_02646_));
 sky130_fd_sc_hd__or3_1 _06699_ (.A(_02646_),
    .B(_02489_),
    .C(\mem[92][1] ),
    .X(_02647_));
 sky130_fd_sc_hd__o221a_1 _06700_ (.A1(\mem[94][1] ),
    .A2(_02643_),
    .B1(_02644_),
    .B2(\mem[95][1] ),
    .C1(_02647_),
    .X(_02648_));
 sky130_fd_sc_hd__buf_4 _06701_ (.A(_02379_),
    .X(_02649_));
 sky130_fd_sc_hd__buf_4 _06702_ (.A(_02649_),
    .X(_02650_));
 sky130_fd_sc_hd__buf_4 _06703_ (.A(_02454_),
    .X(_02651_));
 sky130_fd_sc_hd__buf_6 _06704_ (.A(_02651_),
    .X(_02652_));
 sky130_fd_sc_hd__o21a_1 _06705_ (.A1(\mem[80][1] ),
    .A2(_02650_),
    .B1(_02652_),
    .X(_02653_));
 sky130_fd_sc_hd__buf_6 _06706_ (.A(_02639_),
    .X(_02654_));
 sky130_fd_sc_hd__buf_4 _06707_ (.A(_02442_),
    .X(_02655_));
 sky130_fd_sc_hd__buf_6 _06708_ (.A(_02467_),
    .X(_02656_));
 sky130_fd_sc_hd__or3b_1 _06709_ (.A(_02656_),
    .B(\mem[82][1] ),
    .C_N(_02492_),
    .X(_02657_));
 sky130_fd_sc_hd__o221a_1 _06710_ (.A1(\mem[81][1] ),
    .A2(_02654_),
    .B1(_02655_),
    .B2(\mem[83][1] ),
    .C1(_02657_),
    .X(_02658_));
 sky130_fd_sc_hd__a22o_1 _06711_ (.A1(_02642_),
    .A2(_02648_),
    .B1(_02653_),
    .B2(_02658_),
    .X(_02659_));
 sky130_fd_sc_hd__clkbuf_8 _06712_ (.A(_02445_),
    .X(_02660_));
 sky130_fd_sc_hd__buf_6 _06713_ (.A(_02660_),
    .X(_02661_));
 sky130_fd_sc_hd__buf_6 _06714_ (.A(_02439_),
    .X(_02662_));
 sky130_fd_sc_hd__o21a_1 _06715_ (.A1(\mem[88][1] ),
    .A2(_02650_),
    .B1(_02662_),
    .X(_02663_));
 sky130_fd_sc_hd__buf_6 _06716_ (.A(_02408_),
    .X(_02664_));
 sky130_fd_sc_hd__buf_4 _06717_ (.A(_02664_),
    .X(_02665_));
 sky130_fd_sc_hd__buf_6 _06718_ (.A(_02665_),
    .X(_02666_));
 sky130_fd_sc_hd__o22a_1 _06719_ (.A1(\mem[89][1] ),
    .A2(_02640_),
    .B1(_02666_),
    .B2(\mem[91][1] ),
    .X(_02667_));
 sky130_fd_sc_hd__o211a_1 _06720_ (.A1(\mem[90][1] ),
    .A2(_02661_),
    .B1(_02663_),
    .C1(_02667_),
    .X(_02668_));
 sky130_fd_sc_hd__buf_6 _06721_ (.A(_02406_),
    .X(_02669_));
 sky130_fd_sc_hd__buf_6 _06722_ (.A(_02373_),
    .X(_02670_));
 sky130_fd_sc_hd__buf_12 _06723_ (.A(_02670_),
    .X(_02671_));
 sky130_fd_sc_hd__clkbuf_16 _06724_ (.A(_02671_),
    .X(_02672_));
 sky130_fd_sc_hd__buf_6 _06725_ (.A(_02375_),
    .X(_02673_));
 sky130_fd_sc_hd__buf_6 _06726_ (.A(_02673_),
    .X(_02674_));
 sky130_fd_sc_hd__or3_1 _06727_ (.A(_02672_),
    .B(_02674_),
    .C(\mem[84][1] ),
    .X(_02675_));
 sky130_fd_sc_hd__o221a_1 _06728_ (.A1(\mem[86][1] ),
    .A2(_02643_),
    .B1(_02655_),
    .B2(\mem[87][1] ),
    .C1(_02675_),
    .X(_02676_));
 sky130_fd_sc_hd__buf_6 _06729_ (.A(_02417_),
    .X(_02677_));
 sky130_fd_sc_hd__o211a_1 _06730_ (.A1(\mem[85][1] ),
    .A2(_02669_),
    .B1(_02676_),
    .C1(_02677_),
    .X(_02678_));
 sky130_fd_sc_hd__nor4_4 _06731_ (.A(_02638_),
    .B(_02659_),
    .C(_02668_),
    .D(_02678_),
    .Y(_02679_));
 sky130_fd_sc_hd__buf_6 _06732_ (.A(_02453_),
    .X(_02680_));
 sky130_fd_sc_hd__buf_12 _06733_ (.A(_02467_),
    .X(_02681_));
 sky130_fd_sc_hd__buf_6 _06734_ (.A(_02499_),
    .X(_02682_));
 sky130_fd_sc_hd__or3_1 _06735_ (.A(_02681_),
    .B(_02682_),
    .C(\mem[76][1] ),
    .X(_02683_));
 sky130_fd_sc_hd__o221a_1 _06736_ (.A1(\mem[78][1] ),
    .A2(_02643_),
    .B1(_02655_),
    .B2(\mem[79][1] ),
    .C1(_02683_),
    .X(_02684_));
 sky130_fd_sc_hd__o211a_1 _06737_ (.A1(\mem[77][1] ),
    .A2(_02669_),
    .B1(_02684_),
    .C1(_02641_),
    .X(_02685_));
 sky130_fd_sc_hd__o21a_1 _06738_ (.A1(\mem[64][1] ),
    .A2(_02650_),
    .B1(_02652_),
    .X(_02686_));
 sky130_fd_sc_hd__o22a_1 _06739_ (.A1(\mem[65][1] ),
    .A2(_02640_),
    .B1(_02666_),
    .B2(\mem[67][1] ),
    .X(_02687_));
 sky130_fd_sc_hd__o211a_1 _06740_ (.A1(\mem[66][1] ),
    .A2(_02661_),
    .B1(_02686_),
    .C1(_02687_),
    .X(_02688_));
 sky130_fd_sc_hd__or2_1 _06741_ (.A(\mem[72][1] ),
    .B(_02650_),
    .X(_02689_));
 sky130_fd_sc_hd__or3b_1 _06742_ (.A(_02672_),
    .B(\mem[74][1] ),
    .C_N(_02682_),
    .X(_02690_));
 sky130_fd_sc_hd__o221a_1 _06743_ (.A1(\mem[73][1] ),
    .A2(_02654_),
    .B1(_02655_),
    .B2(\mem[75][1] ),
    .C1(_02690_),
    .X(_02691_));
 sky130_fd_sc_hd__o21a_1 _06744_ (.A1(\mem[69][1] ),
    .A2(_02669_),
    .B1(_02677_),
    .X(_02692_));
 sky130_fd_sc_hd__buf_8 _06745_ (.A(_02487_),
    .X(_02693_));
 sky130_fd_sc_hd__or3_1 _06746_ (.A(_02693_),
    .B(_02674_),
    .C(\mem[68][1] ),
    .X(_02694_));
 sky130_fd_sc_hd__o221a_1 _06747_ (.A1(\mem[70][1] ),
    .A2(_02661_),
    .B1(_02666_),
    .B2(\mem[71][1] ),
    .C1(_02694_),
    .X(_02695_));
 sky130_fd_sc_hd__a32o_1 _06748_ (.A1(_02662_),
    .A2(_02689_),
    .A3(_02691_),
    .B1(_02692_),
    .B2(_02695_),
    .X(_02696_));
 sky130_fd_sc_hd__nor4_4 _06749_ (.A(_02680_),
    .B(_02685_),
    .C(_02688_),
    .D(_02696_),
    .Y(_02697_));
 sky130_fd_sc_hd__buf_6 _06750_ (.A(_02646_),
    .X(_02698_));
 sky130_fd_sc_hd__buf_8 _06751_ (.A(_02674_),
    .X(_02699_));
 sky130_fd_sc_hd__mux4_1 _06752_ (.A0(\mem[124][1] ),
    .A1(\mem[125][1] ),
    .A2(\mem[126][1] ),
    .A3(\mem[127][1] ),
    .S0(_02698_),
    .S1(_02699_),
    .X(_02700_));
 sky130_fd_sc_hd__mux4_1 _06753_ (.A0(\mem[112][1] ),
    .A1(\mem[113][1] ),
    .A2(\mem[114][1] ),
    .A3(\mem[115][1] ),
    .S0(_02698_),
    .S1(_02699_),
    .X(_02701_));
 sky130_fd_sc_hd__buf_8 _06754_ (.A(_02497_),
    .X(_02702_));
 sky130_fd_sc_hd__buf_8 _06755_ (.A(_02488_),
    .X(_02703_));
 sky130_fd_sc_hd__buf_8 _06756_ (.A(_02703_),
    .X(_02704_));
 sky130_fd_sc_hd__mux4_1 _06757_ (.A0(\mem[116][1] ),
    .A1(\mem[117][1] ),
    .A2(\mem[118][1] ),
    .A3(\mem[119][1] ),
    .S0(_02681_),
    .S1(_02704_),
    .X(_02705_));
 sky130_fd_sc_hd__mux4_1 _06758_ (.A0(\mem[120][1] ),
    .A1(\mem[121][1] ),
    .A2(\mem[122][1] ),
    .A3(\mem[123][1] ),
    .S0(_02672_),
    .S1(_02704_),
    .X(_02706_));
 sky130_fd_sc_hd__buf_6 _06759_ (.A(_02505_),
    .X(_02707_));
 sky130_fd_sc_hd__o22a_1 _06760_ (.A1(_02702_),
    .A2(_02705_),
    .B1(_02706_),
    .B2(_02707_),
    .X(_02708_));
 sky130_fd_sc_hd__o221a_1 _06761_ (.A1(_02485_),
    .A2(_02700_),
    .B1(_02701_),
    .B2(_02496_),
    .C1(_02708_),
    .X(_02709_));
 sky130_fd_sc_hd__nor2_1 _06762_ (.A(_02638_),
    .B(_02709_),
    .Y(_02710_));
 sky130_fd_sc_hd__buf_6 _06763_ (.A(_02646_),
    .X(_02711_));
 sky130_fd_sc_hd__clkbuf_8 _06764_ (.A(_02682_),
    .X(_02712_));
 sky130_fd_sc_hd__mux4_1 _06765_ (.A0(\mem[96][1] ),
    .A1(\mem[97][1] ),
    .A2(\mem[98][1] ),
    .A3(\mem[99][1] ),
    .S0(_02711_),
    .S1(_02712_),
    .X(_02713_));
 sky130_fd_sc_hd__mux4_1 _06766_ (.A0(\mem[100][1] ),
    .A1(\mem[101][1] ),
    .A2(\mem[102][1] ),
    .A3(\mem[103][1] ),
    .S0(_02711_),
    .S1(_02699_),
    .X(_02714_));
 sky130_fd_sc_hd__a22o_1 _06767_ (.A1(_02652_),
    .A2(_02713_),
    .B1(_02714_),
    .B2(_02677_),
    .X(_02715_));
 sky130_fd_sc_hd__buf_4 _06768_ (.A(_02472_),
    .X(_02716_));
 sky130_fd_sc_hd__mux4_1 _06769_ (.A0(\mem[108][1] ),
    .A1(\mem[109][1] ),
    .A2(\mem[110][1] ),
    .A3(\mem[111][1] ),
    .S0(_02711_),
    .S1(_02712_),
    .X(_02717_));
 sky130_fd_sc_hd__clkbuf_4 _06770_ (.A(_02475_),
    .X(_02718_));
 sky130_fd_sc_hd__mux4_1 _06771_ (.A0(\mem[104][1] ),
    .A1(\mem[105][1] ),
    .A2(\mem[106][1] ),
    .A3(\mem[107][1] ),
    .S0(_02646_),
    .S1(_02674_),
    .X(_02719_));
 sky130_fd_sc_hd__or2_1 _06772_ (.A(_02718_),
    .B(_02719_),
    .X(_02720_));
 sky130_fd_sc_hd__clkbuf_4 _06773_ (.A(_02478_),
    .X(_02721_));
 sky130_fd_sc_hd__o211a_1 _06774_ (.A1(_02716_),
    .A2(_02717_),
    .B1(_02720_),
    .C1(_02721_),
    .X(_02722_));
 sky130_fd_sc_hd__o31ai_1 _06775_ (.A1(_02680_),
    .A2(_02715_),
    .A3(_02722_),
    .B1(_02637_),
    .Y(_02723_));
 sky130_fd_sc_hd__o32a_1 _06776_ (.A1(_02637_),
    .A2(_02679_),
    .A3(_02697_),
    .B1(_02710_),
    .B2(_02723_),
    .X(_02724_));
 sky130_fd_sc_hd__nor2_1 _06777_ (.A(_02638_),
    .B(_02637_),
    .Y(_02725_));
 sky130_fd_sc_hd__buf_6 _06778_ (.A(_02411_),
    .X(_02726_));
 sky130_fd_sc_hd__or3_1 _06779_ (.A(_02726_),
    .B(_02430_),
    .C(\mem[28][1] ),
    .X(_02727_));
 sky130_fd_sc_hd__o221a_1 _06780_ (.A1(\mem[30][1] ),
    .A2(_02660_),
    .B1(_02665_),
    .B2(\mem[31][1] ),
    .C1(_02727_),
    .X(_02728_));
 sky130_fd_sc_hd__o211a_1 _06781_ (.A1(\mem[29][1] ),
    .A2(_02669_),
    .B1(_02728_),
    .C1(_02641_),
    .X(_02729_));
 sky130_fd_sc_hd__o21a_1 _06782_ (.A1(\mem[16][1] ),
    .A2(_02649_),
    .B1(_02651_),
    .X(_02730_));
 sky130_fd_sc_hd__o22a_1 _06783_ (.A1(\mem[17][1] ),
    .A2(_02406_),
    .B1(_02644_),
    .B2(\mem[19][1] ),
    .X(_02731_));
 sky130_fd_sc_hd__o211a_1 _06784_ (.A1(\mem[18][1] ),
    .A2(_02661_),
    .B1(_02730_),
    .C1(_02731_),
    .X(_02732_));
 sky130_fd_sc_hd__or2_1 _06785_ (.A(\mem[24][1] ),
    .B(_02649_),
    .X(_02733_));
 sky130_fd_sc_hd__or3b_1 _06786_ (.A(_02671_),
    .B(\mem[26][1] ),
    .C_N(_02673_),
    .X(_02734_));
 sky130_fd_sc_hd__o221a_1 _06787_ (.A1(\mem[25][1] ),
    .A2(_02639_),
    .B1(_02665_),
    .B2(\mem[27][1] ),
    .C1(_02734_),
    .X(_02735_));
 sky130_fd_sc_hd__buf_6 _06788_ (.A(_02362_),
    .X(_02736_));
 sky130_fd_sc_hd__buf_8 _06789_ (.A(_02736_),
    .X(_02737_));
 sky130_fd_sc_hd__o21a_1 _06790_ (.A1(\mem[21][1] ),
    .A2(_02737_),
    .B1(_02450_),
    .X(_02738_));
 sky130_fd_sc_hd__or3_1 _06791_ (.A(_02491_),
    .B(_02430_),
    .C(\mem[20][1] ),
    .X(_02739_));
 sky130_fd_sc_hd__o221a_1 _06792_ (.A1(\mem[22][1] ),
    .A2(_02660_),
    .B1(_02665_),
    .B2(\mem[23][1] ),
    .C1(_02739_),
    .X(_02740_));
 sky130_fd_sc_hd__a32o_1 _06793_ (.A1(_02662_),
    .A2(_02733_),
    .A3(_02735_),
    .B1(_02738_),
    .B2(_02740_),
    .X(_02741_));
 sky130_fd_sc_hd__or3_1 _06794_ (.A(_02729_),
    .B(_02732_),
    .C(_02741_),
    .X(_02742_));
 sky130_fd_sc_hd__buf_8 _06795_ (.A(_02601_),
    .X(_02743_));
 sky130_fd_sc_hd__mux4_1 _06796_ (.A0(\mem[8][1] ),
    .A1(\mem[9][1] ),
    .A2(\mem[10][1] ),
    .A3(\mem[11][1] ),
    .S0(_02646_),
    .S1(_02743_),
    .X(_02744_));
 sky130_fd_sc_hd__or2_1 _06797_ (.A(_02718_),
    .B(_02744_),
    .X(_02745_));
 sky130_fd_sc_hd__buf_4 _06798_ (.A(_02617_),
    .X(_02746_));
 sky130_fd_sc_hd__buf_4 _06799_ (.A(_02746_),
    .X(_02747_));
 sky130_fd_sc_hd__buf_4 _06800_ (.A(_02747_),
    .X(_02748_));
 sky130_fd_sc_hd__clkbuf_16 _06801_ (.A(_02428_),
    .X(_02749_));
 sky130_fd_sc_hd__mux2_1 _06802_ (.A0(\mem[14][1] ),
    .A1(\mem[15][1] ),
    .S(_02749_),
    .X(_02750_));
 sky130_fd_sc_hd__mux2_1 _06803_ (.A0(\mem[12][1] ),
    .A1(\mem[13][1] ),
    .S(_02428_),
    .X(_02751_));
 sky130_fd_sc_hd__and2b_1 _06804_ (.A_N(_02747_),
    .B(_02751_),
    .X(_02752_));
 sky130_fd_sc_hd__a211o_1 _06805_ (.A1(_02748_),
    .A2(_02750_),
    .B1(_02752_),
    .C1(_02716_),
    .X(_02753_));
 sky130_fd_sc_hd__mux2_2 _06806_ (.A0(\mem[6][1] ),
    .A1(\mem[7][1] ),
    .S(_02749_),
    .X(_02754_));
 sky130_fd_sc_hd__mux2_1 _06807_ (.A0(\mem[4][1] ),
    .A1(\mem[5][1] ),
    .S(_02428_),
    .X(_02755_));
 sky130_fd_sc_hd__and2b_1 _06808_ (.A_N(_02712_),
    .B(_02755_),
    .X(_02756_));
 sky130_fd_sc_hd__a211o_1 _06809_ (.A1(_02748_),
    .A2(_02754_),
    .B1(_02756_),
    .C1(_02716_),
    .X(_02757_));
 sky130_fd_sc_hd__mux4_1 _06810_ (.A0(\mem[0][1] ),
    .A1(\mem[1][1] ),
    .A2(\mem[2][1] ),
    .A3(\mem[3][1] ),
    .S0(_02693_),
    .S1(_02704_),
    .X(_02758_));
 sky130_fd_sc_hd__o21ba_1 _06811_ (.A1(_02718_),
    .A2(_02758_),
    .B1_N(_02721_),
    .X(_02759_));
 sky130_fd_sc_hd__a32o_1 _06812_ (.A1(_02721_),
    .A2(_02745_),
    .A3(_02753_),
    .B1(_02757_),
    .B2(_02759_),
    .X(_02760_));
 sky130_fd_sc_hd__nor2_1 _06813_ (.A(_02680_),
    .B(_02510_),
    .Y(_02761_));
 sky130_fd_sc_hd__a221o_1 _06814_ (.A1(_02725_),
    .A2(_02742_),
    .B1(_02760_),
    .B2(_02761_),
    .C1(_02634_),
    .X(_02762_));
 sky130_fd_sc_hd__mux4_1 _06815_ (.A0(\mem[60][1] ),
    .A1(\mem[61][1] ),
    .A2(\mem[62][1] ),
    .A3(\mem[63][1] ),
    .S0(_02698_),
    .S1(_02748_),
    .X(_02763_));
 sky130_fd_sc_hd__mux4_1 _06816_ (.A0(\mem[48][1] ),
    .A1(\mem[49][1] ),
    .A2(\mem[50][1] ),
    .A3(\mem[51][1] ),
    .S0(_02698_),
    .S1(_02748_),
    .X(_02764_));
 sky130_fd_sc_hd__mux4_1 _06817_ (.A0(\mem[52][1] ),
    .A1(\mem[53][1] ),
    .A2(\mem[54][1] ),
    .A3(\mem[55][1] ),
    .S0(_02693_),
    .S1(_02747_),
    .X(_02765_));
 sky130_fd_sc_hd__mux4_1 _06818_ (.A0(\mem[56][1] ),
    .A1(\mem[57][1] ),
    .A2(\mem[58][1] ),
    .A3(\mem[59][1] ),
    .S0(_02749_),
    .S1(_02747_),
    .X(_02766_));
 sky130_fd_sc_hd__o22a_1 _06819_ (.A1(_02702_),
    .A2(_02765_),
    .B1(_02766_),
    .B2(_02707_),
    .X(_02767_));
 sky130_fd_sc_hd__o221a_1 _06820_ (.A1(_02485_),
    .A2(_02763_),
    .B1(_02764_),
    .B2(_02496_),
    .C1(_02767_),
    .X(_02768_));
 sky130_fd_sc_hd__mux4_1 _06821_ (.A0(\mem[32][1] ),
    .A1(\mem[33][1] ),
    .A2(\mem[34][1] ),
    .A3(\mem[35][1] ),
    .S0(_02656_),
    .S1(_02743_),
    .X(_02769_));
 sky130_fd_sc_hd__mux4_1 _06822_ (.A0(\mem[36][1] ),
    .A1(\mem[37][1] ),
    .A2(\mem[38][1] ),
    .A3(\mem[39][1] ),
    .S0(_02672_),
    .S1(_02704_),
    .X(_02770_));
 sky130_fd_sc_hd__a22o_1 _06823_ (.A1(_02652_),
    .A2(_02769_),
    .B1(_02770_),
    .B2(_02677_),
    .X(_02771_));
 sky130_fd_sc_hd__mux4_1 _06824_ (.A0(\mem[44][1] ),
    .A1(\mem[45][1] ),
    .A2(\mem[46][1] ),
    .A3(\mem[47][1] ),
    .S0(_02681_),
    .S1(_02743_),
    .X(_02772_));
 sky130_fd_sc_hd__mux4_1 _06825_ (.A0(\mem[40][1] ),
    .A1(\mem[41][1] ),
    .A2(\mem[42][1] ),
    .A3(\mem[43][1] ),
    .S0(_02645_),
    .S1(_02430_),
    .X(_02773_));
 sky130_fd_sc_hd__or2_1 _06826_ (.A(_02718_),
    .B(_02773_),
    .X(_02774_));
 sky130_fd_sc_hd__o211a_1 _06827_ (.A1(_02716_),
    .A2(_02772_),
    .B1(_02774_),
    .C1(_02721_),
    .X(_02775_));
 sky130_fd_sc_hd__or3_1 _06828_ (.A(_02680_),
    .B(_02771_),
    .C(_02775_),
    .X(_02776_));
 sky130_fd_sc_hd__o211a_1 _06829_ (.A1(_02638_),
    .A2(_02768_),
    .B1(_02776_),
    .C1(_02637_),
    .X(_02777_));
 sky130_fd_sc_hd__o2bb2a_1 _06830_ (.A1_N(_02635_),
    .A2_N(_02724_),
    .B1(_02762_),
    .B2(_02777_),
    .X(_00007_));
 sky130_fd_sc_hd__o21a_1 _06831_ (.A1(\mem[29][2] ),
    .A2(_02363_),
    .B1(_02366_),
    .X(_02778_));
 sky130_fd_sc_hd__clkbuf_4 _06832_ (.A(_02388_),
    .X(_02779_));
 sky130_fd_sc_hd__or3_1 _06833_ (.A(_02374_),
    .B(_02779_),
    .C(\mem[28][2] ),
    .X(_02780_));
 sky130_fd_sc_hd__o221a_1 _06834_ (.A1(\mem[30][2] ),
    .A2(_02370_),
    .B1(_02372_),
    .B2(\mem[31][2] ),
    .C1(_02780_),
    .X(_02781_));
 sky130_fd_sc_hd__o21a_1 _06835_ (.A1(\mem[16][2] ),
    .A2(_02380_),
    .B1(_02383_),
    .X(_02782_));
 sky130_fd_sc_hd__clkbuf_4 _06836_ (.A(_02359_),
    .X(_02783_));
 sky130_fd_sc_hd__or3b_1 _06837_ (.A(_02387_),
    .B(\mem[18][2] ),
    .C_N(_02783_),
    .X(_02784_));
 sky130_fd_sc_hd__o221a_1 _06838_ (.A1(\mem[17][2] ),
    .A2(_02385_),
    .B1(_02386_),
    .B2(\mem[19][2] ),
    .C1(_02784_),
    .X(_02785_));
 sky130_fd_sc_hd__a22o_1 _06839_ (.A1(_02778_),
    .A2(_02781_),
    .B1(_02782_),
    .B2(_02785_),
    .X(_02786_));
 sky130_fd_sc_hd__buf_4 _06840_ (.A(_02393_),
    .X(_02787_));
 sky130_fd_sc_hd__buf_4 _06841_ (.A(_02379_),
    .X(_02788_));
 sky130_fd_sc_hd__o21a_1 _06842_ (.A1(\mem[24][2] ),
    .A2(_02788_),
    .B1(_02397_),
    .X(_02789_));
 sky130_fd_sc_hd__buf_4 _06843_ (.A(_02362_),
    .X(_02790_));
 sky130_fd_sc_hd__o22a_1 _06844_ (.A1(\mem[25][2] ),
    .A2(_02790_),
    .B1(_02401_),
    .B2(\mem[27][2] ),
    .X(_02791_));
 sky130_fd_sc_hd__o211a_1 _06845_ (.A1(\mem[26][2] ),
    .A2(_02787_),
    .B1(_02789_),
    .C1(_02791_),
    .X(_02792_));
 sky130_fd_sc_hd__clkbuf_4 _06846_ (.A(_02410_),
    .X(_02793_));
 sky130_fd_sc_hd__or3_1 _06847_ (.A(_02793_),
    .B(_02412_),
    .C(\mem[20][2] ),
    .X(_02794_));
 sky130_fd_sc_hd__o221a_1 _06848_ (.A1(\mem[22][2] ),
    .A2(_02407_),
    .B1(_02409_),
    .B2(\mem[23][2] ),
    .C1(_02794_),
    .X(_02795_));
 sky130_fd_sc_hd__o211a_1 _06849_ (.A1(\mem[21][2] ),
    .A2(_02406_),
    .B1(_02795_),
    .C1(_02417_),
    .X(_02796_));
 sky130_fd_sc_hd__or4_2 _06850_ (.A(_02358_),
    .B(_02786_),
    .C(_02792_),
    .D(_02796_),
    .X(_02797_));
 sky130_fd_sc_hd__clkbuf_2 _06851_ (.A(_02420_),
    .X(_02798_));
 sky130_fd_sc_hd__clkbuf_4 _06852_ (.A(_02399_),
    .X(_02799_));
 sky130_fd_sc_hd__clkbuf_8 _06853_ (.A(_02369_),
    .X(_02800_));
 sky130_fd_sc_hd__buf_4 _06854_ (.A(_02408_),
    .X(_02801_));
 sky130_fd_sc_hd__clkbuf_4 _06855_ (.A(_02373_),
    .X(_02802_));
 sky130_fd_sc_hd__clkbuf_4 _06856_ (.A(_02388_),
    .X(_02803_));
 sky130_fd_sc_hd__or3_1 _06857_ (.A(_02802_),
    .B(_02803_),
    .C(\mem[12][2] ),
    .X(_02804_));
 sky130_fd_sc_hd__o221a_1 _06858_ (.A1(\mem[14][2] ),
    .A2(_02800_),
    .B1(_02801_),
    .B2(\mem[15][2] ),
    .C1(_02804_),
    .X(_02805_));
 sky130_fd_sc_hd__clkbuf_4 _06859_ (.A(_02422_),
    .X(_02806_));
 sky130_fd_sc_hd__o211a_1 _06860_ (.A1(\mem[13][2] ),
    .A2(_02799_),
    .B1(_02805_),
    .C1(_02806_),
    .X(_02807_));
 sky130_fd_sc_hd__o21a_1 _06861_ (.A1(\mem[0][2] ),
    .A2(_02438_),
    .B1(_02455_),
    .X(_02808_));
 sky130_fd_sc_hd__o22a_1 _06862_ (.A1(\mem[1][2] ),
    .A2(_02441_),
    .B1(_02442_),
    .B2(\mem[3][2] ),
    .X(_02809_));
 sky130_fd_sc_hd__o211a_1 _06863_ (.A1(\mem[2][2] ),
    .A2(_02437_),
    .B1(_02808_),
    .C1(_02809_),
    .X(_02810_));
 sky130_fd_sc_hd__clkbuf_4 _06864_ (.A(_02439_),
    .X(_02811_));
 sky130_fd_sc_hd__buf_4 _06865_ (.A(_02378_),
    .X(_02812_));
 sky130_fd_sc_hd__or2_1 _06866_ (.A(\mem[8][2] ),
    .B(_02812_),
    .X(_02813_));
 sky130_fd_sc_hd__clkbuf_8 _06867_ (.A(_02408_),
    .X(_02814_));
 sky130_fd_sc_hd__buf_4 _06868_ (.A(_02373_),
    .X(_02815_));
 sky130_fd_sc_hd__buf_2 _06869_ (.A(_02388_),
    .X(_02816_));
 sky130_fd_sc_hd__or3b_1 _06870_ (.A(_02815_),
    .B(\mem[10][2] ),
    .C_N(_02816_),
    .X(_02817_));
 sky130_fd_sc_hd__o221a_1 _06871_ (.A1(\mem[9][2] ),
    .A2(_02736_),
    .B1(_02814_),
    .B2(\mem[11][2] ),
    .C1(_02817_),
    .X(_02818_));
 sky130_fd_sc_hd__clkbuf_4 _06872_ (.A(_02404_),
    .X(_02819_));
 sky130_fd_sc_hd__o21a_1 _06873_ (.A1(\mem[5][2] ),
    .A2(_02819_),
    .B1(_02416_),
    .X(_02820_));
 sky130_fd_sc_hd__or3_1 _06874_ (.A(_02447_),
    .B(_02429_),
    .C(\mem[4][2] ),
    .X(_02821_));
 sky130_fd_sc_hd__o221a_2 _06875_ (.A1(\mem[6][2] ),
    .A2(_02445_),
    .B1(_02446_),
    .B2(\mem[7][2] ),
    .C1(_02821_),
    .X(_02822_));
 sky130_fd_sc_hd__a32o_1 _06876_ (.A1(_02811_),
    .A2(_02813_),
    .A3(_02818_),
    .B1(_02820_),
    .B2(_02822_),
    .X(_02823_));
 sky130_fd_sc_hd__or4_1 _06877_ (.A(_02798_),
    .B(_02807_),
    .C(_02810_),
    .D(_02823_),
    .X(_02824_));
 sky130_fd_sc_hd__buf_4 _06878_ (.A(_02416_),
    .X(_02825_));
 sky130_fd_sc_hd__buf_6 _06879_ (.A(_02457_),
    .X(_02826_));
 sky130_fd_sc_hd__mux4_1 _06880_ (.A0(\mem[36][2] ),
    .A1(\mem[37][2] ),
    .A2(\mem[38][2] ),
    .A3(\mem[39][2] ),
    .S0(_02826_),
    .S1(_02461_),
    .X(_02827_));
 sky130_fd_sc_hd__mux4_1 _06881_ (.A0(\mem[32][2] ),
    .A1(\mem[33][2] ),
    .A2(\mem[34][2] ),
    .A3(\mem[35][2] ),
    .S0(_02671_),
    .S1(_02703_),
    .X(_02828_));
 sky130_fd_sc_hd__a22o_1 _06882_ (.A1(_02825_),
    .A2(_02827_),
    .B1(_02828_),
    .B2(_02596_),
    .X(_02829_));
 sky130_fd_sc_hd__mux4_1 _06883_ (.A0(\mem[44][2] ),
    .A1(\mem[45][2] ),
    .A2(\mem[46][2] ),
    .A3(\mem[47][2] ),
    .S0(_02467_),
    .S1(_02468_),
    .X(_02830_));
 sky130_fd_sc_hd__mux4_1 _06884_ (.A0(\mem[40][2] ),
    .A1(\mem[41][2] ),
    .A2(\mem[42][2] ),
    .A3(\mem[43][2] ),
    .S0(_02457_),
    .S1(_02460_),
    .X(_02831_));
 sky130_fd_sc_hd__or2_1 _06885_ (.A(_02475_),
    .B(_02831_),
    .X(_02832_));
 sky130_fd_sc_hd__o211a_1 _06886_ (.A1(_02472_),
    .A2(_02830_),
    .B1(_02832_),
    .C1(_02479_),
    .X(_02833_));
 sky130_fd_sc_hd__or3_2 _06887_ (.A(_02453_),
    .B(_02829_),
    .C(_02833_),
    .X(_02834_));
 sky130_fd_sc_hd__mux4_1 _06888_ (.A0(\mem[60][2] ),
    .A1(\mem[61][2] ),
    .A2(\mem[62][2] ),
    .A3(\mem[63][2] ),
    .S0(_02487_),
    .S1(_02489_),
    .X(_02835_));
 sky130_fd_sc_hd__mux4_1 _06889_ (.A0(\mem[48][2] ),
    .A1(\mem[49][2] ),
    .A2(\mem[50][2] ),
    .A3(\mem[51][2] ),
    .S0(_02491_),
    .S1(_02492_),
    .X(_02836_));
 sky130_fd_sc_hd__clkbuf_4 _06890_ (.A(_02375_),
    .X(_02837_));
 sky130_fd_sc_hd__mux4_1 _06891_ (.A0(\mem[52][2] ),
    .A1(\mem[53][2] ),
    .A2(\mem[54][2] ),
    .A3(\mem[55][2] ),
    .S0(_02427_),
    .S1(_02837_),
    .X(_02838_));
 sky130_fd_sc_hd__mux4_1 _06892_ (.A0(\mem[56][2] ),
    .A1(\mem[57][2] ),
    .A2(\mem[58][2] ),
    .A3(\mem[59][2] ),
    .S0(_02502_),
    .S1(_02503_),
    .X(_02839_));
 sky130_fd_sc_hd__o22a_1 _06893_ (.A1(_02498_),
    .A2(_02838_),
    .B1(_02839_),
    .B2(_02506_),
    .X(_02840_));
 sky130_fd_sc_hd__o221a_1 _06894_ (.A1(_02485_),
    .A2(_02835_),
    .B1(_02836_),
    .B2(_02496_),
    .C1(_02840_),
    .X(_02841_));
 sky130_fd_sc_hd__o21a_1 _06895_ (.A1(_02482_),
    .A2(_02841_),
    .B1(_02510_),
    .X(_02842_));
 sky130_fd_sc_hd__a32o_1 _06896_ (.A1(_02356_),
    .A2(_02797_),
    .A3(_02824_),
    .B1(_02834_),
    .B2(_02842_),
    .X(_02843_));
 sky130_fd_sc_hd__o21a_1 _06897_ (.A1(\mem[93][2] ),
    .A2(_02515_),
    .B1(_02516_),
    .X(_02844_));
 sky130_fd_sc_hd__or3_1 _06898_ (.A(_02520_),
    .B(_02521_),
    .C(\mem[92][2] ),
    .X(_02845_));
 sky130_fd_sc_hd__o221a_1 _06899_ (.A1(\mem[94][2] ),
    .A2(_02518_),
    .B1(_02519_),
    .B2(\mem[95][2] ),
    .C1(_02845_),
    .X(_02846_));
 sky130_fd_sc_hd__o21a_1 _06900_ (.A1(\mem[80][2] ),
    .A2(_02524_),
    .B1(_02525_),
    .X(_02847_));
 sky130_fd_sc_hd__or3b_1 _06901_ (.A(_02529_),
    .B(\mem[82][2] ),
    .C_N(_02530_),
    .X(_02848_));
 sky130_fd_sc_hd__o221a_1 _06902_ (.A1(\mem[81][2] ),
    .A2(_02527_),
    .B1(_02528_),
    .B2(\mem[83][2] ),
    .C1(_02848_),
    .X(_02849_));
 sky130_fd_sc_hd__a22o_1 _06903_ (.A1(_02844_),
    .A2(_02846_),
    .B1(_02847_),
    .B2(_02849_),
    .X(_02850_));
 sky130_fd_sc_hd__o21a_1 _06904_ (.A1(\mem[88][2] ),
    .A2(_02535_),
    .B1(_02536_),
    .X(_02851_));
 sky130_fd_sc_hd__o22a_1 _06905_ (.A1(\mem[89][2] ),
    .A2(_02538_),
    .B1(_02539_),
    .B2(\mem[91][2] ),
    .X(_02852_));
 sky130_fd_sc_hd__o211a_1 _06906_ (.A1(\mem[90][2] ),
    .A2(_02534_),
    .B1(_02851_),
    .C1(_02852_),
    .X(_02853_));
 sky130_fd_sc_hd__or3_1 _06907_ (.A(_02545_),
    .B(_02546_),
    .C(\mem[84][2] ),
    .X(_02854_));
 sky130_fd_sc_hd__o221a_1 _06908_ (.A1(\mem[86][2] ),
    .A2(_02543_),
    .B1(_02544_),
    .B2(\mem[87][2] ),
    .C1(_02854_),
    .X(_02855_));
 sky130_fd_sc_hd__o211a_1 _06909_ (.A1(\mem[85][2] ),
    .A2(_02542_),
    .B1(_02855_),
    .C1(_02549_),
    .X(_02856_));
 sky130_fd_sc_hd__or4_4 _06910_ (.A(_02514_),
    .B(_02850_),
    .C(_02853_),
    .D(_02856_),
    .X(_02857_));
 sky130_fd_sc_hd__or3_1 _06911_ (.A(_02556_),
    .B(_02433_),
    .C(\mem[76][2] ),
    .X(_02858_));
 sky130_fd_sc_hd__o221a_1 _06912_ (.A1(\mem[78][2] ),
    .A2(_02554_),
    .B1(_02555_),
    .B2(\mem[79][2] ),
    .C1(_02858_),
    .X(_02859_));
 sky130_fd_sc_hd__o211a_1 _06913_ (.A1(\mem[77][2] ),
    .A2(_02553_),
    .B1(_02859_),
    .C1(_02559_),
    .X(_02860_));
 sky130_fd_sc_hd__o21a_1 _06914_ (.A1(\mem[64][2] ),
    .A2(_02562_),
    .B1(_02563_),
    .X(_02861_));
 sky130_fd_sc_hd__o22a_1 _06915_ (.A1(\mem[65][2] ),
    .A2(_02565_),
    .B1(_02566_),
    .B2(\mem[67][2] ),
    .X(_02862_));
 sky130_fd_sc_hd__o211a_1 _06916_ (.A1(\mem[66][2] ),
    .A2(_02561_),
    .B1(_02861_),
    .C1(_02862_),
    .X(_02863_));
 sky130_fd_sc_hd__or2_1 _06917_ (.A(\mem[72][2] ),
    .B(_02570_),
    .X(_02864_));
 sky130_fd_sc_hd__or3b_1 _06918_ (.A(_02574_),
    .B(\mem[74][2] ),
    .C_N(_02575_),
    .X(_02865_));
 sky130_fd_sc_hd__o221a_1 _06919_ (.A1(\mem[73][2] ),
    .A2(_02572_),
    .B1(_02573_),
    .B2(\mem[75][2] ),
    .C1(_02865_),
    .X(_02866_));
 sky130_fd_sc_hd__o21a_1 _06920_ (.A1(\mem[69][2] ),
    .A2(_02578_),
    .B1(_02579_),
    .X(_02867_));
 sky130_fd_sc_hd__buf_2 _06921_ (.A(_02388_),
    .X(_02868_));
 sky130_fd_sc_hd__or3_1 _06922_ (.A(_02583_),
    .B(_02868_),
    .C(\mem[68][2] ),
    .X(_02869_));
 sky130_fd_sc_hd__o221a_1 _06923_ (.A1(\mem[70][2] ),
    .A2(_02581_),
    .B1(_02582_),
    .B2(\mem[71][2] ),
    .C1(_02869_),
    .X(_02870_));
 sky130_fd_sc_hd__a32o_2 _06924_ (.A1(_02569_),
    .A2(_02864_),
    .A3(_02866_),
    .B1(_02867_),
    .B2(_02870_),
    .X(_02871_));
 sky130_fd_sc_hd__or4_4 _06925_ (.A(_02552_),
    .B(_02860_),
    .C(_02863_),
    .D(_02871_),
    .X(_02872_));
 sky130_fd_sc_hd__mux4_1 _06926_ (.A0(\mem[96][2] ),
    .A1(\mem[97][2] ),
    .A2(\mem[98][2] ),
    .A3(\mem[99][2] ),
    .S0(_02590_),
    .S1(_02591_),
    .X(_02873_));
 sky130_fd_sc_hd__mux4_1 _06927_ (.A0(\mem[100][2] ),
    .A1(\mem[101][2] ),
    .A2(\mem[102][2] ),
    .A3(\mem[103][2] ),
    .S0(_02593_),
    .S1(_02594_),
    .X(_02874_));
 sky130_fd_sc_hd__a22o_1 _06928_ (.A1(_02456_),
    .A2(_02873_),
    .B1(_02874_),
    .B2(_02465_),
    .X(_02875_));
 sky130_fd_sc_hd__mux4_2 _06929_ (.A0(\mem[108][2] ),
    .A1(\mem[109][2] ),
    .A2(\mem[110][2] ),
    .A3(\mem[111][2] ),
    .S0(_02600_),
    .S1(_02601_),
    .X(_02876_));
 sky130_fd_sc_hd__clkbuf_4 _06930_ (.A(_02459_),
    .X(_02877_));
 sky130_fd_sc_hd__mux4_1 _06931_ (.A0(\mem[104][2] ),
    .A1(\mem[105][2] ),
    .A2(\mem[106][2] ),
    .A3(\mem[107][2] ),
    .S0(_02604_),
    .S1(_02877_),
    .X(_02878_));
 sky130_fd_sc_hd__or2_1 _06932_ (.A(_02603_),
    .B(_02878_),
    .X(_02879_));
 sky130_fd_sc_hd__o211a_1 _06933_ (.A1(_02599_),
    .A2(_02876_),
    .B1(_02879_),
    .C1(_02608_),
    .X(_02880_));
 sky130_fd_sc_hd__or3_2 _06934_ (.A(_02589_),
    .B(_02875_),
    .C(_02880_),
    .X(_02881_));
 sky130_fd_sc_hd__mux4_1 _06935_ (.A0(\mem[124][2] ),
    .A1(\mem[125][2] ),
    .A2(\mem[126][2] ),
    .A3(\mem[127][2] ),
    .S0(_02613_),
    .S1(_02614_),
    .X(_02882_));
 sky130_fd_sc_hd__mux4_1 _06936_ (.A0(\mem[112][2] ),
    .A1(\mem[113][2] ),
    .A2(\mem[114][2] ),
    .A3(\mem[115][2] ),
    .S0(_02616_),
    .S1(_02618_),
    .X(_02883_));
 sky130_fd_sc_hd__buf_4 _06937_ (.A(_02495_),
    .X(_02884_));
 sky130_fd_sc_hd__buf_4 _06938_ (.A(_02497_),
    .X(_02885_));
 sky130_fd_sc_hd__mux4_1 _06939_ (.A0(\mem[116][2] ),
    .A1(\mem[117][2] ),
    .A2(\mem[118][2] ),
    .A3(\mem[119][2] ),
    .S0(_02622_),
    .S1(_02623_),
    .X(_02886_));
 sky130_fd_sc_hd__buf_6 _06940_ (.A(_02410_),
    .X(_02887_));
 sky130_fd_sc_hd__mux4_1 _06941_ (.A0(\mem[120][2] ),
    .A1(\mem[121][2] ),
    .A2(\mem[122][2] ),
    .A3(\mem[123][2] ),
    .S0(_02887_),
    .S1(_02626_),
    .X(_02888_));
 sky130_fd_sc_hd__buf_4 _06942_ (.A(_02505_),
    .X(_02889_));
 sky130_fd_sc_hd__o22a_1 _06943_ (.A1(_02885_),
    .A2(_02886_),
    .B1(_02888_),
    .B2(_02889_),
    .X(_02890_));
 sky130_fd_sc_hd__o221a_1 _06944_ (.A1(_02612_),
    .A2(_02882_),
    .B1(_02883_),
    .B2(_02884_),
    .C1(_02890_),
    .X(_02891_));
 sky130_fd_sc_hd__o21a_1 _06945_ (.A1(_02611_),
    .A2(_02891_),
    .B1(_02631_),
    .X(_02892_));
 sky130_fd_sc_hd__a32o_1 _06946_ (.A1(_02513_),
    .A2(_02857_),
    .A3(_02872_),
    .B1(_02881_),
    .B2(_02892_),
    .X(_02893_));
 sky130_fd_sc_hd__mux2_1 _06947_ (.A0(_02843_),
    .A1(_02893_),
    .S(_02635_),
    .X(_02894_));
 sky130_fd_sc_hd__clkbuf_1 _06948_ (.A(_02894_),
    .X(_00008_));
 sky130_fd_sc_hd__o21a_1 _06949_ (.A1(\mem[29][3] ),
    .A2(_02363_),
    .B1(_02366_),
    .X(_02895_));
 sky130_fd_sc_hd__or3_1 _06950_ (.A(_02374_),
    .B(_02779_),
    .C(\mem[28][3] ),
    .X(_02896_));
 sky130_fd_sc_hd__o221a_1 _06951_ (.A1(\mem[30][3] ),
    .A2(_02370_),
    .B1(_02372_),
    .B2(\mem[31][3] ),
    .C1(_02896_),
    .X(_02897_));
 sky130_fd_sc_hd__o21a_1 _06952_ (.A1(\mem[16][3] ),
    .A2(_02380_),
    .B1(_02383_),
    .X(_02898_));
 sky130_fd_sc_hd__clkbuf_4 _06953_ (.A(_02362_),
    .X(_02899_));
 sky130_fd_sc_hd__or3b_1 _06954_ (.A(_02387_),
    .B(\mem[18][3] ),
    .C_N(_02783_),
    .X(_02900_));
 sky130_fd_sc_hd__o221a_1 _06955_ (.A1(\mem[17][3] ),
    .A2(_02899_),
    .B1(_02386_),
    .B2(\mem[19][3] ),
    .C1(_02900_),
    .X(_02901_));
 sky130_fd_sc_hd__a22o_1 _06956_ (.A1(_02895_),
    .A2(_02897_),
    .B1(_02898_),
    .B2(_02901_),
    .X(_02902_));
 sky130_fd_sc_hd__o21a_1 _06957_ (.A1(\mem[24][3] ),
    .A2(_02788_),
    .B1(_02397_),
    .X(_02903_));
 sky130_fd_sc_hd__o22a_1 _06958_ (.A1(\mem[25][3] ),
    .A2(_02790_),
    .B1(_02401_),
    .B2(\mem[27][3] ),
    .X(_02904_));
 sky130_fd_sc_hd__o211a_1 _06959_ (.A1(\mem[26][3] ),
    .A2(_02787_),
    .B1(_02903_),
    .C1(_02904_),
    .X(_02905_));
 sky130_fd_sc_hd__or3_1 _06960_ (.A(_02793_),
    .B(_02412_),
    .C(\mem[20][3] ),
    .X(_02906_));
 sky130_fd_sc_hd__o221a_1 _06961_ (.A1(\mem[22][3] ),
    .A2(_02407_),
    .B1(_02409_),
    .B2(\mem[23][3] ),
    .C1(_02906_),
    .X(_02907_));
 sky130_fd_sc_hd__o211a_1 _06962_ (.A1(\mem[21][3] ),
    .A2(_02406_),
    .B1(_02907_),
    .C1(_02417_),
    .X(_02908_));
 sky130_fd_sc_hd__or4_2 _06963_ (.A(_02358_),
    .B(_02902_),
    .C(_02905_),
    .D(_02908_),
    .X(_02909_));
 sky130_fd_sc_hd__or3_1 _06964_ (.A(_02802_),
    .B(_02803_),
    .C(\mem[12][3] ),
    .X(_02910_));
 sky130_fd_sc_hd__o221a_1 _06965_ (.A1(\mem[14][3] ),
    .A2(_02800_),
    .B1(_02801_),
    .B2(\mem[15][3] ),
    .C1(_02910_),
    .X(_02911_));
 sky130_fd_sc_hd__o211a_1 _06966_ (.A1(\mem[13][3] ),
    .A2(_02799_),
    .B1(_02911_),
    .C1(_02806_),
    .X(_02912_));
 sky130_fd_sc_hd__o21a_1 _06967_ (.A1(\mem[0][3] ),
    .A2(_02438_),
    .B1(_02455_),
    .X(_02913_));
 sky130_fd_sc_hd__clkbuf_4 _06968_ (.A(_02400_),
    .X(_02914_));
 sky130_fd_sc_hd__o22a_1 _06969_ (.A1(\mem[1][3] ),
    .A2(_02441_),
    .B1(_02914_),
    .B2(\mem[3][3] ),
    .X(_02915_));
 sky130_fd_sc_hd__o211a_1 _06970_ (.A1(\mem[2][3] ),
    .A2(_02437_),
    .B1(_02913_),
    .C1(_02915_),
    .X(_02916_));
 sky130_fd_sc_hd__clkbuf_2 _06971_ (.A(_02378_),
    .X(_02917_));
 sky130_fd_sc_hd__or2_1 _06972_ (.A(\mem[8][3] ),
    .B(_02917_),
    .X(_02918_));
 sky130_fd_sc_hd__or3b_1 _06973_ (.A(_02815_),
    .B(\mem[10][3] ),
    .C_N(_02816_),
    .X(_02919_));
 sky130_fd_sc_hd__o221a_1 _06974_ (.A1(\mem[9][3] ),
    .A2(_02736_),
    .B1(_02814_),
    .B2(\mem[11][3] ),
    .C1(_02919_),
    .X(_02920_));
 sky130_fd_sc_hd__o21a_1 _06975_ (.A1(\mem[5][3] ),
    .A2(_02819_),
    .B1(_02416_),
    .X(_02921_));
 sky130_fd_sc_hd__or3_1 _06976_ (.A(_02447_),
    .B(_02429_),
    .C(\mem[4][3] ),
    .X(_02922_));
 sky130_fd_sc_hd__o221a_2 _06977_ (.A1(\mem[6][3] ),
    .A2(_02445_),
    .B1(_02446_),
    .B2(\mem[7][3] ),
    .C1(_02922_),
    .X(_02923_));
 sky130_fd_sc_hd__a32o_1 _06978_ (.A1(_02811_),
    .A2(_02918_),
    .A3(_02920_),
    .B1(_02921_),
    .B2(_02923_),
    .X(_02924_));
 sky130_fd_sc_hd__or4_1 _06979_ (.A(_02798_),
    .B(_02912_),
    .C(_02916_),
    .D(_02924_),
    .X(_02925_));
 sky130_fd_sc_hd__buf_4 _06980_ (.A(_02460_),
    .X(_02926_));
 sky130_fd_sc_hd__mux4_1 _06981_ (.A0(\mem[36][3] ),
    .A1(\mem[37][3] ),
    .A2(\mem[38][3] ),
    .A3(\mem[39][3] ),
    .S0(_02826_),
    .S1(_02926_),
    .X(_02927_));
 sky130_fd_sc_hd__buf_6 _06982_ (.A(_02374_),
    .X(_02928_));
 sky130_fd_sc_hd__buf_4 _06983_ (.A(_02488_),
    .X(_02929_));
 sky130_fd_sc_hd__mux4_1 _06984_ (.A0(\mem[32][3] ),
    .A1(\mem[33][3] ),
    .A2(\mem[34][3] ),
    .A3(\mem[35][3] ),
    .S0(_02928_),
    .S1(_02929_),
    .X(_02930_));
 sky130_fd_sc_hd__a22o_1 _06985_ (.A1(_02825_),
    .A2(_02927_),
    .B1(_02930_),
    .B2(_02596_),
    .X(_02931_));
 sky130_fd_sc_hd__mux4_1 _06986_ (.A0(\mem[44][3] ),
    .A1(\mem[45][3] ),
    .A2(\mem[46][3] ),
    .A3(\mem[47][3] ),
    .S0(_02467_),
    .S1(_02468_),
    .X(_02932_));
 sky130_fd_sc_hd__mux4_1 _06987_ (.A0(\mem[40][3] ),
    .A1(\mem[41][3] ),
    .A2(\mem[42][3] ),
    .A3(\mem[43][3] ),
    .S0(_02457_),
    .S1(_02460_),
    .X(_02933_));
 sky130_fd_sc_hd__or2_1 _06988_ (.A(_02475_),
    .B(_02933_),
    .X(_02934_));
 sky130_fd_sc_hd__o211a_1 _06989_ (.A1(_02472_),
    .A2(_02932_),
    .B1(_02934_),
    .C1(_02479_),
    .X(_02935_));
 sky130_fd_sc_hd__or3_4 _06990_ (.A(_02453_),
    .B(_02931_),
    .C(_02935_),
    .X(_02936_));
 sky130_fd_sc_hd__mux4_1 _06991_ (.A0(\mem[60][3] ),
    .A1(\mem[61][3] ),
    .A2(\mem[62][3] ),
    .A3(\mem[63][3] ),
    .S0(_02487_),
    .S1(_02489_),
    .X(_02937_));
 sky130_fd_sc_hd__mux4_1 _06992_ (.A0(\mem[48][3] ),
    .A1(\mem[49][3] ),
    .A2(\mem[50][3] ),
    .A3(\mem[51][3] ),
    .S0(_02491_),
    .S1(_02492_),
    .X(_02938_));
 sky130_fd_sc_hd__mux4_1 _06993_ (.A0(\mem[52][3] ),
    .A1(\mem[53][3] ),
    .A2(\mem[54][3] ),
    .A3(\mem[55][3] ),
    .S0(_02427_),
    .S1(_02837_),
    .X(_02939_));
 sky130_fd_sc_hd__mux4_1 _06994_ (.A0(\mem[56][3] ),
    .A1(\mem[57][3] ),
    .A2(\mem[58][3] ),
    .A3(\mem[59][3] ),
    .S0(_02502_),
    .S1(_02503_),
    .X(_02940_));
 sky130_fd_sc_hd__o22a_1 _06995_ (.A1(_02498_),
    .A2(_02939_),
    .B1(_02940_),
    .B2(_02506_),
    .X(_02941_));
 sky130_fd_sc_hd__o221a_1 _06996_ (.A1(_02485_),
    .A2(_02937_),
    .B1(_02938_),
    .B2(_02496_),
    .C1(_02941_),
    .X(_02942_));
 sky130_fd_sc_hd__o21a_1 _06997_ (.A1(_02482_),
    .A2(_02942_),
    .B1(_02510_),
    .X(_02943_));
 sky130_fd_sc_hd__a32o_1 _06998_ (.A1(_02356_),
    .A2(_02909_),
    .A3(_02925_),
    .B1(_02936_),
    .B2(_02943_),
    .X(_02944_));
 sky130_fd_sc_hd__o21a_1 _06999_ (.A1(\mem[93][3] ),
    .A2(_02515_),
    .B1(_02516_),
    .X(_02945_));
 sky130_fd_sc_hd__or3_1 _07000_ (.A(_02466_),
    .B(_02521_),
    .C(\mem[92][3] ),
    .X(_02946_));
 sky130_fd_sc_hd__o221a_1 _07001_ (.A1(\mem[94][3] ),
    .A2(_02518_),
    .B1(_02519_),
    .B2(\mem[95][3] ),
    .C1(_02946_),
    .X(_02947_));
 sky130_fd_sc_hd__o21a_1 _07002_ (.A1(\mem[80][3] ),
    .A2(_02524_),
    .B1(_02525_),
    .X(_02948_));
 sky130_fd_sc_hd__or3b_1 _07003_ (.A(_02529_),
    .B(\mem[82][3] ),
    .C_N(_02530_),
    .X(_02949_));
 sky130_fd_sc_hd__o221a_1 _07004_ (.A1(\mem[81][3] ),
    .A2(_02527_),
    .B1(_02424_),
    .B2(\mem[83][3] ),
    .C1(_02949_),
    .X(_02950_));
 sky130_fd_sc_hd__a22o_1 _07005_ (.A1(_02945_),
    .A2(_02947_),
    .B1(_02948_),
    .B2(_02950_),
    .X(_02951_));
 sky130_fd_sc_hd__o21a_1 _07006_ (.A1(\mem[88][3] ),
    .A2(_02535_),
    .B1(_02536_),
    .X(_02952_));
 sky130_fd_sc_hd__o22a_1 _07007_ (.A1(\mem[89][3] ),
    .A2(_02538_),
    .B1(_02539_),
    .B2(\mem[91][3] ),
    .X(_02953_));
 sky130_fd_sc_hd__o211a_1 _07008_ (.A1(\mem[90][3] ),
    .A2(_02534_),
    .B1(_02952_),
    .C1(_02953_),
    .X(_02954_));
 sky130_fd_sc_hd__buf_4 _07009_ (.A(_02441_),
    .X(_02955_));
 sky130_fd_sc_hd__buf_4 _07010_ (.A(_02369_),
    .X(_02956_));
 sky130_fd_sc_hd__or3_1 _07011_ (.A(_02545_),
    .B(_02546_),
    .C(\mem[84][3] ),
    .X(_02957_));
 sky130_fd_sc_hd__o221a_1 _07012_ (.A1(\mem[86][3] ),
    .A2(_02956_),
    .B1(_02544_),
    .B2(\mem[87][3] ),
    .C1(_02957_),
    .X(_02958_));
 sky130_fd_sc_hd__o211a_1 _07013_ (.A1(\mem[85][3] ),
    .A2(_02955_),
    .B1(_02958_),
    .C1(_02549_),
    .X(_02959_));
 sky130_fd_sc_hd__or4_4 _07014_ (.A(_02514_),
    .B(_02951_),
    .C(_02954_),
    .D(_02959_),
    .X(_02960_));
 sky130_fd_sc_hd__or3_1 _07015_ (.A(_02556_),
    .B(_02433_),
    .C(\mem[76][3] ),
    .X(_02961_));
 sky130_fd_sc_hd__o221a_1 _07016_ (.A1(\mem[78][3] ),
    .A2(_02554_),
    .B1(_02555_),
    .B2(\mem[79][3] ),
    .C1(_02961_),
    .X(_02962_));
 sky130_fd_sc_hd__o211a_1 _07017_ (.A1(\mem[77][3] ),
    .A2(_02553_),
    .B1(_02962_),
    .C1(_02559_),
    .X(_02963_));
 sky130_fd_sc_hd__o21a_1 _07018_ (.A1(\mem[64][3] ),
    .A2(_02395_),
    .B1(_02563_),
    .X(_02964_));
 sky130_fd_sc_hd__o22a_1 _07019_ (.A1(\mem[65][3] ),
    .A2(_02565_),
    .B1(_02566_),
    .B2(\mem[67][3] ),
    .X(_02965_));
 sky130_fd_sc_hd__o211a_1 _07020_ (.A1(\mem[66][3] ),
    .A2(_02394_),
    .B1(_02964_),
    .C1(_02965_),
    .X(_02966_));
 sky130_fd_sc_hd__or2_1 _07021_ (.A(\mem[72][3] ),
    .B(_02570_),
    .X(_02967_));
 sky130_fd_sc_hd__or3b_1 _07022_ (.A(_02574_),
    .B(\mem[74][3] ),
    .C_N(_02575_),
    .X(_02968_));
 sky130_fd_sc_hd__o221a_1 _07023_ (.A1(\mem[73][3] ),
    .A2(_02572_),
    .B1(_02573_),
    .B2(\mem[75][3] ),
    .C1(_02968_),
    .X(_02969_));
 sky130_fd_sc_hd__o21a_1 _07024_ (.A1(\mem[69][3] ),
    .A2(_02578_),
    .B1(_02463_),
    .X(_02970_));
 sky130_fd_sc_hd__or3_1 _07025_ (.A(_02583_),
    .B(_02868_),
    .C(\mem[68][3] ),
    .X(_02971_));
 sky130_fd_sc_hd__o221a_1 _07026_ (.A1(\mem[70][3] ),
    .A2(_02581_),
    .B1(_02582_),
    .B2(\mem[71][3] ),
    .C1(_02971_),
    .X(_02972_));
 sky130_fd_sc_hd__a32o_1 _07027_ (.A1(_02569_),
    .A2(_02967_),
    .A3(_02969_),
    .B1(_02970_),
    .B2(_02972_),
    .X(_02973_));
 sky130_fd_sc_hd__or4_4 _07028_ (.A(_02552_),
    .B(_02963_),
    .C(_02966_),
    .D(_02973_),
    .X(_02974_));
 sky130_fd_sc_hd__mux4_1 _07029_ (.A0(\mem[96][3] ),
    .A1(\mem[97][3] ),
    .A2(\mem[98][3] ),
    .A3(\mem[99][3] ),
    .S0(_02590_),
    .S1(_02591_),
    .X(_02975_));
 sky130_fd_sc_hd__mux4_1 _07030_ (.A0(\mem[100][3] ),
    .A1(\mem[101][3] ),
    .A2(\mem[102][3] ),
    .A3(\mem[103][3] ),
    .S0(_02593_),
    .S1(_02594_),
    .X(_02976_));
 sky130_fd_sc_hd__a22o_1 _07031_ (.A1(_02456_),
    .A2(_02975_),
    .B1(_02976_),
    .B2(_02825_),
    .X(_02977_));
 sky130_fd_sc_hd__mux4_2 _07032_ (.A0(\mem[108][3] ),
    .A1(\mem[109][3] ),
    .A2(\mem[110][3] ),
    .A3(\mem[111][3] ),
    .S0(_02458_),
    .S1(_02601_),
    .X(_02978_));
 sky130_fd_sc_hd__mux4_1 _07033_ (.A0(\mem[104][3] ),
    .A1(\mem[105][3] ),
    .A2(\mem[106][3] ),
    .A3(\mem[107][3] ),
    .S0(_02604_),
    .S1(_02877_),
    .X(_02979_));
 sky130_fd_sc_hd__or2_1 _07034_ (.A(_02474_),
    .B(_02979_),
    .X(_02980_));
 sky130_fd_sc_hd__o211a_1 _07035_ (.A1(_02599_),
    .A2(_02978_),
    .B1(_02980_),
    .C1(_02608_),
    .X(_02981_));
 sky130_fd_sc_hd__or3_1 _07036_ (.A(_02589_),
    .B(_02977_),
    .C(_02981_),
    .X(_02982_));
 sky130_fd_sc_hd__mux4_1 _07037_ (.A0(\mem[124][3] ),
    .A1(\mem[125][3] ),
    .A2(\mem[126][3] ),
    .A3(\mem[127][3] ),
    .S0(_02613_),
    .S1(_02614_),
    .X(_02983_));
 sky130_fd_sc_hd__mux4_1 _07038_ (.A0(\mem[112][3] ),
    .A1(\mem[113][3] ),
    .A2(\mem[114][3] ),
    .A3(\mem[115][3] ),
    .S0(_02616_),
    .S1(_02618_),
    .X(_02984_));
 sky130_fd_sc_hd__buf_6 _07039_ (.A(_02410_),
    .X(_02985_));
 sky130_fd_sc_hd__mux4_1 _07040_ (.A0(\mem[116][3] ),
    .A1(\mem[117][3] ),
    .A2(\mem[118][3] ),
    .A3(\mem[119][3] ),
    .S0(_02985_),
    .S1(_02623_),
    .X(_02986_));
 sky130_fd_sc_hd__mux4_1 _07041_ (.A0(\mem[120][3] ),
    .A1(\mem[121][3] ),
    .A2(\mem[122][3] ),
    .A3(\mem[123][3] ),
    .S0(_02887_),
    .S1(_02626_),
    .X(_02987_));
 sky130_fd_sc_hd__o22a_1 _07042_ (.A1(_02885_),
    .A2(_02986_),
    .B1(_02987_),
    .B2(_02889_),
    .X(_02988_));
 sky130_fd_sc_hd__o221a_1 _07043_ (.A1(_02612_),
    .A2(_02983_),
    .B1(_02984_),
    .B2(_02884_),
    .C1(_02988_),
    .X(_02989_));
 sky130_fd_sc_hd__o21a_1 _07044_ (.A1(_02611_),
    .A2(_02989_),
    .B1(_02631_),
    .X(_02990_));
 sky130_fd_sc_hd__a32o_1 _07045_ (.A1(_02513_),
    .A2(_02960_),
    .A3(_02974_),
    .B1(_02982_),
    .B2(_02990_),
    .X(_02991_));
 sky130_fd_sc_hd__mux2_1 _07046_ (.A0(_02944_),
    .A1(_02991_),
    .S(_02635_),
    .X(_02992_));
 sky130_fd_sc_hd__clkbuf_1 _07047_ (.A(_02992_),
    .X(_00009_));
 sky130_fd_sc_hd__clkbuf_4 _07048_ (.A(_02357_),
    .X(_02993_));
 sky130_fd_sc_hd__o21a_1 _07049_ (.A1(\mem[29][4] ),
    .A2(_02363_),
    .B1(_02366_),
    .X(_02994_));
 sky130_fd_sc_hd__clkbuf_4 _07050_ (.A(_02368_),
    .X(_02995_));
 sky130_fd_sc_hd__or3_1 _07051_ (.A(_02374_),
    .B(_02779_),
    .C(\mem[28][4] ),
    .X(_02996_));
 sky130_fd_sc_hd__o221a_1 _07052_ (.A1(\mem[30][4] ),
    .A2(_02995_),
    .B1(_02372_),
    .B2(\mem[31][4] ),
    .C1(_02996_),
    .X(_02997_));
 sky130_fd_sc_hd__o21a_1 _07053_ (.A1(\mem[16][4] ),
    .A2(_02380_),
    .B1(_02383_),
    .X(_02998_));
 sky130_fd_sc_hd__or3b_1 _07054_ (.A(_02387_),
    .B(\mem[18][4] ),
    .C_N(_02783_),
    .X(_02999_));
 sky130_fd_sc_hd__o221a_1 _07055_ (.A1(\mem[17][4] ),
    .A2(_02899_),
    .B1(_02386_),
    .B2(\mem[19][4] ),
    .C1(_02999_),
    .X(_03000_));
 sky130_fd_sc_hd__a22o_1 _07056_ (.A1(_02994_),
    .A2(_02997_),
    .B1(_02998_),
    .B2(_03000_),
    .X(_03001_));
 sky130_fd_sc_hd__o21a_1 _07057_ (.A1(\mem[24][4] ),
    .A2(_02788_),
    .B1(_02397_),
    .X(_03002_));
 sky130_fd_sc_hd__o22a_1 _07058_ (.A1(\mem[25][4] ),
    .A2(_02790_),
    .B1(_02401_),
    .B2(\mem[27][4] ),
    .X(_03003_));
 sky130_fd_sc_hd__o211a_1 _07059_ (.A1(\mem[26][4] ),
    .A2(_02787_),
    .B1(_03002_),
    .C1(_03003_),
    .X(_03004_));
 sky130_fd_sc_hd__or3_1 _07060_ (.A(_02793_),
    .B(_02412_),
    .C(\mem[20][4] ),
    .X(_03005_));
 sky130_fd_sc_hd__o221a_1 _07061_ (.A1(\mem[22][4] ),
    .A2(_02407_),
    .B1(_02409_),
    .B2(\mem[23][4] ),
    .C1(_03005_),
    .X(_03006_));
 sky130_fd_sc_hd__o211a_1 _07062_ (.A1(\mem[21][4] ),
    .A2(_02406_),
    .B1(_03006_),
    .C1(_02417_),
    .X(_03007_));
 sky130_fd_sc_hd__or4_2 _07063_ (.A(_02993_),
    .B(_03001_),
    .C(_03004_),
    .D(_03007_),
    .X(_03008_));
 sky130_fd_sc_hd__buf_4 _07064_ (.A(_02408_),
    .X(_03009_));
 sky130_fd_sc_hd__or3_1 _07065_ (.A(_02802_),
    .B(_02803_),
    .C(\mem[12][4] ),
    .X(_03010_));
 sky130_fd_sc_hd__o221a_1 _07066_ (.A1(\mem[14][4] ),
    .A2(_02800_),
    .B1(_03009_),
    .B2(\mem[15][4] ),
    .C1(_03010_),
    .X(_03011_));
 sky130_fd_sc_hd__o211a_1 _07067_ (.A1(\mem[13][4] ),
    .A2(_02799_),
    .B1(_03011_),
    .C1(_02806_),
    .X(_03012_));
 sky130_fd_sc_hd__clkbuf_4 _07068_ (.A(_02454_),
    .X(_03013_));
 sky130_fd_sc_hd__o21a_1 _07069_ (.A1(\mem[0][4] ),
    .A2(_02438_),
    .B1(_03013_),
    .X(_03014_));
 sky130_fd_sc_hd__o22a_1 _07070_ (.A1(\mem[1][4] ),
    .A2(_02441_),
    .B1(_02914_),
    .B2(\mem[3][4] ),
    .X(_03015_));
 sky130_fd_sc_hd__o211a_1 _07071_ (.A1(\mem[2][4] ),
    .A2(_02437_),
    .B1(_03014_),
    .C1(_03015_),
    .X(_03016_));
 sky130_fd_sc_hd__or2_1 _07072_ (.A(\mem[8][4] ),
    .B(_02917_),
    .X(_03017_));
 sky130_fd_sc_hd__or3b_1 _07073_ (.A(_02815_),
    .B(\mem[10][4] ),
    .C_N(_02816_),
    .X(_03018_));
 sky130_fd_sc_hd__o221a_1 _07074_ (.A1(\mem[9][4] ),
    .A2(_02736_),
    .B1(_02814_),
    .B2(\mem[11][4] ),
    .C1(_03018_),
    .X(_03019_));
 sky130_fd_sc_hd__o21a_1 _07075_ (.A1(\mem[5][4] ),
    .A2(_02819_),
    .B1(_02416_),
    .X(_03020_));
 sky130_fd_sc_hd__or3_1 _07076_ (.A(_02447_),
    .B(_02429_),
    .C(\mem[4][4] ),
    .X(_03021_));
 sky130_fd_sc_hd__o221a_2 _07077_ (.A1(\mem[6][4] ),
    .A2(_02445_),
    .B1(_02446_),
    .B2(\mem[7][4] ),
    .C1(_03021_),
    .X(_03022_));
 sky130_fd_sc_hd__a32o_1 _07078_ (.A1(_02811_),
    .A2(_03017_),
    .A3(_03019_),
    .B1(_03020_),
    .B2(_03022_),
    .X(_03023_));
 sky130_fd_sc_hd__or4_1 _07079_ (.A(_02798_),
    .B(_03012_),
    .C(_03016_),
    .D(_03023_),
    .X(_03024_));
 sky130_fd_sc_hd__mux4_1 _07080_ (.A0(\mem[36][4] ),
    .A1(\mem[37][4] ),
    .A2(\mem[38][4] ),
    .A3(\mem[39][4] ),
    .S0(_02826_),
    .S1(_02926_),
    .X(_03025_));
 sky130_fd_sc_hd__mux4_1 _07081_ (.A0(\mem[32][4] ),
    .A1(\mem[33][4] ),
    .A2(\mem[34][4] ),
    .A3(\mem[35][4] ),
    .S0(_02928_),
    .S1(_02929_),
    .X(_03026_));
 sky130_fd_sc_hd__a22o_1 _07082_ (.A1(_02825_),
    .A2(_03025_),
    .B1(_03026_),
    .B2(_02596_),
    .X(_03027_));
 sky130_fd_sc_hd__mux4_1 _07083_ (.A0(\mem[44][4] ),
    .A1(\mem[45][4] ),
    .A2(\mem[46][4] ),
    .A3(\mem[47][4] ),
    .S0(_02467_),
    .S1(_02468_),
    .X(_03028_));
 sky130_fd_sc_hd__mux4_1 _07084_ (.A0(\mem[40][4] ),
    .A1(\mem[41][4] ),
    .A2(\mem[42][4] ),
    .A3(\mem[43][4] ),
    .S0(_02457_),
    .S1(_02460_),
    .X(_03029_));
 sky130_fd_sc_hd__or2_1 _07085_ (.A(_02475_),
    .B(_03029_),
    .X(_03030_));
 sky130_fd_sc_hd__o211a_1 _07086_ (.A1(_02472_),
    .A2(_03028_),
    .B1(_03030_),
    .C1(_02479_),
    .X(_03031_));
 sky130_fd_sc_hd__or3_4 _07087_ (.A(_02453_),
    .B(_03027_),
    .C(_03031_),
    .X(_03032_));
 sky130_fd_sc_hd__clkbuf_4 _07088_ (.A(_02484_),
    .X(_03033_));
 sky130_fd_sc_hd__mux4_1 _07089_ (.A0(\mem[60][4] ),
    .A1(\mem[61][4] ),
    .A2(\mem[62][4] ),
    .A3(\mem[63][4] ),
    .S0(_02487_),
    .S1(_02489_),
    .X(_03034_));
 sky130_fd_sc_hd__mux4_1 _07090_ (.A0(\mem[48][4] ),
    .A1(\mem[49][4] ),
    .A2(\mem[50][4] ),
    .A3(\mem[51][4] ),
    .S0(_02491_),
    .S1(_02492_),
    .X(_03035_));
 sky130_fd_sc_hd__mux4_1 _07091_ (.A0(\mem[52][4] ),
    .A1(\mem[53][4] ),
    .A2(\mem[54][4] ),
    .A3(\mem[55][4] ),
    .S0(_02427_),
    .S1(_02837_),
    .X(_03036_));
 sky130_fd_sc_hd__mux4_1 _07092_ (.A0(\mem[56][4] ),
    .A1(\mem[57][4] ),
    .A2(\mem[58][4] ),
    .A3(\mem[59][4] ),
    .S0(_02502_),
    .S1(_02503_),
    .X(_03037_));
 sky130_fd_sc_hd__o22a_1 _07093_ (.A1(_02498_),
    .A2(_03036_),
    .B1(_03037_),
    .B2(_02506_),
    .X(_03038_));
 sky130_fd_sc_hd__o221a_1 _07094_ (.A1(_03033_),
    .A2(_03034_),
    .B1(_03035_),
    .B2(_02496_),
    .C1(_03038_),
    .X(_03039_));
 sky130_fd_sc_hd__o21a_1 _07095_ (.A1(_02482_),
    .A2(_03039_),
    .B1(_02510_),
    .X(_03040_));
 sky130_fd_sc_hd__a32o_1 _07096_ (.A1(_02356_),
    .A2(_03008_),
    .A3(_03024_),
    .B1(_03032_),
    .B2(_03040_),
    .X(_03041_));
 sky130_fd_sc_hd__clkbuf_8 _07097_ (.A(_02362_),
    .X(_03042_));
 sky130_fd_sc_hd__o21a_1 _07098_ (.A1(\mem[93][4] ),
    .A2(_03042_),
    .B1(_02516_),
    .X(_03043_));
 sky130_fd_sc_hd__or3_1 _07099_ (.A(_02466_),
    .B(_02521_),
    .C(\mem[92][4] ),
    .X(_03044_));
 sky130_fd_sc_hd__o221a_1 _07100_ (.A1(\mem[94][4] ),
    .A2(_02518_),
    .B1(_02519_),
    .B2(\mem[95][4] ),
    .C1(_03044_),
    .X(_03045_));
 sky130_fd_sc_hd__o21a_1 _07101_ (.A1(\mem[80][4] ),
    .A2(_02524_),
    .B1(_02525_),
    .X(_03046_));
 sky130_fd_sc_hd__or3b_1 _07102_ (.A(_02529_),
    .B(\mem[82][4] ),
    .C_N(_02530_),
    .X(_03047_));
 sky130_fd_sc_hd__o221a_1 _07103_ (.A1(\mem[81][4] ),
    .A2(_02527_),
    .B1(_02424_),
    .B2(\mem[83][4] ),
    .C1(_03047_),
    .X(_03048_));
 sky130_fd_sc_hd__a22o_1 _07104_ (.A1(_03043_),
    .A2(_03045_),
    .B1(_03046_),
    .B2(_03048_),
    .X(_03049_));
 sky130_fd_sc_hd__o21a_1 _07105_ (.A1(\mem[88][4] ),
    .A2(_02535_),
    .B1(_02536_),
    .X(_03050_));
 sky130_fd_sc_hd__o22a_1 _07106_ (.A1(\mem[89][4] ),
    .A2(_02538_),
    .B1(_02539_),
    .B2(\mem[91][4] ),
    .X(_03051_));
 sky130_fd_sc_hd__o211a_1 _07107_ (.A1(\mem[90][4] ),
    .A2(_02534_),
    .B1(_03050_),
    .C1(_03051_),
    .X(_03052_));
 sky130_fd_sc_hd__or3_1 _07108_ (.A(_02545_),
    .B(_02546_),
    .C(\mem[84][4] ),
    .X(_03053_));
 sky130_fd_sc_hd__o221a_1 _07109_ (.A1(\mem[86][4] ),
    .A2(_02956_),
    .B1(_02664_),
    .B2(\mem[87][4] ),
    .C1(_03053_),
    .X(_03054_));
 sky130_fd_sc_hd__o211a_1 _07110_ (.A1(\mem[85][4] ),
    .A2(_02955_),
    .B1(_03054_),
    .C1(_02549_),
    .X(_03055_));
 sky130_fd_sc_hd__or4_4 _07111_ (.A(_02514_),
    .B(_03049_),
    .C(_03052_),
    .D(_03055_),
    .X(_03056_));
 sky130_fd_sc_hd__or3_1 _07112_ (.A(_02556_),
    .B(_02433_),
    .C(\mem[76][4] ),
    .X(_03057_));
 sky130_fd_sc_hd__o221a_1 _07113_ (.A1(\mem[78][4] ),
    .A2(_02554_),
    .B1(_02555_),
    .B2(\mem[79][4] ),
    .C1(_03057_),
    .X(_03058_));
 sky130_fd_sc_hd__o211a_1 _07114_ (.A1(\mem[77][4] ),
    .A2(_02553_),
    .B1(_03058_),
    .C1(_02559_),
    .X(_03059_));
 sky130_fd_sc_hd__o21a_1 _07115_ (.A1(\mem[64][4] ),
    .A2(_02395_),
    .B1(_02563_),
    .X(_03060_));
 sky130_fd_sc_hd__o22a_1 _07116_ (.A1(\mem[65][4] ),
    .A2(_02399_),
    .B1(_02566_),
    .B2(\mem[67][4] ),
    .X(_03061_));
 sky130_fd_sc_hd__o211a_1 _07117_ (.A1(\mem[66][4] ),
    .A2(_02394_),
    .B1(_03060_),
    .C1(_03061_),
    .X(_03062_));
 sky130_fd_sc_hd__or2_1 _07118_ (.A(\mem[72][4] ),
    .B(_02570_),
    .X(_03063_));
 sky130_fd_sc_hd__or3b_1 _07119_ (.A(_02574_),
    .B(\mem[74][4] ),
    .C_N(_02575_),
    .X(_03064_));
 sky130_fd_sc_hd__o221a_1 _07120_ (.A1(\mem[73][4] ),
    .A2(_02572_),
    .B1(_02801_),
    .B2(\mem[75][4] ),
    .C1(_03064_),
    .X(_03065_));
 sky130_fd_sc_hd__o21a_1 _07121_ (.A1(\mem[69][4] ),
    .A2(_02578_),
    .B1(_02463_),
    .X(_03066_));
 sky130_fd_sc_hd__or3_1 _07122_ (.A(_02583_),
    .B(_02868_),
    .C(\mem[68][4] ),
    .X(_03067_));
 sky130_fd_sc_hd__o221a_1 _07123_ (.A1(\mem[70][4] ),
    .A2(_02581_),
    .B1(_02582_),
    .B2(\mem[71][4] ),
    .C1(_03067_),
    .X(_03068_));
 sky130_fd_sc_hd__a32o_1 _07124_ (.A1(_02569_),
    .A2(_03063_),
    .A3(_03065_),
    .B1(_03066_),
    .B2(_03068_),
    .X(_03069_));
 sky130_fd_sc_hd__or4_4 _07125_ (.A(_02552_),
    .B(_03059_),
    .C(_03062_),
    .D(_03069_),
    .X(_03070_));
 sky130_fd_sc_hd__mux4_1 _07126_ (.A0(\mem[100][4] ),
    .A1(\mem[101][4] ),
    .A2(\mem[102][4] ),
    .A3(\mem[103][4] ),
    .S0(_02590_),
    .S1(_02591_),
    .X(_03071_));
 sky130_fd_sc_hd__mux4_1 _07127_ (.A0(\mem[96][4] ),
    .A1(\mem[97][4] ),
    .A2(\mem[98][4] ),
    .A3(\mem[99][4] ),
    .S0(_02593_),
    .S1(_02594_),
    .X(_03072_));
 sky130_fd_sc_hd__a22o_1 _07128_ (.A1(_02450_),
    .A2(_03071_),
    .B1(_03072_),
    .B2(_02596_),
    .X(_03073_));
 sky130_fd_sc_hd__mux4_1 _07129_ (.A0(\mem[108][4] ),
    .A1(\mem[109][4] ),
    .A2(\mem[110][4] ),
    .A3(\mem[111][4] ),
    .S0(_02458_),
    .S1(_02461_),
    .X(_03074_));
 sky130_fd_sc_hd__mux4_1 _07130_ (.A0(\mem[104][4] ),
    .A1(\mem[105][4] ),
    .A2(\mem[106][4] ),
    .A3(\mem[107][4] ),
    .S0(_02501_),
    .S1(_02877_),
    .X(_03075_));
 sky130_fd_sc_hd__or2_1 _07131_ (.A(_02474_),
    .B(_03075_),
    .X(_03076_));
 sky130_fd_sc_hd__o211a_1 _07132_ (.A1(_02599_),
    .A2(_03074_),
    .B1(_03076_),
    .C1(_02478_),
    .X(_03077_));
 sky130_fd_sc_hd__or3_1 _07133_ (.A(_02589_),
    .B(_03073_),
    .C(_03077_),
    .X(_03078_));
 sky130_fd_sc_hd__mux4_1 _07134_ (.A0(\mem[124][4] ),
    .A1(\mem[125][4] ),
    .A2(\mem[126][4] ),
    .A3(\mem[127][4] ),
    .S0(_02613_),
    .S1(_02703_),
    .X(_03079_));
 sky130_fd_sc_hd__mux4_1 _07135_ (.A0(\mem[112][4] ),
    .A1(\mem[113][4] ),
    .A2(\mem[114][4] ),
    .A3(\mem[115][4] ),
    .S0(_02616_),
    .S1(_02618_),
    .X(_03080_));
 sky130_fd_sc_hd__mux4_1 _07136_ (.A0(\mem[116][4] ),
    .A1(\mem[117][4] ),
    .A2(\mem[118][4] ),
    .A3(\mem[119][4] ),
    .S0(_02985_),
    .S1(_02623_),
    .X(_03081_));
 sky130_fd_sc_hd__mux4_1 _07137_ (.A0(\mem[120][4] ),
    .A1(\mem[121][4] ),
    .A2(\mem[122][4] ),
    .A3(\mem[123][4] ),
    .S0(_02887_),
    .S1(_02626_),
    .X(_03082_));
 sky130_fd_sc_hd__o22a_1 _07138_ (.A1(_02885_),
    .A2(_03081_),
    .B1(_03082_),
    .B2(_02889_),
    .X(_03083_));
 sky130_fd_sc_hd__o221a_1 _07139_ (.A1(_02612_),
    .A2(_03079_),
    .B1(_03080_),
    .B2(_02884_),
    .C1(_03083_),
    .X(_03084_));
 sky130_fd_sc_hd__o21a_1 _07140_ (.A1(_02611_),
    .A2(_03084_),
    .B1(_02631_),
    .X(_03085_));
 sky130_fd_sc_hd__a32o_1 _07141_ (.A1(_02513_),
    .A2(_03056_),
    .A3(_03070_),
    .B1(_03078_),
    .B2(_03085_),
    .X(_03086_));
 sky130_fd_sc_hd__mux2_1 _07142_ (.A0(_03041_),
    .A1(_03086_),
    .S(_02635_),
    .X(_03087_));
 sky130_fd_sc_hd__clkbuf_1 _07143_ (.A(_03087_),
    .X(_00010_));
 sky130_fd_sc_hd__o21a_1 _07144_ (.A1(\mem[93][5] ),
    .A2(_02640_),
    .B1(_02641_),
    .X(_03088_));
 sky130_fd_sc_hd__or3_1 _07145_ (.A(_02646_),
    .B(_02489_),
    .C(\mem[92][5] ),
    .X(_03089_));
 sky130_fd_sc_hd__o221a_1 _07146_ (.A1(\mem[94][5] ),
    .A2(_02643_),
    .B1(_02644_),
    .B2(\mem[95][5] ),
    .C1(_03089_),
    .X(_03090_));
 sky130_fd_sc_hd__o21a_1 _07147_ (.A1(\mem[80][5] ),
    .A2(_02650_),
    .B1(_02596_),
    .X(_03091_));
 sky130_fd_sc_hd__buf_8 _07148_ (.A(_02442_),
    .X(_03092_));
 sky130_fd_sc_hd__or3b_1 _07149_ (.A(_02656_),
    .B(\mem[82][5] ),
    .C_N(_02492_),
    .X(_03093_));
 sky130_fd_sc_hd__o221a_1 _07150_ (.A1(\mem[81][5] ),
    .A2(_02654_),
    .B1(_03092_),
    .B2(\mem[83][5] ),
    .C1(_03093_),
    .X(_03094_));
 sky130_fd_sc_hd__a22o_1 _07151_ (.A1(_03088_),
    .A2(_03090_),
    .B1(_03091_),
    .B2(_03094_),
    .X(_03095_));
 sky130_fd_sc_hd__o21a_1 _07152_ (.A1(\mem[88][5] ),
    .A2(_02650_),
    .B1(_02662_),
    .X(_03096_));
 sky130_fd_sc_hd__o22a_1 _07153_ (.A1(\mem[89][5] ),
    .A2(_02640_),
    .B1(_02666_),
    .B2(\mem[91][5] ),
    .X(_03097_));
 sky130_fd_sc_hd__o211a_1 _07154_ (.A1(\mem[90][5] ),
    .A2(_02661_),
    .B1(_03096_),
    .C1(_03097_),
    .X(_03098_));
 sky130_fd_sc_hd__or3_1 _07155_ (.A(_02672_),
    .B(_02682_),
    .C(\mem[84][5] ),
    .X(_03099_));
 sky130_fd_sc_hd__o221a_1 _07156_ (.A1(\mem[86][5] ),
    .A2(_02643_),
    .B1(_02655_),
    .B2(\mem[87][5] ),
    .C1(_03099_),
    .X(_03100_));
 sky130_fd_sc_hd__o211a_1 _07157_ (.A1(\mem[85][5] ),
    .A2(_02669_),
    .B1(_03100_),
    .C1(_02677_),
    .X(_03101_));
 sky130_fd_sc_hd__nor4_4 _07158_ (.A(_02638_),
    .B(_03095_),
    .C(_03098_),
    .D(_03101_),
    .Y(_03102_));
 sky130_fd_sc_hd__or3_1 _07159_ (.A(_02681_),
    .B(_02682_),
    .C(\mem[76][5] ),
    .X(_03103_));
 sky130_fd_sc_hd__o221a_1 _07160_ (.A1(\mem[78][5] ),
    .A2(_02643_),
    .B1(_02655_),
    .B2(\mem[79][5] ),
    .C1(_03103_),
    .X(_03104_));
 sky130_fd_sc_hd__o211a_1 _07161_ (.A1(\mem[77][5] ),
    .A2(_02669_),
    .B1(_03104_),
    .C1(_02641_),
    .X(_03105_));
 sky130_fd_sc_hd__o21a_1 _07162_ (.A1(\mem[64][5] ),
    .A2(_02650_),
    .B1(_02652_),
    .X(_03106_));
 sky130_fd_sc_hd__o22a_1 _07163_ (.A1(\mem[65][5] ),
    .A2(_02640_),
    .B1(_02666_),
    .B2(\mem[67][5] ),
    .X(_03107_));
 sky130_fd_sc_hd__o211a_1 _07164_ (.A1(\mem[66][5] ),
    .A2(_02661_),
    .B1(_03106_),
    .C1(_03107_),
    .X(_03108_));
 sky130_fd_sc_hd__or2_1 _07165_ (.A(\mem[72][5] ),
    .B(_02649_),
    .X(_03109_));
 sky130_fd_sc_hd__or3b_1 _07166_ (.A(_02672_),
    .B(\mem[74][5] ),
    .C_N(_02682_),
    .X(_03110_));
 sky130_fd_sc_hd__o221a_1 _07167_ (.A1(\mem[73][5] ),
    .A2(_02654_),
    .B1(_02655_),
    .B2(\mem[75][5] ),
    .C1(_03110_),
    .X(_03111_));
 sky130_fd_sc_hd__o21a_1 _07168_ (.A1(\mem[69][5] ),
    .A2(_02669_),
    .B1(_02465_),
    .X(_03112_));
 sky130_fd_sc_hd__or3_1 _07169_ (.A(_02693_),
    .B(_02674_),
    .C(\mem[68][5] ),
    .X(_03113_));
 sky130_fd_sc_hd__o221a_1 _07170_ (.A1(\mem[70][5] ),
    .A2(_02643_),
    .B1(_02666_),
    .B2(\mem[71][5] ),
    .C1(_03113_),
    .X(_03114_));
 sky130_fd_sc_hd__a32o_1 _07171_ (.A1(_02662_),
    .A2(_03109_),
    .A3(_03111_),
    .B1(_03112_),
    .B2(_03114_),
    .X(_03115_));
 sky130_fd_sc_hd__nor4_4 _07172_ (.A(_02680_),
    .B(_03105_),
    .C(_03108_),
    .D(_03115_),
    .Y(_03116_));
 sky130_fd_sc_hd__mux4_1 _07173_ (.A0(\mem[124][5] ),
    .A1(\mem[125][5] ),
    .A2(\mem[126][5] ),
    .A3(\mem[127][5] ),
    .S0(_02711_),
    .S1(_02699_),
    .X(_03117_));
 sky130_fd_sc_hd__mux4_1 _07174_ (.A0(\mem[112][5] ),
    .A1(\mem[113][5] ),
    .A2(\mem[114][5] ),
    .A3(\mem[115][5] ),
    .S0(_02698_),
    .S1(_02699_),
    .X(_03118_));
 sky130_fd_sc_hd__mux4_1 _07175_ (.A0(\mem[116][5] ),
    .A1(\mem[117][5] ),
    .A2(\mem[118][5] ),
    .A3(\mem[119][5] ),
    .S0(_02681_),
    .S1(_02743_),
    .X(_03119_));
 sky130_fd_sc_hd__mux4_1 _07176_ (.A0(\mem[120][5] ),
    .A1(\mem[121][5] ),
    .A2(\mem[122][5] ),
    .A3(\mem[123][5] ),
    .S0(_02672_),
    .S1(_02704_),
    .X(_03120_));
 sky130_fd_sc_hd__o22a_1 _07177_ (.A1(_02702_),
    .A2(_03119_),
    .B1(_03120_),
    .B2(_02707_),
    .X(_03121_));
 sky130_fd_sc_hd__o221a_1 _07178_ (.A1(_02485_),
    .A2(_03117_),
    .B1(_03118_),
    .B2(_02496_),
    .C1(_03121_),
    .X(_03122_));
 sky130_fd_sc_hd__nor2_1 _07179_ (.A(_02638_),
    .B(_03122_),
    .Y(_03123_));
 sky130_fd_sc_hd__mux4_1 _07180_ (.A0(\mem[100][5] ),
    .A1(\mem[101][5] ),
    .A2(\mem[102][5] ),
    .A3(\mem[103][5] ),
    .S0(_02711_),
    .S1(_02712_),
    .X(_03124_));
 sky130_fd_sc_hd__mux4_1 _07181_ (.A0(\mem[96][5] ),
    .A1(\mem[97][5] ),
    .A2(\mem[98][5] ),
    .A3(\mem[99][5] ),
    .S0(_02711_),
    .S1(_02699_),
    .X(_03125_));
 sky130_fd_sc_hd__a22o_1 _07182_ (.A1(_02677_),
    .A2(_03124_),
    .B1(_03125_),
    .B2(_02652_),
    .X(_03126_));
 sky130_fd_sc_hd__mux4_1 _07183_ (.A0(\mem[108][5] ),
    .A1(\mem[109][5] ),
    .A2(\mem[110][5] ),
    .A3(\mem[111][5] ),
    .S0(_02711_),
    .S1(_02712_),
    .X(_03127_));
 sky130_fd_sc_hd__mux4_1 _07184_ (.A0(\mem[104][5] ),
    .A1(\mem[105][5] ),
    .A2(\mem[106][5] ),
    .A3(\mem[107][5] ),
    .S0(_02428_),
    .S1(_02674_),
    .X(_03128_));
 sky130_fd_sc_hd__or2_1 _07185_ (.A(_02718_),
    .B(_03128_),
    .X(_03129_));
 sky130_fd_sc_hd__o211a_1 _07186_ (.A1(_02716_),
    .A2(_03127_),
    .B1(_03129_),
    .C1(_02721_),
    .X(_03130_));
 sky130_fd_sc_hd__o31ai_1 _07187_ (.A1(_02680_),
    .A2(_03126_),
    .A3(_03130_),
    .B1(_02637_),
    .Y(_03131_));
 sky130_fd_sc_hd__o32a_1 _07188_ (.A1(_02637_),
    .A2(_03102_),
    .A3(_03116_),
    .B1(_03123_),
    .B2(_03131_),
    .X(_03132_));
 sky130_fd_sc_hd__or3_1 _07189_ (.A(_02726_),
    .B(_02673_),
    .C(\mem[28][5] ),
    .X(_03133_));
 sky130_fd_sc_hd__o221a_1 _07190_ (.A1(\mem[30][5] ),
    .A2(_02660_),
    .B1(_02665_),
    .B2(\mem[31][5] ),
    .C1(_03133_),
    .X(_03134_));
 sky130_fd_sc_hd__o211a_1 _07191_ (.A1(\mem[29][5] ),
    .A2(_02640_),
    .B1(_03134_),
    .C1(_02641_),
    .X(_03135_));
 sky130_fd_sc_hd__o21a_1 _07192_ (.A1(\mem[16][5] ),
    .A2(_02649_),
    .B1(_02651_),
    .X(_03136_));
 sky130_fd_sc_hd__o22a_1 _07193_ (.A1(\mem[17][5] ),
    .A2(_02406_),
    .B1(_02644_),
    .B2(\mem[19][5] ),
    .X(_03137_));
 sky130_fd_sc_hd__o211a_1 _07194_ (.A1(\mem[18][5] ),
    .A2(_02661_),
    .B1(_03136_),
    .C1(_03137_),
    .X(_03138_));
 sky130_fd_sc_hd__or2_1 _07195_ (.A(\mem[24][5] ),
    .B(_02649_),
    .X(_03139_));
 sky130_fd_sc_hd__or3b_1 _07196_ (.A(_02671_),
    .B(\mem[26][5] ),
    .C_N(_02673_),
    .X(_03140_));
 sky130_fd_sc_hd__o221a_1 _07197_ (.A1(\mem[25][5] ),
    .A2(_02639_),
    .B1(_02665_),
    .B2(\mem[27][5] ),
    .C1(_03140_),
    .X(_03141_));
 sky130_fd_sc_hd__o21a_1 _07198_ (.A1(\mem[21][5] ),
    .A2(_02737_),
    .B1(_02417_),
    .X(_03142_));
 sky130_fd_sc_hd__or3_1 _07199_ (.A(_02491_),
    .B(_02430_),
    .C(\mem[20][5] ),
    .X(_03143_));
 sky130_fd_sc_hd__o221a_1 _07200_ (.A1(\mem[22][5] ),
    .A2(_02660_),
    .B1(_02665_),
    .B2(\mem[23][5] ),
    .C1(_03143_),
    .X(_03144_));
 sky130_fd_sc_hd__a32o_1 _07201_ (.A1(_02662_),
    .A2(_03139_),
    .A3(_03141_),
    .B1(_03142_),
    .B2(_03144_),
    .X(_03145_));
 sky130_fd_sc_hd__or3_1 _07202_ (.A(_03135_),
    .B(_03138_),
    .C(_03145_),
    .X(_03146_));
 sky130_fd_sc_hd__mux4_1 _07203_ (.A0(\mem[8][5] ),
    .A1(\mem[9][5] ),
    .A2(\mem[10][5] ),
    .A3(\mem[11][5] ),
    .S0(_02646_),
    .S1(_02743_),
    .X(_03147_));
 sky130_fd_sc_hd__or2_1 _07204_ (.A(_02718_),
    .B(_03147_),
    .X(_03148_));
 sky130_fd_sc_hd__mux2_1 _07205_ (.A0(\mem[14][5] ),
    .A1(\mem[15][5] ),
    .S(_02749_),
    .X(_03149_));
 sky130_fd_sc_hd__mux2_1 _07206_ (.A0(\mem[12][5] ),
    .A1(\mem[13][5] ),
    .S(_02428_),
    .X(_03150_));
 sky130_fd_sc_hd__and2b_1 _07207_ (.A_N(_02747_),
    .B(_03150_),
    .X(_03151_));
 sky130_fd_sc_hd__a211o_1 _07208_ (.A1(_02748_),
    .A2(_03149_),
    .B1(_03151_),
    .C1(_02716_),
    .X(_03152_));
 sky130_fd_sc_hd__mux2_2 _07209_ (.A0(\mem[6][5] ),
    .A1(\mem[7][5] ),
    .S(_02749_),
    .X(_03153_));
 sky130_fd_sc_hd__mux2_1 _07210_ (.A0(\mem[4][5] ),
    .A1(\mem[5][5] ),
    .S(_02428_),
    .X(_03154_));
 sky130_fd_sc_hd__and2b_1 _07211_ (.A_N(_02712_),
    .B(_03154_),
    .X(_03155_));
 sky130_fd_sc_hd__a211o_1 _07212_ (.A1(_02748_),
    .A2(_03153_),
    .B1(_03155_),
    .C1(_02716_),
    .X(_03156_));
 sky130_fd_sc_hd__mux4_1 _07213_ (.A0(\mem[0][5] ),
    .A1(\mem[1][5] ),
    .A2(\mem[2][5] ),
    .A3(\mem[3][5] ),
    .S0(_02693_),
    .S1(_02704_),
    .X(_03157_));
 sky130_fd_sc_hd__o21ba_1 _07214_ (.A1(_02718_),
    .A2(_03157_),
    .B1_N(_02479_),
    .X(_03158_));
 sky130_fd_sc_hd__a32o_1 _07215_ (.A1(_02721_),
    .A2(_03148_),
    .A3(_03152_),
    .B1(_03156_),
    .B2(_03158_),
    .X(_03159_));
 sky130_fd_sc_hd__a221o_1 _07216_ (.A1(_02725_),
    .A2(_03146_),
    .B1(_03159_),
    .B2(_02761_),
    .C1(_02634_),
    .X(_03160_));
 sky130_fd_sc_hd__mux4_1 _07217_ (.A0(\mem[60][5] ),
    .A1(\mem[61][5] ),
    .A2(\mem[62][5] ),
    .A3(\mem[63][5] ),
    .S0(_02698_),
    .S1(_02699_),
    .X(_03161_));
 sky130_fd_sc_hd__mux4_1 _07218_ (.A0(\mem[48][5] ),
    .A1(\mem[49][5] ),
    .A2(\mem[50][5] ),
    .A3(\mem[51][5] ),
    .S0(_02698_),
    .S1(_02748_),
    .X(_03162_));
 sky130_fd_sc_hd__mux4_1 _07219_ (.A0(\mem[52][5] ),
    .A1(\mem[53][5] ),
    .A2(\mem[54][5] ),
    .A3(\mem[55][5] ),
    .S0(_02693_),
    .S1(_02747_),
    .X(_03163_));
 sky130_fd_sc_hd__mux4_1 _07220_ (.A0(\mem[56][5] ),
    .A1(\mem[57][5] ),
    .A2(\mem[58][5] ),
    .A3(\mem[59][5] ),
    .S0(_02749_),
    .S1(_02747_),
    .X(_03164_));
 sky130_fd_sc_hd__o22a_1 _07221_ (.A1(_02702_),
    .A2(_03163_),
    .B1(_03164_),
    .B2(_02707_),
    .X(_03165_));
 sky130_fd_sc_hd__o221a_1 _07222_ (.A1(_02485_),
    .A2(_03161_),
    .B1(_03162_),
    .B2(_02496_),
    .C1(_03165_),
    .X(_03166_));
 sky130_fd_sc_hd__mux4_1 _07223_ (.A0(\mem[36][5] ),
    .A1(\mem[37][5] ),
    .A2(\mem[38][5] ),
    .A3(\mem[39][5] ),
    .S0(_02656_),
    .S1(_02743_),
    .X(_03167_));
 sky130_fd_sc_hd__mux4_1 _07224_ (.A0(\mem[32][5] ),
    .A1(\mem[33][5] ),
    .A2(\mem[34][5] ),
    .A3(\mem[35][5] ),
    .S0(_02681_),
    .S1(_02704_),
    .X(_03168_));
 sky130_fd_sc_hd__a22o_1 _07225_ (.A1(_02677_),
    .A2(_03167_),
    .B1(_03168_),
    .B2(_02652_),
    .X(_03169_));
 sky130_fd_sc_hd__mux4_1 _07226_ (.A0(\mem[44][5] ),
    .A1(\mem[45][5] ),
    .A2(\mem[46][5] ),
    .A3(\mem[47][5] ),
    .S0(_02656_),
    .S1(_02743_),
    .X(_03170_));
 sky130_fd_sc_hd__mux4_1 _07227_ (.A0(\mem[40][5] ),
    .A1(\mem[41][5] ),
    .A2(\mem[42][5] ),
    .A3(\mem[43][5] ),
    .S0(_02645_),
    .S1(_02430_),
    .X(_03171_));
 sky130_fd_sc_hd__or2_1 _07228_ (.A(_02475_),
    .B(_03171_),
    .X(_03172_));
 sky130_fd_sc_hd__o211a_1 _07229_ (.A1(_02472_),
    .A2(_03170_),
    .B1(_03172_),
    .C1(_02721_),
    .X(_03173_));
 sky130_fd_sc_hd__or3_1 _07230_ (.A(_02680_),
    .B(_03169_),
    .C(_03173_),
    .X(_03174_));
 sky130_fd_sc_hd__o211a_1 _07231_ (.A1(_02638_),
    .A2(_03166_),
    .B1(_03174_),
    .C1(_02637_),
    .X(_03175_));
 sky130_fd_sc_hd__o2bb2a_1 _07232_ (.A1_N(_02635_),
    .A2_N(_03132_),
    .B1(_03160_),
    .B2(_03175_),
    .X(_00011_));
 sky130_fd_sc_hd__o21a_1 _07233_ (.A1(\mem[29][6] ),
    .A2(_02363_),
    .B1(_02366_),
    .X(_03176_));
 sky130_fd_sc_hd__or3_1 _07234_ (.A(_02374_),
    .B(_02779_),
    .C(\mem[28][6] ),
    .X(_03177_));
 sky130_fd_sc_hd__o221a_1 _07235_ (.A1(\mem[30][6] ),
    .A2(_02995_),
    .B1(_02372_),
    .B2(\mem[31][6] ),
    .C1(_03177_),
    .X(_03178_));
 sky130_fd_sc_hd__o21a_1 _07236_ (.A1(\mem[16][6] ),
    .A2(_02380_),
    .B1(_02383_),
    .X(_03179_));
 sky130_fd_sc_hd__or3b_1 _07237_ (.A(_02387_),
    .B(\mem[18][6] ),
    .C_N(_02783_),
    .X(_03180_));
 sky130_fd_sc_hd__o221a_1 _07238_ (.A1(\mem[17][6] ),
    .A2(_02899_),
    .B1(_02386_),
    .B2(\mem[19][6] ),
    .C1(_03180_),
    .X(_03181_));
 sky130_fd_sc_hd__a22o_1 _07239_ (.A1(_03176_),
    .A2(_03178_),
    .B1(_03179_),
    .B2(_03181_),
    .X(_03182_));
 sky130_fd_sc_hd__o21a_1 _07240_ (.A1(\mem[24][6] ),
    .A2(_02788_),
    .B1(_02397_),
    .X(_03183_));
 sky130_fd_sc_hd__o22a_1 _07241_ (.A1(\mem[25][6] ),
    .A2(_02790_),
    .B1(_02401_),
    .B2(\mem[27][6] ),
    .X(_03184_));
 sky130_fd_sc_hd__o211a_1 _07242_ (.A1(\mem[26][6] ),
    .A2(_02787_),
    .B1(_03183_),
    .C1(_03184_),
    .X(_03185_));
 sky130_fd_sc_hd__or3_1 _07243_ (.A(_02793_),
    .B(_02412_),
    .C(\mem[20][6] ),
    .X(_03186_));
 sky130_fd_sc_hd__o221a_1 _07244_ (.A1(\mem[22][6] ),
    .A2(_02407_),
    .B1(_02409_),
    .B2(\mem[23][6] ),
    .C1(_03186_),
    .X(_03187_));
 sky130_fd_sc_hd__o211a_1 _07245_ (.A1(\mem[21][6] ),
    .A2(_02406_),
    .B1(_03187_),
    .C1(_02417_),
    .X(_03188_));
 sky130_fd_sc_hd__or4_2 _07246_ (.A(_02993_),
    .B(_03182_),
    .C(_03185_),
    .D(_03188_),
    .X(_03189_));
 sky130_fd_sc_hd__or3_1 _07247_ (.A(_02802_),
    .B(_02803_),
    .C(\mem[12][6] ),
    .X(_03190_));
 sky130_fd_sc_hd__o221a_1 _07248_ (.A1(\mem[14][6] ),
    .A2(_02800_),
    .B1(_03009_),
    .B2(\mem[15][6] ),
    .C1(_03190_),
    .X(_03191_));
 sky130_fd_sc_hd__o211a_1 _07249_ (.A1(\mem[13][6] ),
    .A2(_02799_),
    .B1(_03191_),
    .C1(_02806_),
    .X(_03192_));
 sky130_fd_sc_hd__o21a_1 _07250_ (.A1(\mem[0][6] ),
    .A2(_02438_),
    .B1(_03013_),
    .X(_03193_));
 sky130_fd_sc_hd__o22a_1 _07251_ (.A1(\mem[1][6] ),
    .A2(_02441_),
    .B1(_02914_),
    .B2(\mem[3][6] ),
    .X(_03194_));
 sky130_fd_sc_hd__o211a_1 _07252_ (.A1(\mem[2][6] ),
    .A2(_02437_),
    .B1(_03193_),
    .C1(_03194_),
    .X(_03195_));
 sky130_fd_sc_hd__or2_1 _07253_ (.A(\mem[8][6] ),
    .B(_02917_),
    .X(_03196_));
 sky130_fd_sc_hd__or3b_1 _07254_ (.A(_02815_),
    .B(\mem[10][6] ),
    .C_N(_02816_),
    .X(_03197_));
 sky130_fd_sc_hd__o221a_1 _07255_ (.A1(\mem[9][6] ),
    .A2(_02736_),
    .B1(_02814_),
    .B2(\mem[11][6] ),
    .C1(_03197_),
    .X(_03198_));
 sky130_fd_sc_hd__o21a_1 _07256_ (.A1(\mem[5][6] ),
    .A2(_02819_),
    .B1(_02416_),
    .X(_03199_));
 sky130_fd_sc_hd__or3_1 _07257_ (.A(_02447_),
    .B(_02584_),
    .C(\mem[4][6] ),
    .X(_03200_));
 sky130_fd_sc_hd__o221a_1 _07258_ (.A1(\mem[6][6] ),
    .A2(_02445_),
    .B1(_02446_),
    .B2(\mem[7][6] ),
    .C1(_03200_),
    .X(_03201_));
 sky130_fd_sc_hd__a32o_1 _07259_ (.A1(_02811_),
    .A2(_03196_),
    .A3(_03198_),
    .B1(_03199_),
    .B2(_03201_),
    .X(_03202_));
 sky130_fd_sc_hd__or4_1 _07260_ (.A(_02798_),
    .B(_03192_),
    .C(_03195_),
    .D(_03202_),
    .X(_03203_));
 sky130_fd_sc_hd__mux4_1 _07261_ (.A0(\mem[36][6] ),
    .A1(\mem[37][6] ),
    .A2(\mem[38][6] ),
    .A3(\mem[39][6] ),
    .S0(_02826_),
    .S1(_02926_),
    .X(_03204_));
 sky130_fd_sc_hd__mux4_1 _07262_ (.A0(\mem[32][6] ),
    .A1(\mem[33][6] ),
    .A2(\mem[34][6] ),
    .A3(\mem[35][6] ),
    .S0(_02928_),
    .S1(_02929_),
    .X(_03205_));
 sky130_fd_sc_hd__a22o_1 _07263_ (.A1(_02450_),
    .A2(_03204_),
    .B1(_03205_),
    .B2(_02596_),
    .X(_03206_));
 sky130_fd_sc_hd__mux4_1 _07264_ (.A0(\mem[44][6] ),
    .A1(\mem[45][6] ),
    .A2(\mem[46][6] ),
    .A3(\mem[47][6] ),
    .S0(_02467_),
    .S1(_02468_),
    .X(_03207_));
 sky130_fd_sc_hd__mux4_1 _07265_ (.A0(\mem[40][6] ),
    .A1(\mem[41][6] ),
    .A2(\mem[42][6] ),
    .A3(\mem[43][6] ),
    .S0(_02457_),
    .S1(_02605_),
    .X(_03208_));
 sky130_fd_sc_hd__or2_1 _07266_ (.A(_02475_),
    .B(_03208_),
    .X(_03209_));
 sky130_fd_sc_hd__o211a_1 _07267_ (.A1(_02472_),
    .A2(_03207_),
    .B1(_03209_),
    .C1(_02479_),
    .X(_03210_));
 sky130_fd_sc_hd__or3_4 _07268_ (.A(_02453_),
    .B(_03206_),
    .C(_03210_),
    .X(_03211_));
 sky130_fd_sc_hd__mux4_1 _07269_ (.A0(\mem[60][6] ),
    .A1(\mem[61][6] ),
    .A2(\mem[62][6] ),
    .A3(\mem[63][6] ),
    .S0(_02487_),
    .S1(_02489_),
    .X(_03212_));
 sky130_fd_sc_hd__mux4_1 _07270_ (.A0(\mem[48][6] ),
    .A1(\mem[49][6] ),
    .A2(\mem[50][6] ),
    .A3(\mem[51][6] ),
    .S0(_02491_),
    .S1(_02746_),
    .X(_03213_));
 sky130_fd_sc_hd__mux4_1 _07271_ (.A0(\mem[52][6] ),
    .A1(\mem[53][6] ),
    .A2(\mem[54][6] ),
    .A3(\mem[55][6] ),
    .S0(_02427_),
    .S1(_02837_),
    .X(_03214_));
 sky130_fd_sc_hd__mux4_1 _07272_ (.A0(\mem[56][6] ),
    .A1(\mem[57][6] ),
    .A2(\mem[58][6] ),
    .A3(\mem[59][6] ),
    .S0(_02625_),
    .S1(_02503_),
    .X(_03215_));
 sky130_fd_sc_hd__o22a_1 _07273_ (.A1(_02621_),
    .A2(_03214_),
    .B1(_03215_),
    .B2(_02628_),
    .X(_03216_));
 sky130_fd_sc_hd__o221a_1 _07274_ (.A1(_03033_),
    .A2(_03212_),
    .B1(_03213_),
    .B2(_02620_),
    .C1(_03216_),
    .X(_03217_));
 sky130_fd_sc_hd__o21a_1 _07275_ (.A1(_02482_),
    .A2(_03217_),
    .B1(_02510_),
    .X(_03218_));
 sky130_fd_sc_hd__a32o_1 _07276_ (.A1(_02356_),
    .A2(_03189_),
    .A3(_03203_),
    .B1(_03211_),
    .B2(_03218_),
    .X(_03219_));
 sky130_fd_sc_hd__o21a_1 _07277_ (.A1(\mem[93][6] ),
    .A2(_02565_),
    .B1(_02422_),
    .X(_03220_));
 sky130_fd_sc_hd__or3_1 _07278_ (.A(_02387_),
    .B(_02389_),
    .C(\mem[92][6] ),
    .X(_03221_));
 sky130_fd_sc_hd__o221a_1 _07279_ (.A1(\mem[94][6] ),
    .A2(_02370_),
    .B1(_02386_),
    .B2(\mem[95][6] ),
    .C1(_03221_),
    .X(_03222_));
 sky130_fd_sc_hd__o21a_1 _07280_ (.A1(\mem[80][6] ),
    .A2(_02438_),
    .B1(_02455_),
    .X(_03223_));
 sky130_fd_sc_hd__buf_4 _07281_ (.A(_02388_),
    .X(_03224_));
 sky130_fd_sc_hd__or3b_1 _07282_ (.A(_02815_),
    .B(\mem[82][6] ),
    .C_N(_03224_),
    .X(_03225_));
 sky130_fd_sc_hd__o221a_1 _07283_ (.A1(\mem[81][6] ),
    .A2(_02736_),
    .B1(_02814_),
    .B2(\mem[83][6] ),
    .C1(_03225_),
    .X(_03226_));
 sky130_fd_sc_hd__a22o_1 _07284_ (.A1(_03220_),
    .A2(_03222_),
    .B1(_03223_),
    .B2(_03226_),
    .X(_03227_));
 sky130_fd_sc_hd__o21a_1 _07285_ (.A1(\mem[88][6] ),
    .A2(_02649_),
    .B1(_02439_),
    .X(_03228_));
 sky130_fd_sc_hd__o22a_1 _07286_ (.A1(\mem[89][6] ),
    .A2(_02405_),
    .B1(_02442_),
    .B2(\mem[91][6] ),
    .X(_03229_));
 sky130_fd_sc_hd__o211a_1 _07287_ (.A1(\mem[90][6] ),
    .A2(_02437_),
    .B1(_03228_),
    .C1(_03229_),
    .X(_03230_));
 sky130_fd_sc_hd__buf_4 _07288_ (.A(_02408_),
    .X(_03231_));
 sky130_fd_sc_hd__or3_1 _07289_ (.A(_02427_),
    .B(_02429_),
    .C(\mem[84][6] ),
    .X(_03232_));
 sky130_fd_sc_hd__o221a_1 _07290_ (.A1(\mem[86][6] ),
    .A2(_02393_),
    .B1(_03231_),
    .B2(\mem[87][6] ),
    .C1(_03232_),
    .X(_03233_));
 sky130_fd_sc_hd__o211a_1 _07291_ (.A1(\mem[85][6] ),
    .A2(_02737_),
    .B1(_03233_),
    .C1(_02450_),
    .X(_03234_));
 sky130_fd_sc_hd__or4_2 _07292_ (.A(_02358_),
    .B(_03227_),
    .C(_03230_),
    .D(_03234_),
    .X(_03235_));
 sky130_fd_sc_hd__or3_1 _07293_ (.A(_02486_),
    .B(_03224_),
    .C(\mem[76][6] ),
    .X(_03236_));
 sky130_fd_sc_hd__o221a_1 _07294_ (.A1(\mem[78][6] ),
    .A2(_02956_),
    .B1(_02814_),
    .B2(\mem[79][6] ),
    .C1(_03236_),
    .X(_03237_));
 sky130_fd_sc_hd__o211a_1 _07295_ (.A1(\mem[77][6] ),
    .A2(_02955_),
    .B1(_03237_),
    .C1(_02641_),
    .X(_03238_));
 sky130_fd_sc_hd__o21a_1 _07296_ (.A1(\mem[64][6] ),
    .A2(_02438_),
    .B1(_02455_),
    .X(_03239_));
 sky130_fd_sc_hd__o22a_1 _07297_ (.A1(\mem[65][6] ),
    .A2(_02405_),
    .B1(_02442_),
    .B2(\mem[67][6] ),
    .X(_03240_));
 sky130_fd_sc_hd__o211a_1 _07298_ (.A1(\mem[66][6] ),
    .A2(_02437_),
    .B1(_03239_),
    .C1(_03240_),
    .X(_03241_));
 sky130_fd_sc_hd__or2_1 _07299_ (.A(\mem[72][6] ),
    .B(_02812_),
    .X(_03242_));
 sky130_fd_sc_hd__or3b_1 _07300_ (.A(_02486_),
    .B(\mem[74][6] ),
    .C_N(_03224_),
    .X(_03243_));
 sky130_fd_sc_hd__o221a_1 _07301_ (.A1(\mem[73][6] ),
    .A2(_03042_),
    .B1(_02664_),
    .B2(\mem[75][6] ),
    .C1(_03243_),
    .X(_03244_));
 sky130_fd_sc_hd__o21a_1 _07302_ (.A1(\mem[69][6] ),
    .A2(_02819_),
    .B1(_02416_),
    .X(_03245_));
 sky130_fd_sc_hd__or3_1 _07303_ (.A(_02985_),
    .B(_02429_),
    .C(\mem[68][6] ),
    .X(_03246_));
 sky130_fd_sc_hd__o221a_1 _07304_ (.A1(\mem[70][6] ),
    .A2(_02393_),
    .B1(_03231_),
    .B2(\mem[71][6] ),
    .C1(_03246_),
    .X(_03247_));
 sky130_fd_sc_hd__a32o_1 _07305_ (.A1(_02662_),
    .A2(_03242_),
    .A3(_03244_),
    .B1(_03245_),
    .B2(_03247_),
    .X(_03248_));
 sky130_fd_sc_hd__or4_2 _07306_ (.A(_02421_),
    .B(_03238_),
    .C(_03241_),
    .D(_03248_),
    .X(_03249_));
 sky130_fd_sc_hd__mux4_1 _07307_ (.A0(\mem[104][6] ),
    .A1(\mem[105][6] ),
    .A2(\mem[106][6] ),
    .A3(\mem[107][6] ),
    .S0(_02670_),
    .S1(_02488_),
    .X(_03250_));
 sky130_fd_sc_hd__or2_1 _07308_ (.A(_02475_),
    .B(_03250_),
    .X(_03251_));
 sky130_fd_sc_hd__mux4_1 _07309_ (.A0(\mem[108][6] ),
    .A1(\mem[109][6] ),
    .A2(\mem[110][6] ),
    .A3(\mem[111][6] ),
    .S0(_02374_),
    .S1(_02488_),
    .X(_03252_));
 sky130_fd_sc_hd__or2_1 _07310_ (.A(_02598_),
    .B(_03252_),
    .X(_03253_));
 sky130_fd_sc_hd__mux4_1 _07311_ (.A0(\mem[100][6] ),
    .A1(\mem[101][6] ),
    .A2(\mem[102][6] ),
    .A3(\mem[103][6] ),
    .S0(_02432_),
    .S1(_02488_),
    .X(_03254_));
 sky130_fd_sc_hd__mux4_1 _07312_ (.A0(\mem[96][6] ),
    .A1(\mem[97][6] ),
    .A2(\mem[98][6] ),
    .A3(\mem[99][6] ),
    .S0(_02411_),
    .S1(_02617_),
    .X(_03255_));
 sky130_fd_sc_hd__a22o_1 _07313_ (.A1(_02464_),
    .A2(_03254_),
    .B1(_03255_),
    .B2(_02455_),
    .X(_03256_));
 sky130_fd_sc_hd__a31o_1 _07314_ (.A1(_02479_),
    .A2(_03251_),
    .A3(_03253_),
    .B1(_03256_),
    .X(_03257_));
 sky130_fd_sc_hd__mux4_1 _07315_ (.A0(\mem[116][6] ),
    .A1(\mem[117][6] ),
    .A2(\mem[118][6] ),
    .A3(\mem[119][6] ),
    .S0(_02502_),
    .S1(_02503_),
    .X(_03258_));
 sky130_fd_sc_hd__mux4_1 _07316_ (.A0(\mem[120][6] ),
    .A1(\mem[121][6] ),
    .A2(\mem[122][6] ),
    .A3(\mem[123][6] ),
    .S0(_02502_),
    .S1(_02673_),
    .X(_03259_));
 sky130_fd_sc_hd__o22a_1 _07317_ (.A1(_02498_),
    .A2(_03258_),
    .B1(_03259_),
    .B2(_02506_),
    .X(_03260_));
 sky130_fd_sc_hd__mux4_1 _07318_ (.A0(\mem[124][6] ),
    .A1(\mem[125][6] ),
    .A2(\mem[126][6] ),
    .A3(\mem[127][6] ),
    .S0(_02427_),
    .S1(_02499_),
    .X(_03261_));
 sky130_fd_sc_hd__mux4_1 _07319_ (.A0(\mem[112][6] ),
    .A1(\mem[113][6] ),
    .A2(\mem[114][6] ),
    .A3(\mem[115][6] ),
    .S0(_02502_),
    .S1(_02673_),
    .X(_03262_));
 sky130_fd_sc_hd__o22a_1 _07320_ (.A1(_02484_),
    .A2(_03261_),
    .B1(_03262_),
    .B2(_02495_),
    .X(_03263_));
 sky130_fd_sc_hd__a21o_1 _07321_ (.A1(_03260_),
    .A2(_03263_),
    .B1(_02357_),
    .X(_03264_));
 sky130_fd_sc_hd__o211a_1 _07322_ (.A1(_02453_),
    .A2(_03257_),
    .B1(_03264_),
    .C1(_02509_),
    .X(_03265_));
 sky130_fd_sc_hd__a31o_1 _07323_ (.A1(_02356_),
    .A2(_03235_),
    .A3(_03249_),
    .B1(_03265_),
    .X(_03266_));
 sky130_fd_sc_hd__mux2_1 _07324_ (.A0(_03219_),
    .A1(_03266_),
    .S(_02635_),
    .X(_03267_));
 sky130_fd_sc_hd__clkbuf_1 _07325_ (.A(_03267_),
    .X(_00012_));
 sky130_fd_sc_hd__o21a_1 _07326_ (.A1(\mem[29][7] ),
    .A2(_02363_),
    .B1(_02366_),
    .X(_03268_));
 sky130_fd_sc_hd__or3_1 _07327_ (.A(_02520_),
    .B(_02779_),
    .C(\mem[28][7] ),
    .X(_03269_));
 sky130_fd_sc_hd__o221a_1 _07328_ (.A1(\mem[30][7] ),
    .A2(_02995_),
    .B1(_02372_),
    .B2(\mem[31][7] ),
    .C1(_03269_),
    .X(_03270_));
 sky130_fd_sc_hd__o21a_1 _07329_ (.A1(\mem[16][7] ),
    .A2(_02380_),
    .B1(_02383_),
    .X(_03271_));
 sky130_fd_sc_hd__or3b_1 _07330_ (.A(_02387_),
    .B(\mem[18][7] ),
    .C_N(_02783_),
    .X(_03272_));
 sky130_fd_sc_hd__o221a_1 _07331_ (.A1(\mem[17][7] ),
    .A2(_02899_),
    .B1(_02528_),
    .B2(\mem[19][7] ),
    .C1(_03272_),
    .X(_03273_));
 sky130_fd_sc_hd__a22o_1 _07332_ (.A1(_03268_),
    .A2(_03270_),
    .B1(_03271_),
    .B2(_03273_),
    .X(_03274_));
 sky130_fd_sc_hd__o21a_1 _07333_ (.A1(\mem[24][7] ),
    .A2(_02788_),
    .B1(_02397_),
    .X(_03275_));
 sky130_fd_sc_hd__o22a_1 _07334_ (.A1(\mem[25][7] ),
    .A2(_02790_),
    .B1(_02401_),
    .B2(\mem[27][7] ),
    .X(_03276_));
 sky130_fd_sc_hd__o211a_1 _07335_ (.A1(\mem[26][7] ),
    .A2(_02787_),
    .B1(_03275_),
    .C1(_03276_),
    .X(_03277_));
 sky130_fd_sc_hd__or3_1 _07336_ (.A(_02793_),
    .B(_02412_),
    .C(\mem[20][7] ),
    .X(_03278_));
 sky130_fd_sc_hd__o221a_1 _07337_ (.A1(\mem[22][7] ),
    .A2(_02543_),
    .B1(_02409_),
    .B2(\mem[23][7] ),
    .C1(_03278_),
    .X(_03279_));
 sky130_fd_sc_hd__o211a_1 _07338_ (.A1(\mem[21][7] ),
    .A2(_02542_),
    .B1(_03279_),
    .C1(_02417_),
    .X(_03280_));
 sky130_fd_sc_hd__or4_2 _07339_ (.A(_02993_),
    .B(_03274_),
    .C(_03277_),
    .D(_03280_),
    .X(_03281_));
 sky130_fd_sc_hd__or3_1 _07340_ (.A(_02802_),
    .B(_02803_),
    .C(\mem[12][7] ),
    .X(_03282_));
 sky130_fd_sc_hd__o221a_1 _07341_ (.A1(\mem[14][7] ),
    .A2(_02800_),
    .B1(_03009_),
    .B2(\mem[15][7] ),
    .C1(_03282_),
    .X(_03283_));
 sky130_fd_sc_hd__o211a_1 _07342_ (.A1(\mem[13][7] ),
    .A2(_02799_),
    .B1(_03283_),
    .C1(_02806_),
    .X(_03284_));
 sky130_fd_sc_hd__o21a_1 _07343_ (.A1(\mem[0][7] ),
    .A2(_02562_),
    .B1(_03013_),
    .X(_03285_));
 sky130_fd_sc_hd__o22a_1 _07344_ (.A1(\mem[1][7] ),
    .A2(_02441_),
    .B1(_02914_),
    .B2(\mem[3][7] ),
    .X(_03286_));
 sky130_fd_sc_hd__o211a_1 _07345_ (.A1(\mem[2][7] ),
    .A2(_02561_),
    .B1(_03285_),
    .C1(_03286_),
    .X(_03287_));
 sky130_fd_sc_hd__or2_1 _07346_ (.A(\mem[8][7] ),
    .B(_02917_),
    .X(_03288_));
 sky130_fd_sc_hd__or3b_1 _07347_ (.A(_02815_),
    .B(\mem[10][7] ),
    .C_N(_02816_),
    .X(_03289_));
 sky130_fd_sc_hd__o221a_1 _07348_ (.A1(\mem[9][7] ),
    .A2(_02736_),
    .B1(_02814_),
    .B2(\mem[11][7] ),
    .C1(_03289_),
    .X(_03290_));
 sky130_fd_sc_hd__o21a_1 _07349_ (.A1(\mem[5][7] ),
    .A2(_02819_),
    .B1(_02579_),
    .X(_03291_));
 sky130_fd_sc_hd__or3_1 _07350_ (.A(_02447_),
    .B(_02584_),
    .C(\mem[4][7] ),
    .X(_03292_));
 sky130_fd_sc_hd__o221a_2 _07351_ (.A1(\mem[6][7] ),
    .A2(_02445_),
    .B1(_02446_),
    .B2(\mem[7][7] ),
    .C1(_03292_),
    .X(_03293_));
 sky130_fd_sc_hd__a32o_1 _07352_ (.A1(_02811_),
    .A2(_03288_),
    .A3(_03290_),
    .B1(_03291_),
    .B2(_03293_),
    .X(_03294_));
 sky130_fd_sc_hd__or4_1 _07353_ (.A(_02798_),
    .B(_03284_),
    .C(_03287_),
    .D(_03294_),
    .X(_03295_));
 sky130_fd_sc_hd__mux4_1 _07354_ (.A0(\mem[32][7] ),
    .A1(\mem[33][7] ),
    .A2(\mem[34][7] ),
    .A3(\mem[35][7] ),
    .S0(_02826_),
    .S1(_02926_),
    .X(_03296_));
 sky130_fd_sc_hd__mux4_1 _07355_ (.A0(\mem[36][7] ),
    .A1(\mem[37][7] ),
    .A2(\mem[38][7] ),
    .A3(\mem[39][7] ),
    .S0(_02928_),
    .S1(_02929_),
    .X(_03297_));
 sky130_fd_sc_hd__a22o_1 _07356_ (.A1(_02456_),
    .A2(_03296_),
    .B1(_03297_),
    .B2(_02465_),
    .X(_03298_));
 sky130_fd_sc_hd__mux4_1 _07357_ (.A0(\mem[44][7] ),
    .A1(\mem[45][7] ),
    .A2(\mem[46][7] ),
    .A3(\mem[47][7] ),
    .S0(_02600_),
    .S1(_02468_),
    .X(_03299_));
 sky130_fd_sc_hd__mux4_1 _07358_ (.A0(\mem[40][7] ),
    .A1(\mem[41][7] ),
    .A2(\mem[42][7] ),
    .A3(\mem[43][7] ),
    .S0(_02457_),
    .S1(_02605_),
    .X(_03300_));
 sky130_fd_sc_hd__or2_1 _07359_ (.A(_02603_),
    .B(_03300_),
    .X(_03301_));
 sky130_fd_sc_hd__o211a_1 _07360_ (.A1(_02472_),
    .A2(_03299_),
    .B1(_03301_),
    .C1(_02479_),
    .X(_03302_));
 sky130_fd_sc_hd__or3_2 _07361_ (.A(_02453_),
    .B(_03298_),
    .C(_03302_),
    .X(_03303_));
 sky130_fd_sc_hd__mux4_1 _07362_ (.A0(\mem[60][7] ),
    .A1(\mem[61][7] ),
    .A2(\mem[62][7] ),
    .A3(\mem[63][7] ),
    .S0(_02487_),
    .S1(_02489_),
    .X(_03304_));
 sky130_fd_sc_hd__mux4_1 _07363_ (.A0(\mem[48][7] ),
    .A1(\mem[49][7] ),
    .A2(\mem[50][7] ),
    .A3(\mem[51][7] ),
    .S0(_02491_),
    .S1(_02746_),
    .X(_03305_));
 sky130_fd_sc_hd__mux4_1 _07364_ (.A0(\mem[52][7] ),
    .A1(\mem[53][7] ),
    .A2(\mem[54][7] ),
    .A3(\mem[55][7] ),
    .S0(_02622_),
    .S1(_02837_),
    .X(_03306_));
 sky130_fd_sc_hd__mux4_1 _07365_ (.A0(\mem[56][7] ),
    .A1(\mem[57][7] ),
    .A2(\mem[58][7] ),
    .A3(\mem[59][7] ),
    .S0(_02625_),
    .S1(_02503_),
    .X(_03307_));
 sky130_fd_sc_hd__o22a_1 _07366_ (.A1(_02621_),
    .A2(_03306_),
    .B1(_03307_),
    .B2(_02628_),
    .X(_03308_));
 sky130_fd_sc_hd__o221a_1 _07367_ (.A1(_03033_),
    .A2(_03304_),
    .B1(_03305_),
    .B2(_02620_),
    .C1(_03308_),
    .X(_03309_));
 sky130_fd_sc_hd__o21a_1 _07368_ (.A1(_02482_),
    .A2(_03309_),
    .B1(_02510_),
    .X(_03310_));
 sky130_fd_sc_hd__a32o_1 _07369_ (.A1(_02356_),
    .A2(_03281_),
    .A3(_03295_),
    .B1(_03303_),
    .B2(_03310_),
    .X(_03311_));
 sky130_fd_sc_hd__o21a_1 _07370_ (.A1(\mem[93][7] ),
    .A2(_03042_),
    .B1(_02516_),
    .X(_03312_));
 sky130_fd_sc_hd__or3_1 _07371_ (.A(_02466_),
    .B(_02521_),
    .C(\mem[92][7] ),
    .X(_03313_));
 sky130_fd_sc_hd__o221a_1 _07372_ (.A1(\mem[94][7] ),
    .A2(_02518_),
    .B1(_02519_),
    .B2(\mem[95][7] ),
    .C1(_03313_),
    .X(_03314_));
 sky130_fd_sc_hd__o21a_1 _07373_ (.A1(\mem[80][7] ),
    .A2(_02812_),
    .B1(_02525_),
    .X(_03315_));
 sky130_fd_sc_hd__or3b_1 _07374_ (.A(_02670_),
    .B(\mem[82][7] ),
    .C_N(_02530_),
    .X(_03316_));
 sky130_fd_sc_hd__o221a_1 _07375_ (.A1(\mem[81][7] ),
    .A2(_02527_),
    .B1(_02424_),
    .B2(\mem[83][7] ),
    .C1(_03316_),
    .X(_03317_));
 sky130_fd_sc_hd__a22o_1 _07376_ (.A1(_03312_),
    .A2(_03314_),
    .B1(_03315_),
    .B2(_03317_),
    .X(_03318_));
 sky130_fd_sc_hd__o21a_1 _07377_ (.A1(\mem[88][7] ),
    .A2(_02535_),
    .B1(_02536_),
    .X(_03319_));
 sky130_fd_sc_hd__o22a_1 _07378_ (.A1(\mem[89][7] ),
    .A2(_02538_),
    .B1(_02539_),
    .B2(\mem[91][7] ),
    .X(_03320_));
 sky130_fd_sc_hd__o211a_1 _07379_ (.A1(\mem[90][7] ),
    .A2(_02534_),
    .B1(_03319_),
    .C1(_03320_),
    .X(_03321_));
 sky130_fd_sc_hd__or3_1 _07380_ (.A(_02545_),
    .B(_02546_),
    .C(\mem[84][7] ),
    .X(_03322_));
 sky130_fd_sc_hd__o221a_1 _07381_ (.A1(\mem[86][7] ),
    .A2(_02956_),
    .B1(_02664_),
    .B2(\mem[87][7] ),
    .C1(_03322_),
    .X(_03323_));
 sky130_fd_sc_hd__o211a_1 _07382_ (.A1(\mem[85][7] ),
    .A2(_02955_),
    .B1(_03323_),
    .C1(_02464_),
    .X(_03324_));
 sky130_fd_sc_hd__or4_4 _07383_ (.A(_02514_),
    .B(_03318_),
    .C(_03321_),
    .D(_03324_),
    .X(_03325_));
 sky130_fd_sc_hd__or3_1 _07384_ (.A(_02556_),
    .B(_02389_),
    .C(\mem[76][7] ),
    .X(_03326_));
 sky130_fd_sc_hd__o221a_1 _07385_ (.A1(\mem[78][7] ),
    .A2(_02554_),
    .B1(_02555_),
    .B2(\mem[79][7] ),
    .C1(_03326_),
    .X(_03327_));
 sky130_fd_sc_hd__o211a_1 _07386_ (.A1(\mem[77][7] ),
    .A2(_02553_),
    .B1(_03327_),
    .C1(_02559_),
    .X(_03328_));
 sky130_fd_sc_hd__o21a_1 _07387_ (.A1(\mem[64][7] ),
    .A2(_02395_),
    .B1(_02563_),
    .X(_03329_));
 sky130_fd_sc_hd__o22a_1 _07388_ (.A1(\mem[65][7] ),
    .A2(_02399_),
    .B1(_02566_),
    .B2(\mem[67][7] ),
    .X(_03330_));
 sky130_fd_sc_hd__o211a_1 _07389_ (.A1(\mem[66][7] ),
    .A2(_02394_),
    .B1(_03329_),
    .C1(_03330_),
    .X(_03331_));
 sky130_fd_sc_hd__or2_1 _07390_ (.A(\mem[72][7] ),
    .B(_02570_),
    .X(_03332_));
 sky130_fd_sc_hd__or3b_1 _07391_ (.A(_02574_),
    .B(\mem[74][7] ),
    .C_N(_02575_),
    .X(_03333_));
 sky130_fd_sc_hd__o221a_1 _07392_ (.A1(\mem[73][7] ),
    .A2(_02572_),
    .B1(_02801_),
    .B2(\mem[75][7] ),
    .C1(_03333_),
    .X(_03334_));
 sky130_fd_sc_hd__o21a_1 _07393_ (.A1(\mem[69][7] ),
    .A2(_02578_),
    .B1(_02463_),
    .X(_03335_));
 sky130_fd_sc_hd__or3_1 _07394_ (.A(_02583_),
    .B(_02868_),
    .C(\mem[68][7] ),
    .X(_03336_));
 sky130_fd_sc_hd__o221a_1 _07395_ (.A1(\mem[70][7] ),
    .A2(_02581_),
    .B1(_02582_),
    .B2(\mem[71][7] ),
    .C1(_03336_),
    .X(_03337_));
 sky130_fd_sc_hd__a32o_1 _07396_ (.A1(_02569_),
    .A2(_03332_),
    .A3(_03334_),
    .B1(_03335_),
    .B2(_03337_),
    .X(_03338_));
 sky130_fd_sc_hd__or4_4 _07397_ (.A(_02552_),
    .B(_03328_),
    .C(_03331_),
    .D(_03338_),
    .X(_03339_));
 sky130_fd_sc_hd__mux4_1 _07398_ (.A0(\mem[96][7] ),
    .A1(\mem[97][7] ),
    .A2(\mem[98][7] ),
    .A3(\mem[99][7] ),
    .S0(_02590_),
    .S1(_02591_),
    .X(_03340_));
 sky130_fd_sc_hd__mux4_1 _07399_ (.A0(\mem[100][7] ),
    .A1(\mem[101][7] ),
    .A2(\mem[102][7] ),
    .A3(\mem[103][7] ),
    .S0(_02593_),
    .S1(_02594_),
    .X(_03341_));
 sky130_fd_sc_hd__a22o_1 _07400_ (.A1(_02651_),
    .A2(_03340_),
    .B1(_03341_),
    .B2(_02825_),
    .X(_03342_));
 sky130_fd_sc_hd__mux4_1 _07401_ (.A0(\mem[108][7] ),
    .A1(\mem[109][7] ),
    .A2(\mem[110][7] ),
    .A3(\mem[111][7] ),
    .S0(_02458_),
    .S1(_02461_),
    .X(_03343_));
 sky130_fd_sc_hd__mux4_1 _07402_ (.A0(\mem[104][7] ),
    .A1(\mem[105][7] ),
    .A2(\mem[106][7] ),
    .A3(\mem[107][7] ),
    .S0(_02501_),
    .S1(_02877_),
    .X(_03344_));
 sky130_fd_sc_hd__or2_1 _07403_ (.A(_02474_),
    .B(_03344_),
    .X(_03345_));
 sky130_fd_sc_hd__o211a_1 _07404_ (.A1(_02598_),
    .A2(_03343_),
    .B1(_03345_),
    .C1(_02478_),
    .X(_03346_));
 sky130_fd_sc_hd__or3_1 _07405_ (.A(_02421_),
    .B(_03342_),
    .C(_03346_),
    .X(_03347_));
 sky130_fd_sc_hd__mux4_1 _07406_ (.A0(\mem[124][7] ),
    .A1(\mem[125][7] ),
    .A2(\mem[126][7] ),
    .A3(\mem[127][7] ),
    .S0(_02613_),
    .S1(_02703_),
    .X(_03348_));
 sky130_fd_sc_hd__mux4_1 _07407_ (.A0(\mem[112][7] ),
    .A1(\mem[113][7] ),
    .A2(\mem[114][7] ),
    .A3(\mem[115][7] ),
    .S0(_02726_),
    .S1(_02618_),
    .X(_03349_));
 sky130_fd_sc_hd__mux4_1 _07408_ (.A0(\mem[116][7] ),
    .A1(\mem[117][7] ),
    .A2(\mem[118][7] ),
    .A3(\mem[119][7] ),
    .S0(_02985_),
    .S1(_02623_),
    .X(_03350_));
 sky130_fd_sc_hd__mux4_1 _07409_ (.A0(\mem[120][7] ),
    .A1(\mem[121][7] ),
    .A2(\mem[122][7] ),
    .A3(\mem[123][7] ),
    .S0(_02887_),
    .S1(_02626_),
    .X(_03351_));
 sky130_fd_sc_hd__o22a_1 _07410_ (.A1(_02885_),
    .A2(_03350_),
    .B1(_03351_),
    .B2(_02889_),
    .X(_03352_));
 sky130_fd_sc_hd__o221a_1 _07411_ (.A1(_02612_),
    .A2(_03348_),
    .B1(_03349_),
    .B2(_02884_),
    .C1(_03352_),
    .X(_03353_));
 sky130_fd_sc_hd__o21a_1 _07412_ (.A1(_02611_),
    .A2(_03353_),
    .B1(_02631_),
    .X(_03354_));
 sky130_fd_sc_hd__a32o_1 _07413_ (.A1(_02513_),
    .A2(_03325_),
    .A3(_03339_),
    .B1(_03347_),
    .B2(_03354_),
    .X(_03355_));
 sky130_fd_sc_hd__mux2_1 _07414_ (.A0(_03311_),
    .A1(_03355_),
    .S(_02635_),
    .X(_03356_));
 sky130_fd_sc_hd__clkbuf_1 _07415_ (.A(_03356_),
    .X(_00013_));
 sky130_fd_sc_hd__o21a_1 _07416_ (.A1(\mem[29][8] ),
    .A2(_02515_),
    .B1(_02366_),
    .X(_03357_));
 sky130_fd_sc_hd__or3_1 _07417_ (.A(_02520_),
    .B(_02779_),
    .C(\mem[28][8] ),
    .X(_03358_));
 sky130_fd_sc_hd__o221a_1 _07418_ (.A1(\mem[30][8] ),
    .A2(_02995_),
    .B1(_02372_),
    .B2(\mem[31][8] ),
    .C1(_03358_),
    .X(_03359_));
 sky130_fd_sc_hd__o21a_1 _07419_ (.A1(\mem[16][8] ),
    .A2(_02380_),
    .B1(_02383_),
    .X(_03360_));
 sky130_fd_sc_hd__or3b_1 _07420_ (.A(_02387_),
    .B(\mem[18][8] ),
    .C_N(_02783_),
    .X(_03361_));
 sky130_fd_sc_hd__o221a_1 _07421_ (.A1(\mem[17][8] ),
    .A2(_02899_),
    .B1(_02528_),
    .B2(\mem[19][8] ),
    .C1(_03361_),
    .X(_03362_));
 sky130_fd_sc_hd__a22o_1 _07422_ (.A1(_03357_),
    .A2(_03359_),
    .B1(_03360_),
    .B2(_03362_),
    .X(_03363_));
 sky130_fd_sc_hd__o21a_1 _07423_ (.A1(\mem[24][8] ),
    .A2(_02788_),
    .B1(_02397_),
    .X(_03364_));
 sky130_fd_sc_hd__o22a_1 _07424_ (.A1(\mem[25][8] ),
    .A2(_02790_),
    .B1(_02401_),
    .B2(\mem[27][8] ),
    .X(_03365_));
 sky130_fd_sc_hd__o211a_1 _07425_ (.A1(\mem[26][8] ),
    .A2(_02787_),
    .B1(_03364_),
    .C1(_03365_),
    .X(_03366_));
 sky130_fd_sc_hd__or3_1 _07426_ (.A(_02793_),
    .B(_02412_),
    .C(\mem[20][8] ),
    .X(_03367_));
 sky130_fd_sc_hd__o221a_1 _07427_ (.A1(\mem[22][8] ),
    .A2(_02543_),
    .B1(_02544_),
    .B2(\mem[23][8] ),
    .C1(_03367_),
    .X(_03368_));
 sky130_fd_sc_hd__o211a_1 _07428_ (.A1(\mem[21][8] ),
    .A2(_02542_),
    .B1(_03368_),
    .C1(_02417_),
    .X(_03369_));
 sky130_fd_sc_hd__or4_2 _07429_ (.A(_02993_),
    .B(_03363_),
    .C(_03366_),
    .D(_03369_),
    .X(_03370_));
 sky130_fd_sc_hd__or3_1 _07430_ (.A(_02432_),
    .B(_02803_),
    .C(\mem[12][8] ),
    .X(_03371_));
 sky130_fd_sc_hd__o221a_1 _07431_ (.A1(\mem[14][8] ),
    .A2(_02800_),
    .B1(_03009_),
    .B2(\mem[15][8] ),
    .C1(_03371_),
    .X(_03372_));
 sky130_fd_sc_hd__o211a_1 _07432_ (.A1(\mem[13][8] ),
    .A2(_02799_),
    .B1(_03372_),
    .C1(_02806_),
    .X(_03373_));
 sky130_fd_sc_hd__o21a_1 _07433_ (.A1(\mem[0][8] ),
    .A2(_02562_),
    .B1(_03013_),
    .X(_03374_));
 sky130_fd_sc_hd__o22a_1 _07434_ (.A1(\mem[1][8] ),
    .A2(_02441_),
    .B1(_02914_),
    .B2(\mem[3][8] ),
    .X(_03375_));
 sky130_fd_sc_hd__o211a_1 _07435_ (.A1(\mem[2][8] ),
    .A2(_02561_),
    .B1(_03374_),
    .C1(_03375_),
    .X(_03376_));
 sky130_fd_sc_hd__or2_1 _07436_ (.A(\mem[8][8] ),
    .B(_02917_),
    .X(_03377_));
 sky130_fd_sc_hd__or3b_1 _07437_ (.A(_02815_),
    .B(\mem[10][8] ),
    .C_N(_02816_),
    .X(_03378_));
 sky130_fd_sc_hd__o221a_1 _07438_ (.A1(\mem[9][8] ),
    .A2(_02736_),
    .B1(_02573_),
    .B2(\mem[11][8] ),
    .C1(_03378_),
    .X(_03379_));
 sky130_fd_sc_hd__o21a_1 _07439_ (.A1(\mem[5][8] ),
    .A2(_02819_),
    .B1(_02579_),
    .X(_03380_));
 sky130_fd_sc_hd__or3_1 _07440_ (.A(_02447_),
    .B(_02584_),
    .C(\mem[4][8] ),
    .X(_03381_));
 sky130_fd_sc_hd__o221a_2 _07441_ (.A1(\mem[6][8] ),
    .A2(_02445_),
    .B1(_02446_),
    .B2(\mem[7][8] ),
    .C1(_03381_),
    .X(_03382_));
 sky130_fd_sc_hd__a32o_2 _07442_ (.A1(_02811_),
    .A2(_03377_),
    .A3(_03379_),
    .B1(_03380_),
    .B2(_03382_),
    .X(_03383_));
 sky130_fd_sc_hd__or4_1 _07443_ (.A(_02798_),
    .B(_03373_),
    .C(_03376_),
    .D(_03383_),
    .X(_03384_));
 sky130_fd_sc_hd__mux4_1 _07444_ (.A0(\mem[32][8] ),
    .A1(\mem[33][8] ),
    .A2(\mem[34][8] ),
    .A3(\mem[35][8] ),
    .S0(_02826_),
    .S1(_02926_),
    .X(_03385_));
 sky130_fd_sc_hd__mux4_1 _07445_ (.A0(\mem[36][8] ),
    .A1(\mem[37][8] ),
    .A2(\mem[38][8] ),
    .A3(\mem[39][8] ),
    .S0(_02928_),
    .S1(_02929_),
    .X(_03386_));
 sky130_fd_sc_hd__a22o_1 _07446_ (.A1(_02456_),
    .A2(_03385_),
    .B1(_03386_),
    .B2(_02465_),
    .X(_03387_));
 sky130_fd_sc_hd__mux4_1 _07447_ (.A0(\mem[44][8] ),
    .A1(\mem[45][8] ),
    .A2(\mem[46][8] ),
    .A3(\mem[47][8] ),
    .S0(_02600_),
    .S1(_02468_),
    .X(_03388_));
 sky130_fd_sc_hd__mux4_1 _07448_ (.A0(\mem[40][8] ),
    .A1(\mem[41][8] ),
    .A2(\mem[42][8] ),
    .A3(\mem[43][8] ),
    .S0(_02604_),
    .S1(_02605_),
    .X(_03389_));
 sky130_fd_sc_hd__or2_1 _07449_ (.A(_02603_),
    .B(_03389_),
    .X(_03390_));
 sky130_fd_sc_hd__o211a_1 _07450_ (.A1(_02472_),
    .A2(_03388_),
    .B1(_03390_),
    .C1(_02608_),
    .X(_03391_));
 sky130_fd_sc_hd__or3_2 _07451_ (.A(_02453_),
    .B(_03387_),
    .C(_03391_),
    .X(_03392_));
 sky130_fd_sc_hd__mux4_1 _07452_ (.A0(\mem[60][8] ),
    .A1(\mem[61][8] ),
    .A2(\mem[62][8] ),
    .A3(\mem[63][8] ),
    .S0(_02487_),
    .S1(_02614_),
    .X(_03393_));
 sky130_fd_sc_hd__mux4_1 _07453_ (.A0(\mem[48][8] ),
    .A1(\mem[49][8] ),
    .A2(\mem[50][8] ),
    .A3(\mem[51][8] ),
    .S0(_02491_),
    .S1(_02746_),
    .X(_03394_));
 sky130_fd_sc_hd__mux4_1 _07454_ (.A0(\mem[52][8] ),
    .A1(\mem[53][8] ),
    .A2(\mem[54][8] ),
    .A3(\mem[55][8] ),
    .S0(_02622_),
    .S1(_02837_),
    .X(_03395_));
 sky130_fd_sc_hd__mux4_1 _07455_ (.A0(\mem[56][8] ),
    .A1(\mem[57][8] ),
    .A2(\mem[58][8] ),
    .A3(\mem[59][8] ),
    .S0(_02625_),
    .S1(_02503_),
    .X(_03396_));
 sky130_fd_sc_hd__o22a_1 _07456_ (.A1(_02621_),
    .A2(_03395_),
    .B1(_03396_),
    .B2(_02628_),
    .X(_03397_));
 sky130_fd_sc_hd__o221a_1 _07457_ (.A1(_03033_),
    .A2(_03393_),
    .B1(_03394_),
    .B2(_02620_),
    .C1(_03397_),
    .X(_03398_));
 sky130_fd_sc_hd__o21a_1 _07458_ (.A1(_02482_),
    .A2(_03398_),
    .B1(_02510_),
    .X(_03399_));
 sky130_fd_sc_hd__a32o_1 _07459_ (.A1(_02356_),
    .A2(_03370_),
    .A3(_03384_),
    .B1(_03392_),
    .B2(_03399_),
    .X(_03400_));
 sky130_fd_sc_hd__o21a_1 _07460_ (.A1(\mem[93][8] ),
    .A2(_03042_),
    .B1(_02516_),
    .X(_03401_));
 sky130_fd_sc_hd__or3_1 _07461_ (.A(_02466_),
    .B(_02521_),
    .C(\mem[92][8] ),
    .X(_03402_));
 sky130_fd_sc_hd__o221a_1 _07462_ (.A1(\mem[94][8] ),
    .A2(_02518_),
    .B1(_02519_),
    .B2(\mem[95][8] ),
    .C1(_03402_),
    .X(_03403_));
 sky130_fd_sc_hd__o21a_1 _07463_ (.A1(\mem[80][8] ),
    .A2(_02812_),
    .B1(_02454_),
    .X(_03404_));
 sky130_fd_sc_hd__or3b_1 _07464_ (.A(_02670_),
    .B(\mem[82][8] ),
    .C_N(_02530_),
    .X(_03405_));
 sky130_fd_sc_hd__o221a_1 _07465_ (.A1(\mem[81][8] ),
    .A2(_02527_),
    .B1(_02424_),
    .B2(\mem[83][8] ),
    .C1(_03405_),
    .X(_03406_));
 sky130_fd_sc_hd__a22o_1 _07466_ (.A1(_03401_),
    .A2(_03403_),
    .B1(_03404_),
    .B2(_03406_),
    .X(_03407_));
 sky130_fd_sc_hd__o21a_1 _07467_ (.A1(\mem[88][8] ),
    .A2(_02535_),
    .B1(_02536_),
    .X(_03408_));
 sky130_fd_sc_hd__o22a_1 _07468_ (.A1(\mem[89][8] ),
    .A2(_02538_),
    .B1(_03231_),
    .B2(\mem[91][8] ),
    .X(_03409_));
 sky130_fd_sc_hd__o211a_1 _07469_ (.A1(\mem[90][8] ),
    .A2(_02534_),
    .B1(_03408_),
    .C1(_03409_),
    .X(_03410_));
 sky130_fd_sc_hd__or3_1 _07470_ (.A(_02545_),
    .B(_02546_),
    .C(\mem[84][8] ),
    .X(_03411_));
 sky130_fd_sc_hd__o221a_1 _07471_ (.A1(\mem[86][8] ),
    .A2(_02956_),
    .B1(_02664_),
    .B2(\mem[87][8] ),
    .C1(_03411_),
    .X(_03412_));
 sky130_fd_sc_hd__o211a_1 _07472_ (.A1(\mem[85][8] ),
    .A2(_02955_),
    .B1(_03412_),
    .C1(_02464_),
    .X(_03413_));
 sky130_fd_sc_hd__or4_4 _07473_ (.A(_02514_),
    .B(_03407_),
    .C(_03410_),
    .D(_03413_),
    .X(_03414_));
 sky130_fd_sc_hd__or3_1 _07474_ (.A(_02556_),
    .B(_02389_),
    .C(\mem[76][8] ),
    .X(_03415_));
 sky130_fd_sc_hd__o221a_1 _07475_ (.A1(\mem[78][8] ),
    .A2(_02554_),
    .B1(_02555_),
    .B2(\mem[79][8] ),
    .C1(_03415_),
    .X(_03416_));
 sky130_fd_sc_hd__o211a_1 _07476_ (.A1(\mem[77][8] ),
    .A2(_02553_),
    .B1(_03416_),
    .C1(_02559_),
    .X(_03417_));
 sky130_fd_sc_hd__o21a_1 _07477_ (.A1(\mem[64][8] ),
    .A2(_02395_),
    .B1(_02563_),
    .X(_03418_));
 sky130_fd_sc_hd__o22a_1 _07478_ (.A1(\mem[65][8] ),
    .A2(_02399_),
    .B1(_02566_),
    .B2(\mem[67][8] ),
    .X(_03419_));
 sky130_fd_sc_hd__o211a_1 _07479_ (.A1(\mem[66][8] ),
    .A2(_02394_),
    .B1(_03418_),
    .C1(_03419_),
    .X(_03420_));
 sky130_fd_sc_hd__or2_1 _07480_ (.A(\mem[72][8] ),
    .B(_02570_),
    .X(_03421_));
 sky130_fd_sc_hd__or3b_1 _07481_ (.A(_02574_),
    .B(\mem[74][8] ),
    .C_N(_02575_),
    .X(_03422_));
 sky130_fd_sc_hd__o221a_1 _07482_ (.A1(\mem[73][8] ),
    .A2(_02385_),
    .B1(_02801_),
    .B2(\mem[75][8] ),
    .C1(_03422_),
    .X(_03423_));
 sky130_fd_sc_hd__o21a_1 _07483_ (.A1(\mem[69][8] ),
    .A2(_02578_),
    .B1(_02463_),
    .X(_03424_));
 sky130_fd_sc_hd__or3_1 _07484_ (.A(_02411_),
    .B(_02868_),
    .C(\mem[68][8] ),
    .X(_03425_));
 sky130_fd_sc_hd__o221a_1 _07485_ (.A1(\mem[70][8] ),
    .A2(_02581_),
    .B1(_02582_),
    .B2(\mem[71][8] ),
    .C1(_03425_),
    .X(_03426_));
 sky130_fd_sc_hd__a32o_1 _07486_ (.A1(_02569_),
    .A2(_03421_),
    .A3(_03423_),
    .B1(_03424_),
    .B2(_03426_),
    .X(_03427_));
 sky130_fd_sc_hd__or4_4 _07487_ (.A(_02552_),
    .B(_03417_),
    .C(_03420_),
    .D(_03427_),
    .X(_03428_));
 sky130_fd_sc_hd__mux4_1 _07488_ (.A0(\mem[96][8] ),
    .A1(\mem[97][8] ),
    .A2(\mem[98][8] ),
    .A3(\mem[99][8] ),
    .S0(_02590_),
    .S1(_02591_),
    .X(_03429_));
 sky130_fd_sc_hd__mux4_1 _07489_ (.A0(\mem[100][8] ),
    .A1(\mem[101][8] ),
    .A2(\mem[102][8] ),
    .A3(\mem[103][8] ),
    .S0(_02593_),
    .S1(_02594_),
    .X(_03430_));
 sky130_fd_sc_hd__a22o_1 _07490_ (.A1(_02651_),
    .A2(_03429_),
    .B1(_03430_),
    .B2(_02825_),
    .X(_03431_));
 sky130_fd_sc_hd__mux4_1 _07491_ (.A0(\mem[108][8] ),
    .A1(\mem[109][8] ),
    .A2(\mem[110][8] ),
    .A3(\mem[111][8] ),
    .S0(_02458_),
    .S1(_02461_),
    .X(_03432_));
 sky130_fd_sc_hd__mux4_1 _07492_ (.A0(\mem[104][8] ),
    .A1(\mem[105][8] ),
    .A2(\mem[106][8] ),
    .A3(\mem[107][8] ),
    .S0(_02501_),
    .S1(_02877_),
    .X(_03433_));
 sky130_fd_sc_hd__or2_1 _07493_ (.A(_02474_),
    .B(_03433_),
    .X(_03434_));
 sky130_fd_sc_hd__o211a_1 _07494_ (.A1(_02598_),
    .A2(_03432_),
    .B1(_03434_),
    .C1(_02478_),
    .X(_03435_));
 sky130_fd_sc_hd__or3_1 _07495_ (.A(_02421_),
    .B(_03431_),
    .C(_03435_),
    .X(_03436_));
 sky130_fd_sc_hd__mux4_1 _07496_ (.A0(\mem[124][8] ),
    .A1(\mem[125][8] ),
    .A2(\mem[126][8] ),
    .A3(\mem[127][8] ),
    .S0(_02613_),
    .S1(_02703_),
    .X(_03437_));
 sky130_fd_sc_hd__mux4_1 _07497_ (.A0(\mem[112][8] ),
    .A1(\mem[113][8] ),
    .A2(\mem[114][8] ),
    .A3(\mem[115][8] ),
    .S0(_02726_),
    .S1(_02618_),
    .X(_03438_));
 sky130_fd_sc_hd__mux4_1 _07498_ (.A0(\mem[116][8] ),
    .A1(\mem[117][8] ),
    .A2(\mem[118][8] ),
    .A3(\mem[119][8] ),
    .S0(_02985_),
    .S1(_02623_),
    .X(_03439_));
 sky130_fd_sc_hd__mux4_1 _07499_ (.A0(\mem[120][8] ),
    .A1(\mem[121][8] ),
    .A2(\mem[122][8] ),
    .A3(\mem[123][8] ),
    .S0(_02887_),
    .S1(_02499_),
    .X(_03440_));
 sky130_fd_sc_hd__o22a_1 _07500_ (.A1(_02885_),
    .A2(_03439_),
    .B1(_03440_),
    .B2(_02889_),
    .X(_03441_));
 sky130_fd_sc_hd__o221a_1 _07501_ (.A1(_02612_),
    .A2(_03437_),
    .B1(_03438_),
    .B2(_02884_),
    .C1(_03441_),
    .X(_03442_));
 sky130_fd_sc_hd__o21a_1 _07502_ (.A1(_02611_),
    .A2(_03442_),
    .B1(_02509_),
    .X(_03443_));
 sky130_fd_sc_hd__a32o_1 _07503_ (.A1(_02355_),
    .A2(_03414_),
    .A3(_03428_),
    .B1(_03436_),
    .B2(_03443_),
    .X(_03444_));
 sky130_fd_sc_hd__mux2_1 _07504_ (.A0(_03400_),
    .A1(_03444_),
    .S(_02635_),
    .X(_03445_));
 sky130_fd_sc_hd__clkbuf_1 _07505_ (.A(_03445_),
    .X(_00014_));
 sky130_fd_sc_hd__o21a_1 _07506_ (.A1(\mem[29][9] ),
    .A2(_02515_),
    .B1(_02366_),
    .X(_03446_));
 sky130_fd_sc_hd__or3_1 _07507_ (.A(_02520_),
    .B(_02779_),
    .C(\mem[28][9] ),
    .X(_03447_));
 sky130_fd_sc_hd__o221a_1 _07508_ (.A1(\mem[30][9] ),
    .A2(_02995_),
    .B1(_02372_),
    .B2(\mem[31][9] ),
    .C1(_03447_),
    .X(_03448_));
 sky130_fd_sc_hd__o21a_1 _07509_ (.A1(\mem[16][9] ),
    .A2(_02524_),
    .B1(_02383_),
    .X(_03449_));
 sky130_fd_sc_hd__or3b_1 _07510_ (.A(_02529_),
    .B(\mem[18][9] ),
    .C_N(_02783_),
    .X(_03450_));
 sky130_fd_sc_hd__o221a_1 _07511_ (.A1(\mem[17][9] ),
    .A2(_02899_),
    .B1(_02528_),
    .B2(\mem[19][9] ),
    .C1(_03450_),
    .X(_03451_));
 sky130_fd_sc_hd__a22o_1 _07512_ (.A1(_03446_),
    .A2(_03448_),
    .B1(_03449_),
    .B2(_03451_),
    .X(_03452_));
 sky130_fd_sc_hd__o21a_1 _07513_ (.A1(\mem[24][9] ),
    .A2(_02788_),
    .B1(_02397_),
    .X(_03453_));
 sky130_fd_sc_hd__o22a_1 _07514_ (.A1(\mem[25][9] ),
    .A2(_02790_),
    .B1(_02401_),
    .B2(\mem[27][9] ),
    .X(_03454_));
 sky130_fd_sc_hd__o211a_1 _07515_ (.A1(\mem[26][9] ),
    .A2(_02787_),
    .B1(_03453_),
    .C1(_03454_),
    .X(_03455_));
 sky130_fd_sc_hd__or3_1 _07516_ (.A(_02793_),
    .B(_02412_),
    .C(\mem[20][9] ),
    .X(_03456_));
 sky130_fd_sc_hd__o221a_1 _07517_ (.A1(\mem[22][9] ),
    .A2(_02543_),
    .B1(_02544_),
    .B2(\mem[23][9] ),
    .C1(_03456_),
    .X(_03457_));
 sky130_fd_sc_hd__o211a_1 _07518_ (.A1(\mem[21][9] ),
    .A2(_02542_),
    .B1(_03457_),
    .C1(_02549_),
    .X(_03458_));
 sky130_fd_sc_hd__or4_2 _07519_ (.A(_02993_),
    .B(_03452_),
    .C(_03455_),
    .D(_03458_),
    .X(_03459_));
 sky130_fd_sc_hd__or3_1 _07520_ (.A(_02432_),
    .B(_02803_),
    .C(\mem[12][9] ),
    .X(_03460_));
 sky130_fd_sc_hd__o221a_1 _07521_ (.A1(\mem[14][9] ),
    .A2(_02800_),
    .B1(_03009_),
    .B2(\mem[15][9] ),
    .C1(_03460_),
    .X(_03461_));
 sky130_fd_sc_hd__o211a_1 _07522_ (.A1(\mem[13][9] ),
    .A2(_02799_),
    .B1(_03461_),
    .C1(_02806_),
    .X(_03462_));
 sky130_fd_sc_hd__o21a_1 _07523_ (.A1(\mem[0][9] ),
    .A2(_02562_),
    .B1(_03013_),
    .X(_03463_));
 sky130_fd_sc_hd__o22a_1 _07524_ (.A1(\mem[1][9] ),
    .A2(_02441_),
    .B1(_02914_),
    .B2(\mem[3][9] ),
    .X(_03464_));
 sky130_fd_sc_hd__o211a_1 _07525_ (.A1(\mem[2][9] ),
    .A2(_02561_),
    .B1(_03463_),
    .C1(_03464_),
    .X(_03465_));
 sky130_fd_sc_hd__or2_1 _07526_ (.A(\mem[8][9] ),
    .B(_02917_),
    .X(_03466_));
 sky130_fd_sc_hd__or3b_1 _07527_ (.A(_02815_),
    .B(\mem[10][9] ),
    .C_N(_02816_),
    .X(_03467_));
 sky130_fd_sc_hd__o221a_1 _07528_ (.A1(\mem[9][9] ),
    .A2(_02736_),
    .B1(_02573_),
    .B2(\mem[11][9] ),
    .C1(_03467_),
    .X(_03468_));
 sky130_fd_sc_hd__o21a_1 _07529_ (.A1(\mem[5][9] ),
    .A2(_02819_),
    .B1(_02579_),
    .X(_03469_));
 sky130_fd_sc_hd__or3_1 _07530_ (.A(_02447_),
    .B(_02584_),
    .C(\mem[4][9] ),
    .X(_03470_));
 sky130_fd_sc_hd__o221a_1 _07531_ (.A1(\mem[6][9] ),
    .A2(_02445_),
    .B1(_02446_),
    .B2(\mem[7][9] ),
    .C1(_03470_),
    .X(_03471_));
 sky130_fd_sc_hd__a32o_2 _07532_ (.A1(_02811_),
    .A2(_03466_),
    .A3(_03468_),
    .B1(_03469_),
    .B2(_03471_),
    .X(_03472_));
 sky130_fd_sc_hd__or4_1 _07533_ (.A(_02798_),
    .B(_03462_),
    .C(_03465_),
    .D(_03472_),
    .X(_03473_));
 sky130_fd_sc_hd__mux4_1 _07534_ (.A0(\mem[32][9] ),
    .A1(\mem[33][9] ),
    .A2(\mem[34][9] ),
    .A3(\mem[35][9] ),
    .S0(_02826_),
    .S1(_02926_),
    .X(_03474_));
 sky130_fd_sc_hd__mux4_1 _07535_ (.A0(\mem[36][9] ),
    .A1(\mem[37][9] ),
    .A2(\mem[38][9] ),
    .A3(\mem[39][9] ),
    .S0(_02928_),
    .S1(_02929_),
    .X(_03475_));
 sky130_fd_sc_hd__a22o_1 _07536_ (.A1(_02456_),
    .A2(_03474_),
    .B1(_03475_),
    .B2(_02465_),
    .X(_03476_));
 sky130_fd_sc_hd__mux4_1 _07537_ (.A0(\mem[44][9] ),
    .A1(\mem[45][9] ),
    .A2(\mem[46][9] ),
    .A3(\mem[47][9] ),
    .S0(_02600_),
    .S1(_02601_),
    .X(_03477_));
 sky130_fd_sc_hd__mux4_1 _07538_ (.A0(\mem[40][9] ),
    .A1(\mem[41][9] ),
    .A2(\mem[42][9] ),
    .A3(\mem[43][9] ),
    .S0(_02604_),
    .S1(_02605_),
    .X(_03478_));
 sky130_fd_sc_hd__or2_1 _07539_ (.A(_02603_),
    .B(_03478_),
    .X(_03479_));
 sky130_fd_sc_hd__o211a_1 _07540_ (.A1(_02599_),
    .A2(_03477_),
    .B1(_03479_),
    .C1(_02608_),
    .X(_03480_));
 sky130_fd_sc_hd__or3_2 _07541_ (.A(_02589_),
    .B(_03476_),
    .C(_03480_),
    .X(_03481_));
 sky130_fd_sc_hd__mux4_1 _07542_ (.A0(\mem[60][9] ),
    .A1(\mem[61][9] ),
    .A2(\mem[62][9] ),
    .A3(\mem[63][9] ),
    .S0(_02487_),
    .S1(_02614_),
    .X(_03482_));
 sky130_fd_sc_hd__mux4_1 _07543_ (.A0(\mem[48][9] ),
    .A1(\mem[49][9] ),
    .A2(\mem[50][9] ),
    .A3(\mem[51][9] ),
    .S0(_02616_),
    .S1(_02746_),
    .X(_03483_));
 sky130_fd_sc_hd__mux4_1 _07544_ (.A0(\mem[52][9] ),
    .A1(\mem[53][9] ),
    .A2(\mem[54][9] ),
    .A3(\mem[55][9] ),
    .S0(_02622_),
    .S1(_02837_),
    .X(_03484_));
 sky130_fd_sc_hd__mux4_1 _07545_ (.A0(\mem[56][9] ),
    .A1(\mem[57][9] ),
    .A2(\mem[58][9] ),
    .A3(\mem[59][9] ),
    .S0(_02625_),
    .S1(_02503_),
    .X(_03485_));
 sky130_fd_sc_hd__o22a_1 _07546_ (.A1(_02621_),
    .A2(_03484_),
    .B1(_03485_),
    .B2(_02628_),
    .X(_03486_));
 sky130_fd_sc_hd__o221a_1 _07547_ (.A1(_03033_),
    .A2(_03482_),
    .B1(_03483_),
    .B2(_02620_),
    .C1(_03486_),
    .X(_03487_));
 sky130_fd_sc_hd__o21a_1 _07548_ (.A1(_02482_),
    .A2(_03487_),
    .B1(_02510_),
    .X(_03488_));
 sky130_fd_sc_hd__a32o_1 _07549_ (.A1(_02356_),
    .A2(_03459_),
    .A3(_03473_),
    .B1(_03481_),
    .B2(_03488_),
    .X(_03489_));
 sky130_fd_sc_hd__o21a_1 _07550_ (.A1(\mem[93][9] ),
    .A2(_03042_),
    .B1(_02365_),
    .X(_03490_));
 sky130_fd_sc_hd__or3_1 _07551_ (.A(_02466_),
    .B(_02521_),
    .C(\mem[92][9] ),
    .X(_03491_));
 sky130_fd_sc_hd__o221a_1 _07552_ (.A1(\mem[94][9] ),
    .A2(_02518_),
    .B1(_02519_),
    .B2(\mem[95][9] ),
    .C1(_03491_),
    .X(_03492_));
 sky130_fd_sc_hd__o21a_1 _07553_ (.A1(\mem[80][9] ),
    .A2(_02812_),
    .B1(_02454_),
    .X(_03493_));
 sky130_fd_sc_hd__or3b_1 _07554_ (.A(_02670_),
    .B(\mem[82][9] ),
    .C_N(_02530_),
    .X(_03494_));
 sky130_fd_sc_hd__o221a_1 _07555_ (.A1(\mem[81][9] ),
    .A2(_02527_),
    .B1(_02424_),
    .B2(\mem[83][9] ),
    .C1(_03494_),
    .X(_03495_));
 sky130_fd_sc_hd__a22o_1 _07556_ (.A1(_03490_),
    .A2(_03492_),
    .B1(_03493_),
    .B2(_03495_),
    .X(_03496_));
 sky130_fd_sc_hd__o21a_1 _07557_ (.A1(\mem[88][9] ),
    .A2(_02535_),
    .B1(_02536_),
    .X(_03497_));
 sky130_fd_sc_hd__o22a_1 _07558_ (.A1(\mem[89][9] ),
    .A2(_02538_),
    .B1(_03231_),
    .B2(\mem[91][9] ),
    .X(_03498_));
 sky130_fd_sc_hd__o211a_1 _07559_ (.A1(\mem[90][9] ),
    .A2(_02534_),
    .B1(_03497_),
    .C1(_03498_),
    .X(_03499_));
 sky130_fd_sc_hd__or3_1 _07560_ (.A(_02545_),
    .B(_02546_),
    .C(\mem[84][9] ),
    .X(_03500_));
 sky130_fd_sc_hd__o221a_1 _07561_ (.A1(\mem[86][9] ),
    .A2(_02956_),
    .B1(_02664_),
    .B2(\mem[87][9] ),
    .C1(_03500_),
    .X(_03501_));
 sky130_fd_sc_hd__o211a_1 _07562_ (.A1(\mem[85][9] ),
    .A2(_02955_),
    .B1(_03501_),
    .C1(_02464_),
    .X(_03502_));
 sky130_fd_sc_hd__or4_4 _07563_ (.A(_02514_),
    .B(_03496_),
    .C(_03499_),
    .D(_03502_),
    .X(_03503_));
 sky130_fd_sc_hd__or3_1 _07564_ (.A(_02556_),
    .B(_02389_),
    .C(\mem[76][9] ),
    .X(_03504_));
 sky130_fd_sc_hd__o221a_1 _07565_ (.A1(\mem[78][9] ),
    .A2(_02554_),
    .B1(_02555_),
    .B2(\mem[79][9] ),
    .C1(_03504_),
    .X(_03505_));
 sky130_fd_sc_hd__o211a_1 _07566_ (.A1(\mem[77][9] ),
    .A2(_02553_),
    .B1(_03505_),
    .C1(_02559_),
    .X(_03506_));
 sky130_fd_sc_hd__o21a_1 _07567_ (.A1(\mem[64][9] ),
    .A2(_02395_),
    .B1(_02563_),
    .X(_03507_));
 sky130_fd_sc_hd__o22a_1 _07568_ (.A1(\mem[65][9] ),
    .A2(_02399_),
    .B1(_02566_),
    .B2(\mem[67][9] ),
    .X(_03508_));
 sky130_fd_sc_hd__o211a_1 _07569_ (.A1(\mem[66][9] ),
    .A2(_02394_),
    .B1(_03507_),
    .C1(_03508_),
    .X(_03509_));
 sky130_fd_sc_hd__or2_1 _07570_ (.A(\mem[72][9] ),
    .B(_02570_),
    .X(_03510_));
 sky130_fd_sc_hd__or3b_1 _07571_ (.A(_02802_),
    .B(\mem[74][9] ),
    .C_N(_02575_),
    .X(_03511_));
 sky130_fd_sc_hd__o221a_1 _07572_ (.A1(\mem[73][9] ),
    .A2(_02385_),
    .B1(_02801_),
    .B2(\mem[75][9] ),
    .C1(_03511_),
    .X(_03512_));
 sky130_fd_sc_hd__o21a_1 _07573_ (.A1(\mem[69][9] ),
    .A2(_02405_),
    .B1(_02463_),
    .X(_03513_));
 sky130_fd_sc_hd__or3_1 _07574_ (.A(_02411_),
    .B(_02868_),
    .C(\mem[68][9] ),
    .X(_03514_));
 sky130_fd_sc_hd__o221a_1 _07575_ (.A1(\mem[70][9] ),
    .A2(_02407_),
    .B1(_02582_),
    .B2(\mem[71][9] ),
    .C1(_03514_),
    .X(_03515_));
 sky130_fd_sc_hd__a32o_1 _07576_ (.A1(_02569_),
    .A2(_03510_),
    .A3(_03512_),
    .B1(_03513_),
    .B2(_03515_),
    .X(_03516_));
 sky130_fd_sc_hd__or4_2 _07577_ (.A(_02552_),
    .B(_03506_),
    .C(_03509_),
    .D(_03516_),
    .X(_03517_));
 sky130_fd_sc_hd__mux4_1 _07578_ (.A0(\mem[96][9] ),
    .A1(\mem[97][9] ),
    .A2(\mem[98][9] ),
    .A3(\mem[99][9] ),
    .S0(_02590_),
    .S1(_02591_),
    .X(_03518_));
 sky130_fd_sc_hd__mux4_1 _07579_ (.A0(\mem[100][9] ),
    .A1(\mem[101][9] ),
    .A2(\mem[102][9] ),
    .A3(\mem[103][9] ),
    .S0(_02593_),
    .S1(_02594_),
    .X(_03519_));
 sky130_fd_sc_hd__a22o_1 _07580_ (.A1(_02651_),
    .A2(_03518_),
    .B1(_03519_),
    .B2(_02825_),
    .X(_03520_));
 sky130_fd_sc_hd__mux4_2 _07581_ (.A0(\mem[108][9] ),
    .A1(\mem[109][9] ),
    .A2(\mem[110][9] ),
    .A3(\mem[111][9] ),
    .S0(_02458_),
    .S1(_02461_),
    .X(_03521_));
 sky130_fd_sc_hd__mux4_1 _07582_ (.A0(\mem[104][9] ),
    .A1(\mem[105][9] ),
    .A2(\mem[106][9] ),
    .A3(\mem[107][9] ),
    .S0(_02501_),
    .S1(_02877_),
    .X(_03522_));
 sky130_fd_sc_hd__or2_1 _07583_ (.A(_02474_),
    .B(_03522_),
    .X(_03523_));
 sky130_fd_sc_hd__o211a_1 _07584_ (.A1(_02598_),
    .A2(_03521_),
    .B1(_03523_),
    .C1(_02478_),
    .X(_03524_));
 sky130_fd_sc_hd__or3_2 _07585_ (.A(_02421_),
    .B(_03520_),
    .C(_03524_),
    .X(_03525_));
 sky130_fd_sc_hd__mux4_1 _07586_ (.A0(\mem[124][9] ),
    .A1(\mem[125][9] ),
    .A2(\mem[126][9] ),
    .A3(\mem[127][9] ),
    .S0(_02671_),
    .S1(_02703_),
    .X(_03526_));
 sky130_fd_sc_hd__mux4_1 _07587_ (.A0(\mem[112][9] ),
    .A1(\mem[113][9] ),
    .A2(\mem[114][9] ),
    .A3(\mem[115][9] ),
    .S0(_02726_),
    .S1(_02618_),
    .X(_03527_));
 sky130_fd_sc_hd__mux4_1 _07588_ (.A0(\mem[116][9] ),
    .A1(\mem[117][9] ),
    .A2(\mem[118][9] ),
    .A3(\mem[119][9] ),
    .S0(_02985_),
    .S1(_02623_),
    .X(_03528_));
 sky130_fd_sc_hd__mux4_1 _07589_ (.A0(\mem[120][9] ),
    .A1(\mem[121][9] ),
    .A2(\mem[122][9] ),
    .A3(\mem[123][9] ),
    .S0(_02887_),
    .S1(_02499_),
    .X(_03529_));
 sky130_fd_sc_hd__o22a_1 _07590_ (.A1(_02885_),
    .A2(_03528_),
    .B1(_03529_),
    .B2(_02889_),
    .X(_03530_));
 sky130_fd_sc_hd__o221a_2 _07591_ (.A1(_02612_),
    .A2(_03526_),
    .B1(_03527_),
    .B2(_02884_),
    .C1(_03530_),
    .X(_03531_));
 sky130_fd_sc_hd__o21a_1 _07592_ (.A1(_02358_),
    .A2(_03531_),
    .B1(_02509_),
    .X(_03532_));
 sky130_fd_sc_hd__a32o_1 _07593_ (.A1(_02355_),
    .A2(_03503_),
    .A3(_03517_),
    .B1(_03525_),
    .B2(_03532_),
    .X(_03533_));
 sky130_fd_sc_hd__mux2_1 _07594_ (.A0(_03489_),
    .A1(_03533_),
    .S(_02634_),
    .X(_03534_));
 sky130_fd_sc_hd__clkbuf_1 _07595_ (.A(_03534_),
    .X(_00015_));
 sky130_fd_sc_hd__o21a_1 _07596_ (.A1(\mem[29][10] ),
    .A2(_02515_),
    .B1(_02366_),
    .X(_03535_));
 sky130_fd_sc_hd__or3_1 _07597_ (.A(_02520_),
    .B(_02779_),
    .C(\mem[28][10] ),
    .X(_03536_));
 sky130_fd_sc_hd__o221a_1 _07598_ (.A1(\mem[30][10] ),
    .A2(_02995_),
    .B1(_02372_),
    .B2(\mem[31][10] ),
    .C1(_03536_),
    .X(_03537_));
 sky130_fd_sc_hd__o21a_1 _07599_ (.A1(\mem[16][10] ),
    .A2(_02524_),
    .B1(_02525_),
    .X(_03538_));
 sky130_fd_sc_hd__or3b_1 _07600_ (.A(_02529_),
    .B(\mem[18][10] ),
    .C_N(_02783_),
    .X(_03539_));
 sky130_fd_sc_hd__o221a_1 _07601_ (.A1(\mem[17][10] ),
    .A2(_02899_),
    .B1(_02528_),
    .B2(\mem[19][10] ),
    .C1(_03539_),
    .X(_03540_));
 sky130_fd_sc_hd__a22o_1 _07602_ (.A1(_03535_),
    .A2(_03537_),
    .B1(_03538_),
    .B2(_03540_),
    .X(_03541_));
 sky130_fd_sc_hd__o21a_1 _07603_ (.A1(\mem[24][10] ),
    .A2(_02788_),
    .B1(_02397_),
    .X(_03542_));
 sky130_fd_sc_hd__o22a_1 _07604_ (.A1(\mem[25][10] ),
    .A2(_02790_),
    .B1(_02539_),
    .B2(\mem[27][10] ),
    .X(_03543_));
 sky130_fd_sc_hd__o211a_1 _07605_ (.A1(\mem[26][10] ),
    .A2(_02787_),
    .B1(_03542_),
    .C1(_03543_),
    .X(_03544_));
 sky130_fd_sc_hd__or3_1 _07606_ (.A(_02793_),
    .B(_02412_),
    .C(\mem[20][10] ),
    .X(_03545_));
 sky130_fd_sc_hd__o221a_1 _07607_ (.A1(\mem[22][10] ),
    .A2(_02543_),
    .B1(_02544_),
    .B2(\mem[23][10] ),
    .C1(_03545_),
    .X(_03546_));
 sky130_fd_sc_hd__o211a_1 _07608_ (.A1(\mem[21][10] ),
    .A2(_02542_),
    .B1(_03546_),
    .C1(_02549_),
    .X(_03547_));
 sky130_fd_sc_hd__or4_4 _07609_ (.A(_02993_),
    .B(_03541_),
    .C(_03544_),
    .D(_03547_),
    .X(_03548_));
 sky130_fd_sc_hd__or3_1 _07610_ (.A(_02432_),
    .B(_02433_),
    .C(\mem[12][10] ),
    .X(_03549_));
 sky130_fd_sc_hd__o221a_1 _07611_ (.A1(\mem[14][10] ),
    .A2(_02800_),
    .B1(_03009_),
    .B2(\mem[15][10] ),
    .C1(_03549_),
    .X(_03550_));
 sky130_fd_sc_hd__o211a_1 _07612_ (.A1(\mem[13][10] ),
    .A2(_02799_),
    .B1(_03550_),
    .C1(_02806_),
    .X(_03551_));
 sky130_fd_sc_hd__o21a_1 _07613_ (.A1(\mem[0][10] ),
    .A2(_02562_),
    .B1(_03013_),
    .X(_03552_));
 sky130_fd_sc_hd__o22a_1 _07614_ (.A1(\mem[1][10] ),
    .A2(_02565_),
    .B1(_02914_),
    .B2(\mem[3][10] ),
    .X(_03553_));
 sky130_fd_sc_hd__o211a_1 _07615_ (.A1(\mem[2][10] ),
    .A2(_02561_),
    .B1(_03552_),
    .C1(_03553_),
    .X(_03554_));
 sky130_fd_sc_hd__or2_1 _07616_ (.A(\mem[8][10] ),
    .B(_02917_),
    .X(_03555_));
 sky130_fd_sc_hd__or3b_1 _07617_ (.A(_02815_),
    .B(\mem[10][10] ),
    .C_N(_02816_),
    .X(_03556_));
 sky130_fd_sc_hd__o221a_1 _07618_ (.A1(\mem[9][10] ),
    .A2(_02572_),
    .B1(_02573_),
    .B2(\mem[11][10] ),
    .C1(_03556_),
    .X(_03557_));
 sky130_fd_sc_hd__o21a_1 _07619_ (.A1(\mem[5][10] ),
    .A2(_02819_),
    .B1(_02579_),
    .X(_03558_));
 sky130_fd_sc_hd__or3_1 _07620_ (.A(_02583_),
    .B(_02584_),
    .C(\mem[4][10] ),
    .X(_03559_));
 sky130_fd_sc_hd__o221a_1 _07621_ (.A1(\mem[6][10] ),
    .A2(_02445_),
    .B1(_02446_),
    .B2(\mem[7][10] ),
    .C1(_03559_),
    .X(_03560_));
 sky130_fd_sc_hd__a32o_1 _07622_ (.A1(_02811_),
    .A2(_03555_),
    .A3(_03557_),
    .B1(_03558_),
    .B2(_03560_),
    .X(_03561_));
 sky130_fd_sc_hd__or4_1 _07623_ (.A(_02798_),
    .B(_03551_),
    .C(_03554_),
    .D(_03561_),
    .X(_03562_));
 sky130_fd_sc_hd__mux4_1 _07624_ (.A0(\mem[36][10] ),
    .A1(\mem[37][10] ),
    .A2(\mem[38][10] ),
    .A3(\mem[39][10] ),
    .S0(_02826_),
    .S1(_02926_),
    .X(_03563_));
 sky130_fd_sc_hd__mux4_1 _07625_ (.A0(\mem[32][10] ),
    .A1(\mem[33][10] ),
    .A2(\mem[34][10] ),
    .A3(\mem[35][10] ),
    .S0(_02928_),
    .S1(_02929_),
    .X(_03564_));
 sky130_fd_sc_hd__a22o_1 _07626_ (.A1(_02450_),
    .A2(_03563_),
    .B1(_03564_),
    .B2(_02596_),
    .X(_03565_));
 sky130_fd_sc_hd__mux4_1 _07627_ (.A0(\mem[44][10] ),
    .A1(\mem[45][10] ),
    .A2(\mem[46][10] ),
    .A3(\mem[47][10] ),
    .S0(_02600_),
    .S1(_02601_),
    .X(_03566_));
 sky130_fd_sc_hd__mux4_1 _07628_ (.A0(\mem[40][10] ),
    .A1(\mem[41][10] ),
    .A2(\mem[42][10] ),
    .A3(\mem[43][10] ),
    .S0(_02604_),
    .S1(_02605_),
    .X(_03567_));
 sky130_fd_sc_hd__or2_1 _07629_ (.A(_02603_),
    .B(_03567_),
    .X(_03568_));
 sky130_fd_sc_hd__o211a_1 _07630_ (.A1(_02599_),
    .A2(_03566_),
    .B1(_03568_),
    .C1(_02608_),
    .X(_03569_));
 sky130_fd_sc_hd__or3_2 _07631_ (.A(_02589_),
    .B(_03565_),
    .C(_03569_),
    .X(_03570_));
 sky130_fd_sc_hd__mux4_1 _07632_ (.A0(\mem[60][10] ),
    .A1(\mem[61][10] ),
    .A2(\mem[62][10] ),
    .A3(\mem[63][10] ),
    .S0(_02487_),
    .S1(_02614_),
    .X(_03571_));
 sky130_fd_sc_hd__mux4_1 _07633_ (.A0(\mem[48][10] ),
    .A1(\mem[49][10] ),
    .A2(\mem[50][10] ),
    .A3(\mem[51][10] ),
    .S0(_02616_),
    .S1(_02746_),
    .X(_03572_));
 sky130_fd_sc_hd__mux4_1 _07634_ (.A0(\mem[52][10] ),
    .A1(\mem[53][10] ),
    .A2(\mem[54][10] ),
    .A3(\mem[55][10] ),
    .S0(_02622_),
    .S1(_02837_),
    .X(_03573_));
 sky130_fd_sc_hd__mux4_1 _07635_ (.A0(\mem[56][10] ),
    .A1(\mem[57][10] ),
    .A2(\mem[58][10] ),
    .A3(\mem[59][10] ),
    .S0(_02625_),
    .S1(_02626_),
    .X(_03574_));
 sky130_fd_sc_hd__o22a_1 _07636_ (.A1(_02621_),
    .A2(_03573_),
    .B1(_03574_),
    .B2(_02628_),
    .X(_03575_));
 sky130_fd_sc_hd__o221a_1 _07637_ (.A1(_03033_),
    .A2(_03571_),
    .B1(_03572_),
    .B2(_02620_),
    .C1(_03575_),
    .X(_03576_));
 sky130_fd_sc_hd__o21a_1 _07638_ (.A1(_02482_),
    .A2(_03576_),
    .B1(_02631_),
    .X(_03577_));
 sky130_fd_sc_hd__a32o_1 _07639_ (.A1(_02513_),
    .A2(_03548_),
    .A3(_03562_),
    .B1(_03570_),
    .B2(_03577_),
    .X(_03578_));
 sky130_fd_sc_hd__o21a_1 _07640_ (.A1(\mem[93][10] ),
    .A2(_03042_),
    .B1(_02365_),
    .X(_03579_));
 sky130_fd_sc_hd__or3_1 _07641_ (.A(_02466_),
    .B(_02459_),
    .C(\mem[92][10] ),
    .X(_03580_));
 sky130_fd_sc_hd__o221a_1 _07642_ (.A1(\mem[94][10] ),
    .A2(_02518_),
    .B1(_02400_),
    .B2(\mem[95][10] ),
    .C1(_03580_),
    .X(_03581_));
 sky130_fd_sc_hd__o21a_1 _07643_ (.A1(\mem[80][10] ),
    .A2(_02812_),
    .B1(_02454_),
    .X(_03582_));
 sky130_fd_sc_hd__or3b_1 _07644_ (.A(_02670_),
    .B(\mem[82][10] ),
    .C_N(_02530_),
    .X(_03583_));
 sky130_fd_sc_hd__o221a_1 _07645_ (.A1(\mem[81][10] ),
    .A2(_02527_),
    .B1(_02424_),
    .B2(\mem[83][10] ),
    .C1(_03583_),
    .X(_03584_));
 sky130_fd_sc_hd__a22o_1 _07646_ (.A1(_03579_),
    .A2(_03581_),
    .B1(_03582_),
    .B2(_03584_),
    .X(_03585_));
 sky130_fd_sc_hd__o21a_1 _07647_ (.A1(\mem[88][10] ),
    .A2(_02535_),
    .B1(_02396_),
    .X(_03586_));
 sky130_fd_sc_hd__o22a_1 _07648_ (.A1(\mem[89][10] ),
    .A2(_02363_),
    .B1(_03231_),
    .B2(\mem[91][10] ),
    .X(_03587_));
 sky130_fd_sc_hd__o211a_1 _07649_ (.A1(\mem[90][10] ),
    .A2(_02534_),
    .B1(_03586_),
    .C1(_03587_),
    .X(_03588_));
 sky130_fd_sc_hd__or3_1 _07650_ (.A(_02486_),
    .B(_03224_),
    .C(\mem[84][10] ),
    .X(_03589_));
 sky130_fd_sc_hd__o221a_1 _07651_ (.A1(\mem[86][10] ),
    .A2(_02956_),
    .B1(_02664_),
    .B2(\mem[87][10] ),
    .C1(_03589_),
    .X(_03590_));
 sky130_fd_sc_hd__o211a_1 _07652_ (.A1(\mem[85][10] ),
    .A2(_02955_),
    .B1(_03590_),
    .C1(_02464_),
    .X(_03591_));
 sky130_fd_sc_hd__or4_2 _07653_ (.A(_02514_),
    .B(_03585_),
    .C(_03588_),
    .D(_03591_),
    .X(_03592_));
 sky130_fd_sc_hd__or3_1 _07654_ (.A(_02556_),
    .B(_02389_),
    .C(\mem[76][10] ),
    .X(_03593_));
 sky130_fd_sc_hd__o221a_1 _07655_ (.A1(\mem[78][10] ),
    .A2(_02370_),
    .B1(_02555_),
    .B2(\mem[79][10] ),
    .C1(_03593_),
    .X(_03594_));
 sky130_fd_sc_hd__o211a_1 _07656_ (.A1(\mem[77][10] ),
    .A2(_02639_),
    .B1(_03594_),
    .C1(_02422_),
    .X(_03595_));
 sky130_fd_sc_hd__o21a_1 _07657_ (.A1(\mem[64][10] ),
    .A2(_02395_),
    .B1(_02563_),
    .X(_03596_));
 sky130_fd_sc_hd__o22a_1 _07658_ (.A1(\mem[65][10] ),
    .A2(_02399_),
    .B1(_02566_),
    .B2(\mem[67][10] ),
    .X(_03597_));
 sky130_fd_sc_hd__o211a_1 _07659_ (.A1(\mem[66][10] ),
    .A2(_02394_),
    .B1(_03596_),
    .C1(_03597_),
    .X(_03598_));
 sky130_fd_sc_hd__or2_1 _07660_ (.A(\mem[72][10] ),
    .B(_02570_),
    .X(_03599_));
 sky130_fd_sc_hd__or3b_1 _07661_ (.A(_02802_),
    .B(\mem[74][10] ),
    .C_N(_02575_),
    .X(_03600_));
 sky130_fd_sc_hd__o221a_1 _07662_ (.A1(\mem[73][10] ),
    .A2(_02385_),
    .B1(_02801_),
    .B2(\mem[75][10] ),
    .C1(_03600_),
    .X(_03601_));
 sky130_fd_sc_hd__o21a_1 _07663_ (.A1(\mem[69][10] ),
    .A2(_02405_),
    .B1(_02463_),
    .X(_03602_));
 sky130_fd_sc_hd__or3_1 _07664_ (.A(_02411_),
    .B(_02868_),
    .C(\mem[68][10] ),
    .X(_03603_));
 sky130_fd_sc_hd__o221a_1 _07665_ (.A1(\mem[70][10] ),
    .A2(_02407_),
    .B1(_02409_),
    .B2(\mem[71][10] ),
    .C1(_03603_),
    .X(_03604_));
 sky130_fd_sc_hd__a32o_1 _07666_ (.A1(_02439_),
    .A2(_03599_),
    .A3(_03601_),
    .B1(_03602_),
    .B2(_03604_),
    .X(_03605_));
 sky130_fd_sc_hd__or4_1 _07667_ (.A(_02552_),
    .B(_03595_),
    .C(_03598_),
    .D(_03605_),
    .X(_03606_));
 sky130_fd_sc_hd__mux4_1 _07668_ (.A0(\mem[96][10] ),
    .A1(\mem[97][10] ),
    .A2(\mem[98][10] ),
    .A3(\mem[99][10] ),
    .S0(_02590_),
    .S1(_02591_),
    .X(_03607_));
 sky130_fd_sc_hd__mux4_1 _07669_ (.A0(\mem[100][10] ),
    .A1(\mem[101][10] ),
    .A2(\mem[102][10] ),
    .A3(\mem[103][10] ),
    .S0(_02593_),
    .S1(_02594_),
    .X(_03608_));
 sky130_fd_sc_hd__a22o_1 _07670_ (.A1(_02651_),
    .A2(_03607_),
    .B1(_03608_),
    .B2(_02825_),
    .X(_03609_));
 sky130_fd_sc_hd__mux4_1 _07671_ (.A0(\mem[108][10] ),
    .A1(\mem[109][10] ),
    .A2(\mem[110][10] ),
    .A3(\mem[111][10] ),
    .S0(_02458_),
    .S1(_02461_),
    .X(_03610_));
 sky130_fd_sc_hd__mux4_1 _07672_ (.A0(\mem[104][10] ),
    .A1(\mem[105][10] ),
    .A2(\mem[106][10] ),
    .A3(\mem[107][10] ),
    .S0(_02501_),
    .S1(_02877_),
    .X(_03611_));
 sky130_fd_sc_hd__or2_1 _07673_ (.A(_02474_),
    .B(_03611_),
    .X(_03612_));
 sky130_fd_sc_hd__o211a_1 _07674_ (.A1(_02598_),
    .A2(_03610_),
    .B1(_03612_),
    .C1(_02478_),
    .X(_03613_));
 sky130_fd_sc_hd__or3_2 _07675_ (.A(_02421_),
    .B(_03609_),
    .C(_03613_),
    .X(_03614_));
 sky130_fd_sc_hd__mux4_1 _07676_ (.A0(\mem[124][10] ),
    .A1(\mem[125][10] ),
    .A2(\mem[126][10] ),
    .A3(\mem[127][10] ),
    .S0(_02671_),
    .S1(_02703_),
    .X(_03615_));
 sky130_fd_sc_hd__mux4_1 _07677_ (.A0(\mem[112][10] ),
    .A1(\mem[113][10] ),
    .A2(\mem[114][10] ),
    .A3(\mem[115][10] ),
    .S0(_02726_),
    .S1(_02618_),
    .X(_03616_));
 sky130_fd_sc_hd__mux4_1 _07678_ (.A0(\mem[116][10] ),
    .A1(\mem[117][10] ),
    .A2(\mem[118][10] ),
    .A3(\mem[119][10] ),
    .S0(_02985_),
    .S1(_02623_),
    .X(_03617_));
 sky130_fd_sc_hd__mux4_1 _07679_ (.A0(\mem[120][10] ),
    .A1(\mem[121][10] ),
    .A2(\mem[122][10] ),
    .A3(\mem[123][10] ),
    .S0(_02887_),
    .S1(_02499_),
    .X(_03618_));
 sky130_fd_sc_hd__o22a_1 _07680_ (.A1(_02885_),
    .A2(_03617_),
    .B1(_03618_),
    .B2(_02889_),
    .X(_03619_));
 sky130_fd_sc_hd__o221a_2 _07681_ (.A1(_02612_),
    .A2(_03615_),
    .B1(_03616_),
    .B2(_02884_),
    .C1(_03619_),
    .X(_03620_));
 sky130_fd_sc_hd__o21a_1 _07682_ (.A1(_02358_),
    .A2(_03620_),
    .B1(_02509_),
    .X(_03621_));
 sky130_fd_sc_hd__a32o_1 _07683_ (.A1(_02355_),
    .A2(_03592_),
    .A3(_03606_),
    .B1(_03614_),
    .B2(_03621_),
    .X(_03622_));
 sky130_fd_sc_hd__mux2_1 _07684_ (.A0(_03578_),
    .A1(_03622_),
    .S(_02634_),
    .X(_03623_));
 sky130_fd_sc_hd__clkbuf_1 _07685_ (.A(_03623_),
    .X(_00001_));
 sky130_fd_sc_hd__o21a_1 _07686_ (.A1(\mem[29][11] ),
    .A2(_02515_),
    .B1(_02516_),
    .X(_03624_));
 sky130_fd_sc_hd__or3_1 _07687_ (.A(_02520_),
    .B(_02779_),
    .C(\mem[28][11] ),
    .X(_03625_));
 sky130_fd_sc_hd__o221a_1 _07688_ (.A1(\mem[30][11] ),
    .A2(_02995_),
    .B1(_02372_),
    .B2(\mem[31][11] ),
    .C1(_03625_),
    .X(_03626_));
 sky130_fd_sc_hd__o21a_1 _07689_ (.A1(\mem[16][11] ),
    .A2(_02524_),
    .B1(_02525_),
    .X(_03627_));
 sky130_fd_sc_hd__or3b_1 _07690_ (.A(_02529_),
    .B(\mem[18][11] ),
    .C_N(_02783_),
    .X(_03628_));
 sky130_fd_sc_hd__o221a_1 _07691_ (.A1(\mem[17][11] ),
    .A2(_02899_),
    .B1(_02528_),
    .B2(\mem[19][11] ),
    .C1(_03628_),
    .X(_03629_));
 sky130_fd_sc_hd__a22o_1 _07692_ (.A1(_03624_),
    .A2(_03626_),
    .B1(_03627_),
    .B2(_03629_),
    .X(_03630_));
 sky130_fd_sc_hd__o21a_1 _07693_ (.A1(\mem[24][11] ),
    .A2(_02788_),
    .B1(_02397_),
    .X(_03631_));
 sky130_fd_sc_hd__o22a_1 _07694_ (.A1(\mem[25][11] ),
    .A2(_02790_),
    .B1(_02539_),
    .B2(\mem[27][11] ),
    .X(_03632_));
 sky130_fd_sc_hd__o211a_1 _07695_ (.A1(\mem[26][11] ),
    .A2(_02787_),
    .B1(_03631_),
    .C1(_03632_),
    .X(_03633_));
 sky130_fd_sc_hd__or3_1 _07696_ (.A(_02793_),
    .B(_02412_),
    .C(\mem[20][11] ),
    .X(_03634_));
 sky130_fd_sc_hd__o221a_1 _07697_ (.A1(\mem[22][11] ),
    .A2(_02543_),
    .B1(_02544_),
    .B2(\mem[23][11] ),
    .C1(_03634_),
    .X(_03635_));
 sky130_fd_sc_hd__o211a_1 _07698_ (.A1(\mem[21][11] ),
    .A2(_02542_),
    .B1(_03635_),
    .C1(_02549_),
    .X(_03636_));
 sky130_fd_sc_hd__or4_4 _07699_ (.A(_02993_),
    .B(_03630_),
    .C(_03633_),
    .D(_03636_),
    .X(_03637_));
 sky130_fd_sc_hd__or3_1 _07700_ (.A(_02432_),
    .B(_02433_),
    .C(\mem[12][11] ),
    .X(_03638_));
 sky130_fd_sc_hd__o221a_1 _07701_ (.A1(\mem[14][11] ),
    .A2(_02800_),
    .B1(_03009_),
    .B2(\mem[15][11] ),
    .C1(_03638_),
    .X(_03639_));
 sky130_fd_sc_hd__o211a_1 _07702_ (.A1(\mem[13][11] ),
    .A2(_02799_),
    .B1(_03639_),
    .C1(_02806_),
    .X(_03640_));
 sky130_fd_sc_hd__o21a_1 _07703_ (.A1(\mem[0][11] ),
    .A2(_02562_),
    .B1(_03013_),
    .X(_03641_));
 sky130_fd_sc_hd__o22a_1 _07704_ (.A1(\mem[1][11] ),
    .A2(_02565_),
    .B1(_02914_),
    .B2(\mem[3][11] ),
    .X(_03642_));
 sky130_fd_sc_hd__o211a_1 _07705_ (.A1(\mem[2][11] ),
    .A2(_02561_),
    .B1(_03641_),
    .C1(_03642_),
    .X(_03643_));
 sky130_fd_sc_hd__or2_1 _07706_ (.A(\mem[8][11] ),
    .B(_02917_),
    .X(_03644_));
 sky130_fd_sc_hd__or3b_1 _07707_ (.A(_02574_),
    .B(\mem[10][11] ),
    .C_N(_02816_),
    .X(_03645_));
 sky130_fd_sc_hd__o221a_1 _07708_ (.A1(\mem[9][11] ),
    .A2(_02572_),
    .B1(_02573_),
    .B2(\mem[11][11] ),
    .C1(_03645_),
    .X(_03646_));
 sky130_fd_sc_hd__o21a_1 _07709_ (.A1(\mem[5][11] ),
    .A2(_02578_),
    .B1(_02579_),
    .X(_03647_));
 sky130_fd_sc_hd__or3_1 _07710_ (.A(_02583_),
    .B(_02584_),
    .C(\mem[4][11] ),
    .X(_03648_));
 sky130_fd_sc_hd__o221a_1 _07711_ (.A1(\mem[6][11] ),
    .A2(_02581_),
    .B1(_02446_),
    .B2(\mem[7][11] ),
    .C1(_03648_),
    .X(_03649_));
 sky130_fd_sc_hd__a32o_1 _07712_ (.A1(_02811_),
    .A2(_03644_),
    .A3(_03646_),
    .B1(_03647_),
    .B2(_03649_),
    .X(_03650_));
 sky130_fd_sc_hd__or4_1 _07713_ (.A(_02798_),
    .B(_03640_),
    .C(_03643_),
    .D(_03650_),
    .X(_03651_));
 sky130_fd_sc_hd__mux4_1 _07714_ (.A0(\mem[32][11] ),
    .A1(\mem[33][11] ),
    .A2(\mem[34][11] ),
    .A3(\mem[35][11] ),
    .S0(_02826_),
    .S1(_02926_),
    .X(_03652_));
 sky130_fd_sc_hd__mux4_1 _07715_ (.A0(\mem[36][11] ),
    .A1(\mem[37][11] ),
    .A2(\mem[38][11] ),
    .A3(\mem[39][11] ),
    .S0(_02928_),
    .S1(_02929_),
    .X(_03653_));
 sky130_fd_sc_hd__a22o_1 _07716_ (.A1(_02456_),
    .A2(_03652_),
    .B1(_03653_),
    .B2(_02465_),
    .X(_03654_));
 sky130_fd_sc_hd__mux4_1 _07717_ (.A0(\mem[44][11] ),
    .A1(\mem[45][11] ),
    .A2(\mem[46][11] ),
    .A3(\mem[47][11] ),
    .S0(_02600_),
    .S1(_02601_),
    .X(_03655_));
 sky130_fd_sc_hd__mux4_1 _07718_ (.A0(\mem[40][11] ),
    .A1(\mem[41][11] ),
    .A2(\mem[42][11] ),
    .A3(\mem[43][11] ),
    .S0(_02604_),
    .S1(_02605_),
    .X(_03656_));
 sky130_fd_sc_hd__or2_1 _07719_ (.A(_02603_),
    .B(_03656_),
    .X(_03657_));
 sky130_fd_sc_hd__o211a_1 _07720_ (.A1(_02599_),
    .A2(_03655_),
    .B1(_03657_),
    .C1(_02608_),
    .X(_03658_));
 sky130_fd_sc_hd__or3_2 _07721_ (.A(_02589_),
    .B(_03654_),
    .C(_03658_),
    .X(_03659_));
 sky130_fd_sc_hd__mux4_1 _07722_ (.A0(\mem[60][11] ),
    .A1(\mem[61][11] ),
    .A2(\mem[62][11] ),
    .A3(\mem[63][11] ),
    .S0(_02613_),
    .S1(_02614_),
    .X(_03660_));
 sky130_fd_sc_hd__mux4_1 _07723_ (.A0(\mem[48][11] ),
    .A1(\mem[49][11] ),
    .A2(\mem[50][11] ),
    .A3(\mem[51][11] ),
    .S0(_02616_),
    .S1(_02746_),
    .X(_03661_));
 sky130_fd_sc_hd__mux4_1 _07724_ (.A0(\mem[52][11] ),
    .A1(\mem[53][11] ),
    .A2(\mem[54][11] ),
    .A3(\mem[55][11] ),
    .S0(_02622_),
    .S1(_02837_),
    .X(_03662_));
 sky130_fd_sc_hd__mux4_1 _07725_ (.A0(\mem[56][11] ),
    .A1(\mem[57][11] ),
    .A2(\mem[58][11] ),
    .A3(\mem[59][11] ),
    .S0(_02625_),
    .S1(_02626_),
    .X(_03663_));
 sky130_fd_sc_hd__o22a_1 _07726_ (.A1(_02621_),
    .A2(_03662_),
    .B1(_03663_),
    .B2(_02628_),
    .X(_03664_));
 sky130_fd_sc_hd__o221a_1 _07727_ (.A1(_03033_),
    .A2(_03660_),
    .B1(_03661_),
    .B2(_02620_),
    .C1(_03664_),
    .X(_03665_));
 sky130_fd_sc_hd__o21a_1 _07728_ (.A1(_02611_),
    .A2(_03665_),
    .B1(_02631_),
    .X(_03666_));
 sky130_fd_sc_hd__a32o_1 _07729_ (.A1(_02513_),
    .A2(_03637_),
    .A3(_03651_),
    .B1(_03659_),
    .B2(_03666_),
    .X(_03667_));
 sky130_fd_sc_hd__o21a_1 _07730_ (.A1(\mem[93][11] ),
    .A2(_02565_),
    .B1(_02366_),
    .X(_03668_));
 sky130_fd_sc_hd__or3_1 _07731_ (.A(_02387_),
    .B(_02389_),
    .C(\mem[92][11] ),
    .X(_03669_));
 sky130_fd_sc_hd__o221a_1 _07732_ (.A1(\mem[94][11] ),
    .A2(_02370_),
    .B1(_02386_),
    .B2(\mem[95][11] ),
    .C1(_03669_),
    .X(_03670_));
 sky130_fd_sc_hd__o21a_1 _07733_ (.A1(\mem[80][11] ),
    .A2(_02438_),
    .B1(_02455_),
    .X(_03671_));
 sky130_fd_sc_hd__or3b_1 _07734_ (.A(_02815_),
    .B(\mem[82][11] ),
    .C_N(_03224_),
    .X(_03672_));
 sky130_fd_sc_hd__o221a_1 _07735_ (.A1(\mem[81][11] ),
    .A2(_02736_),
    .B1(_02814_),
    .B2(\mem[83][11] ),
    .C1(_03672_),
    .X(_03673_));
 sky130_fd_sc_hd__a22o_1 _07736_ (.A1(_03668_),
    .A2(_03670_),
    .B1(_03671_),
    .B2(_03673_),
    .X(_03674_));
 sky130_fd_sc_hd__o21a_1 _07737_ (.A1(\mem[88][11] ),
    .A2(_02438_),
    .B1(_02439_),
    .X(_03675_));
 sky130_fd_sc_hd__o22a_1 _07738_ (.A1(\mem[89][11] ),
    .A2(_02405_),
    .B1(_02442_),
    .B2(\mem[91][11] ),
    .X(_03676_));
 sky130_fd_sc_hd__o211a_1 _07739_ (.A1(\mem[90][11] ),
    .A2(_02437_),
    .B1(_03675_),
    .C1(_03676_),
    .X(_03677_));
 sky130_fd_sc_hd__or3_1 _07740_ (.A(_02427_),
    .B(_02429_),
    .C(\mem[84][11] ),
    .X(_03678_));
 sky130_fd_sc_hd__o221a_1 _07741_ (.A1(\mem[86][11] ),
    .A2(_02393_),
    .B1(_03231_),
    .B2(\mem[87][11] ),
    .C1(_03678_),
    .X(_03679_));
 sky130_fd_sc_hd__o211a_1 _07742_ (.A1(\mem[85][11] ),
    .A2(_02737_),
    .B1(_03679_),
    .C1(_02450_),
    .X(_03680_));
 sky130_fd_sc_hd__or4_2 _07743_ (.A(_02358_),
    .B(_03674_),
    .C(_03677_),
    .D(_03680_),
    .X(_03681_));
 sky130_fd_sc_hd__or3_1 _07744_ (.A(_02486_),
    .B(_03224_),
    .C(\mem[76][11] ),
    .X(_03682_));
 sky130_fd_sc_hd__o221a_1 _07745_ (.A1(\mem[78][11] ),
    .A2(_02800_),
    .B1(_02814_),
    .B2(\mem[79][11] ),
    .C1(_03682_),
    .X(_03683_));
 sky130_fd_sc_hd__o211a_1 _07746_ (.A1(\mem[77][11] ),
    .A2(_02799_),
    .B1(_03683_),
    .C1(_02806_),
    .X(_03684_));
 sky130_fd_sc_hd__o21a_1 _07747_ (.A1(\mem[64][11] ),
    .A2(_02438_),
    .B1(_02455_),
    .X(_03685_));
 sky130_fd_sc_hd__o22a_1 _07748_ (.A1(\mem[65][11] ),
    .A2(_02441_),
    .B1(_02442_),
    .B2(\mem[67][11] ),
    .X(_03686_));
 sky130_fd_sc_hd__o211a_1 _07749_ (.A1(\mem[66][11] ),
    .A2(_02437_),
    .B1(_03685_),
    .C1(_03686_),
    .X(_03687_));
 sky130_fd_sc_hd__or2_1 _07750_ (.A(\mem[72][11] ),
    .B(_02812_),
    .X(_03688_));
 sky130_fd_sc_hd__or3b_1 _07751_ (.A(_02486_),
    .B(\mem[74][11] ),
    .C_N(_03224_),
    .X(_03689_));
 sky130_fd_sc_hd__o221a_1 _07752_ (.A1(\mem[73][11] ),
    .A2(_03042_),
    .B1(_02814_),
    .B2(\mem[75][11] ),
    .C1(_03689_),
    .X(_03690_));
 sky130_fd_sc_hd__o21a_1 _07753_ (.A1(\mem[69][11] ),
    .A2(_02819_),
    .B1(_02416_),
    .X(_03691_));
 sky130_fd_sc_hd__or3_1 _07754_ (.A(_02447_),
    .B(_02429_),
    .C(\mem[68][11] ),
    .X(_03692_));
 sky130_fd_sc_hd__o221a_1 _07755_ (.A1(\mem[70][11] ),
    .A2(_02393_),
    .B1(_03231_),
    .B2(\mem[71][11] ),
    .C1(_03692_),
    .X(_03693_));
 sky130_fd_sc_hd__a32o_1 _07756_ (.A1(_02811_),
    .A2(_03688_),
    .A3(_03690_),
    .B1(_03691_),
    .B2(_03693_),
    .X(_03694_));
 sky130_fd_sc_hd__or4_1 _07757_ (.A(_02421_),
    .B(_03684_),
    .C(_03687_),
    .D(_03694_),
    .X(_03695_));
 sky130_fd_sc_hd__mux4_1 _07758_ (.A0(\mem[104][11] ),
    .A1(\mem[105][11] ),
    .A2(\mem[106][11] ),
    .A3(\mem[107][11] ),
    .S0(_02670_),
    .S1(_02488_),
    .X(_03696_));
 sky130_fd_sc_hd__or2_1 _07759_ (.A(_02475_),
    .B(_03696_),
    .X(_03697_));
 sky130_fd_sc_hd__mux4_1 _07760_ (.A0(\mem[108][11] ),
    .A1(\mem[109][11] ),
    .A2(\mem[110][11] ),
    .A3(\mem[111][11] ),
    .S0(_02374_),
    .S1(_02460_),
    .X(_03698_));
 sky130_fd_sc_hd__or2_1 _07761_ (.A(_02598_),
    .B(_03698_),
    .X(_03699_));
 sky130_fd_sc_hd__mux4_1 _07762_ (.A0(\mem[96][11] ),
    .A1(\mem[97][11] ),
    .A2(\mem[98][11] ),
    .A3(\mem[99][11] ),
    .S0(_02432_),
    .S1(_02488_),
    .X(_03700_));
 sky130_fd_sc_hd__mux4_1 _07763_ (.A0(\mem[100][11] ),
    .A1(\mem[101][11] ),
    .A2(\mem[102][11] ),
    .A3(\mem[103][11] ),
    .S0(_02411_),
    .S1(_02617_),
    .X(_03701_));
 sky130_fd_sc_hd__a22o_1 _07764_ (.A1(_02455_),
    .A2(_03700_),
    .B1(_03701_),
    .B2(_02464_),
    .X(_03702_));
 sky130_fd_sc_hd__a31o_1 _07765_ (.A1(_02479_),
    .A2(_03697_),
    .A3(_03699_),
    .B1(_03702_),
    .X(_03703_));
 sky130_fd_sc_hd__mux4_1 _07766_ (.A0(\mem[116][11] ),
    .A1(\mem[117][11] ),
    .A2(\mem[118][11] ),
    .A3(\mem[119][11] ),
    .S0(_02502_),
    .S1(_02503_),
    .X(_03704_));
 sky130_fd_sc_hd__mux4_1 _07767_ (.A0(\mem[120][11] ),
    .A1(\mem[121][11] ),
    .A2(\mem[122][11] ),
    .A3(\mem[123][11] ),
    .S0(_02502_),
    .S1(_02673_),
    .X(_03705_));
 sky130_fd_sc_hd__o22a_1 _07768_ (.A1(_02498_),
    .A2(_03704_),
    .B1(_03705_),
    .B2(_02506_),
    .X(_03706_));
 sky130_fd_sc_hd__mux4_1 _07769_ (.A0(\mem[124][11] ),
    .A1(\mem[125][11] ),
    .A2(\mem[126][11] ),
    .A3(\mem[127][11] ),
    .S0(_02427_),
    .S1(_02499_),
    .X(_03707_));
 sky130_fd_sc_hd__mux4_2 _07770_ (.A0(\mem[112][11] ),
    .A1(\mem[113][11] ),
    .A2(\mem[114][11] ),
    .A3(\mem[115][11] ),
    .S0(_02502_),
    .S1(_02673_),
    .X(_03708_));
 sky130_fd_sc_hd__o22a_1 _07771_ (.A1(_02484_),
    .A2(_03707_),
    .B1(_03708_),
    .B2(_02495_),
    .X(_03709_));
 sky130_fd_sc_hd__a21o_2 _07772_ (.A1(_03706_),
    .A2(_03709_),
    .B1(_02357_),
    .X(_03710_));
 sky130_fd_sc_hd__o211a_1 _07773_ (.A1(_02453_),
    .A2(_03703_),
    .B1(_03710_),
    .C1(_02509_),
    .X(_03711_));
 sky130_fd_sc_hd__a31o_1 _07774_ (.A1(_02356_),
    .A2(_03681_),
    .A3(_03695_),
    .B1(_03711_),
    .X(_03712_));
 sky130_fd_sc_hd__mux2_1 _07775_ (.A0(_03667_),
    .A1(_03712_),
    .S(_02634_),
    .X(_03713_));
 sky130_fd_sc_hd__clkbuf_1 _07776_ (.A(_03713_),
    .X(_00002_));
 sky130_fd_sc_hd__o21a_1 _07777_ (.A1(\mem[29][12] ),
    .A2(_02515_),
    .B1(_02516_),
    .X(_03714_));
 sky130_fd_sc_hd__or3_1 _07778_ (.A(_02520_),
    .B(_02779_),
    .C(\mem[28][12] ),
    .X(_03715_));
 sky130_fd_sc_hd__o221a_1 _07779_ (.A1(\mem[30][12] ),
    .A2(_02995_),
    .B1(_02519_),
    .B2(\mem[31][12] ),
    .C1(_03715_),
    .X(_03716_));
 sky130_fd_sc_hd__o21a_1 _07780_ (.A1(\mem[16][12] ),
    .A2(_02524_),
    .B1(_02525_),
    .X(_03717_));
 sky130_fd_sc_hd__or3b_1 _07781_ (.A(_02529_),
    .B(\mem[18][12] ),
    .C_N(_02783_),
    .X(_03718_));
 sky130_fd_sc_hd__o221a_1 _07782_ (.A1(\mem[17][12] ),
    .A2(_02899_),
    .B1(_02528_),
    .B2(\mem[19][12] ),
    .C1(_03718_),
    .X(_03719_));
 sky130_fd_sc_hd__a22o_1 _07783_ (.A1(_03714_),
    .A2(_03716_),
    .B1(_03717_),
    .B2(_03719_),
    .X(_03720_));
 sky130_fd_sc_hd__o21a_1 _07784_ (.A1(\mem[24][12] ),
    .A2(_02788_),
    .B1(_02536_),
    .X(_03721_));
 sky130_fd_sc_hd__o22a_1 _07785_ (.A1(\mem[25][12] ),
    .A2(_02790_),
    .B1(_02539_),
    .B2(\mem[27][12] ),
    .X(_03722_));
 sky130_fd_sc_hd__o211a_1 _07786_ (.A1(\mem[26][12] ),
    .A2(_02787_),
    .B1(_03721_),
    .C1(_03722_),
    .X(_03723_));
 sky130_fd_sc_hd__or3_1 _07787_ (.A(_02793_),
    .B(_02546_),
    .C(\mem[20][12] ),
    .X(_03724_));
 sky130_fd_sc_hd__o221a_1 _07788_ (.A1(\mem[22][12] ),
    .A2(_02543_),
    .B1(_02544_),
    .B2(\mem[23][12] ),
    .C1(_03724_),
    .X(_03725_));
 sky130_fd_sc_hd__o211a_1 _07789_ (.A1(\mem[21][12] ),
    .A2(_02542_),
    .B1(_03725_),
    .C1(_02549_),
    .X(_03726_));
 sky130_fd_sc_hd__or4_4 _07790_ (.A(_02993_),
    .B(_03720_),
    .C(_03723_),
    .D(_03726_),
    .X(_03727_));
 sky130_fd_sc_hd__or3_1 _07791_ (.A(_02432_),
    .B(_02433_),
    .C(\mem[12][12] ),
    .X(_03728_));
 sky130_fd_sc_hd__o221a_1 _07792_ (.A1(\mem[14][12] ),
    .A2(_02554_),
    .B1(_03009_),
    .B2(\mem[15][12] ),
    .C1(_03728_),
    .X(_03729_));
 sky130_fd_sc_hd__o211a_1 _07793_ (.A1(\mem[13][12] ),
    .A2(_02553_),
    .B1(_03729_),
    .C1(_02559_),
    .X(_03730_));
 sky130_fd_sc_hd__o21a_1 _07794_ (.A1(\mem[0][12] ),
    .A2(_02562_),
    .B1(_03013_),
    .X(_03731_));
 sky130_fd_sc_hd__o22a_1 _07795_ (.A1(\mem[1][12] ),
    .A2(_02565_),
    .B1(_02914_),
    .B2(\mem[3][12] ),
    .X(_03732_));
 sky130_fd_sc_hd__o211a_1 _07796_ (.A1(\mem[2][12] ),
    .A2(_02561_),
    .B1(_03731_),
    .C1(_03732_),
    .X(_03733_));
 sky130_fd_sc_hd__or2_1 _07797_ (.A(\mem[8][12] ),
    .B(_02917_),
    .X(_03734_));
 sky130_fd_sc_hd__or3b_1 _07798_ (.A(_02574_),
    .B(\mem[10][12] ),
    .C_N(_02816_),
    .X(_03735_));
 sky130_fd_sc_hd__o221a_1 _07799_ (.A1(\mem[9][12] ),
    .A2(_02572_),
    .B1(_02573_),
    .B2(\mem[11][12] ),
    .C1(_03735_),
    .X(_03736_));
 sky130_fd_sc_hd__o21a_1 _07800_ (.A1(\mem[5][12] ),
    .A2(_02578_),
    .B1(_02579_),
    .X(_03737_));
 sky130_fd_sc_hd__or3_1 _07801_ (.A(_02583_),
    .B(_02584_),
    .C(\mem[4][12] ),
    .X(_03738_));
 sky130_fd_sc_hd__o221a_1 _07802_ (.A1(\mem[6][12] ),
    .A2(_02581_),
    .B1(_02582_),
    .B2(\mem[7][12] ),
    .C1(_03738_),
    .X(_03739_));
 sky130_fd_sc_hd__a32o_2 _07803_ (.A1(_02569_),
    .A2(_03734_),
    .A3(_03736_),
    .B1(_03737_),
    .B2(_03739_),
    .X(_03740_));
 sky130_fd_sc_hd__or4_1 _07804_ (.A(_02798_),
    .B(_03730_),
    .C(_03733_),
    .D(_03740_),
    .X(_03741_));
 sky130_fd_sc_hd__mux4_1 _07805_ (.A0(\mem[36][12] ),
    .A1(\mem[37][12] ),
    .A2(\mem[38][12] ),
    .A3(\mem[39][12] ),
    .S0(_02826_),
    .S1(_02926_),
    .X(_03742_));
 sky130_fd_sc_hd__mux4_1 _07806_ (.A0(\mem[32][12] ),
    .A1(\mem[33][12] ),
    .A2(\mem[34][12] ),
    .A3(\mem[35][12] ),
    .S0(_02928_),
    .S1(_02929_),
    .X(_03743_));
 sky130_fd_sc_hd__a22o_1 _07807_ (.A1(_02450_),
    .A2(_03742_),
    .B1(_03743_),
    .B2(_02596_),
    .X(_03744_));
 sky130_fd_sc_hd__mux4_1 _07808_ (.A0(\mem[44][12] ),
    .A1(\mem[45][12] ),
    .A2(\mem[46][12] ),
    .A3(\mem[47][12] ),
    .S0(_02600_),
    .S1(_02601_),
    .X(_03745_));
 sky130_fd_sc_hd__mux4_1 _07809_ (.A0(\mem[40][12] ),
    .A1(\mem[41][12] ),
    .A2(\mem[42][12] ),
    .A3(\mem[43][12] ),
    .S0(_02604_),
    .S1(_02605_),
    .X(_03746_));
 sky130_fd_sc_hd__or2_1 _07810_ (.A(_02603_),
    .B(_03746_),
    .X(_03747_));
 sky130_fd_sc_hd__o211a_1 _07811_ (.A1(_02599_),
    .A2(_03745_),
    .B1(_03747_),
    .C1(_02608_),
    .X(_03748_));
 sky130_fd_sc_hd__or3_4 _07812_ (.A(_02589_),
    .B(_03744_),
    .C(_03748_),
    .X(_03749_));
 sky130_fd_sc_hd__mux4_1 _07813_ (.A0(\mem[60][12] ),
    .A1(\mem[61][12] ),
    .A2(\mem[62][12] ),
    .A3(\mem[63][12] ),
    .S0(_02613_),
    .S1(_02614_),
    .X(_03750_));
 sky130_fd_sc_hd__mux4_1 _07814_ (.A0(\mem[48][12] ),
    .A1(\mem[49][12] ),
    .A2(\mem[50][12] ),
    .A3(\mem[51][12] ),
    .S0(_02616_),
    .S1(_02746_),
    .X(_03751_));
 sky130_fd_sc_hd__mux4_1 _07815_ (.A0(\mem[52][12] ),
    .A1(\mem[53][12] ),
    .A2(\mem[54][12] ),
    .A3(\mem[55][12] ),
    .S0(_02622_),
    .S1(_02837_),
    .X(_03752_));
 sky130_fd_sc_hd__mux4_1 _07816_ (.A0(\mem[56][12] ),
    .A1(\mem[57][12] ),
    .A2(\mem[58][12] ),
    .A3(\mem[59][12] ),
    .S0(_02625_),
    .S1(_02626_),
    .X(_03753_));
 sky130_fd_sc_hd__o22a_1 _07817_ (.A1(_02621_),
    .A2(_03752_),
    .B1(_03753_),
    .B2(_02628_),
    .X(_03754_));
 sky130_fd_sc_hd__o221a_1 _07818_ (.A1(_03033_),
    .A2(_03750_),
    .B1(_03751_),
    .B2(_02620_),
    .C1(_03754_),
    .X(_03755_));
 sky130_fd_sc_hd__o21a_1 _07819_ (.A1(_02611_),
    .A2(_03755_),
    .B1(_02631_),
    .X(_03756_));
 sky130_fd_sc_hd__a32o_1 _07820_ (.A1(_02513_),
    .A2(_03727_),
    .A3(_03741_),
    .B1(_03749_),
    .B2(_03756_),
    .X(_03757_));
 sky130_fd_sc_hd__o21a_1 _07821_ (.A1(\mem[93][12] ),
    .A2(_03042_),
    .B1(_02365_),
    .X(_03758_));
 sky130_fd_sc_hd__or3_1 _07822_ (.A(_02466_),
    .B(_02459_),
    .C(\mem[92][12] ),
    .X(_03759_));
 sky130_fd_sc_hd__o221a_1 _07823_ (.A1(\mem[94][12] ),
    .A2(_02518_),
    .B1(_02400_),
    .B2(\mem[95][12] ),
    .C1(_03759_),
    .X(_03760_));
 sky130_fd_sc_hd__o21a_1 _07824_ (.A1(\mem[80][12] ),
    .A2(_02812_),
    .B1(_02454_),
    .X(_03761_));
 sky130_fd_sc_hd__or3b_1 _07825_ (.A(_02670_),
    .B(\mem[82][12] ),
    .C_N(_02375_),
    .X(_03762_));
 sky130_fd_sc_hd__o221a_1 _07826_ (.A1(\mem[81][12] ),
    .A2(_02527_),
    .B1(_02424_),
    .B2(\mem[83][12] ),
    .C1(_03762_),
    .X(_03763_));
 sky130_fd_sc_hd__a22o_1 _07827_ (.A1(_03758_),
    .A2(_03760_),
    .B1(_03761_),
    .B2(_03763_),
    .X(_03764_));
 sky130_fd_sc_hd__o21a_1 _07828_ (.A1(\mem[88][12] ),
    .A2(_02380_),
    .B1(_02396_),
    .X(_03765_));
 sky130_fd_sc_hd__o22a_1 _07829_ (.A1(\mem[89][12] ),
    .A2(_02363_),
    .B1(_03231_),
    .B2(\mem[91][12] ),
    .X(_03766_));
 sky130_fd_sc_hd__o211a_1 _07830_ (.A1(\mem[90][12] ),
    .A2(_02660_),
    .B1(_03765_),
    .C1(_03766_),
    .X(_03767_));
 sky130_fd_sc_hd__or3_1 _07831_ (.A(_02486_),
    .B(_03224_),
    .C(\mem[84][12] ),
    .X(_03768_));
 sky130_fd_sc_hd__o221a_1 _07832_ (.A1(\mem[86][12] ),
    .A2(_02956_),
    .B1(_02664_),
    .B2(\mem[87][12] ),
    .C1(_03768_),
    .X(_03769_));
 sky130_fd_sc_hd__o211a_1 _07833_ (.A1(\mem[85][12] ),
    .A2(_02955_),
    .B1(_03769_),
    .C1(_02464_),
    .X(_03770_));
 sky130_fd_sc_hd__or4_2 _07834_ (.A(_02514_),
    .B(_03764_),
    .C(_03767_),
    .D(_03770_),
    .X(_03771_));
 sky130_fd_sc_hd__or3_1 _07835_ (.A(_02556_),
    .B(_02389_),
    .C(\mem[76][12] ),
    .X(_03772_));
 sky130_fd_sc_hd__o221a_1 _07836_ (.A1(\mem[78][12] ),
    .A2(_02370_),
    .B1(_02555_),
    .B2(\mem[79][12] ),
    .C1(_03772_),
    .X(_03773_));
 sky130_fd_sc_hd__o211a_1 _07837_ (.A1(\mem[77][12] ),
    .A2(_02639_),
    .B1(_03773_),
    .C1(_02422_),
    .X(_03774_));
 sky130_fd_sc_hd__o21a_1 _07838_ (.A1(\mem[64][12] ),
    .A2(_02395_),
    .B1(_02563_),
    .X(_03775_));
 sky130_fd_sc_hd__o22a_1 _07839_ (.A1(\mem[65][12] ),
    .A2(_02399_),
    .B1(_02566_),
    .B2(\mem[67][12] ),
    .X(_03776_));
 sky130_fd_sc_hd__o211a_1 _07840_ (.A1(\mem[66][12] ),
    .A2(_02394_),
    .B1(_03775_),
    .C1(_03776_),
    .X(_03777_));
 sky130_fd_sc_hd__or2_1 _07841_ (.A(\mem[72][12] ),
    .B(_02570_),
    .X(_03778_));
 sky130_fd_sc_hd__or3b_1 _07842_ (.A(_02802_),
    .B(\mem[74][12] ),
    .C_N(_02803_),
    .X(_03779_));
 sky130_fd_sc_hd__o221a_1 _07843_ (.A1(\mem[73][12] ),
    .A2(_02385_),
    .B1(_02801_),
    .B2(\mem[75][12] ),
    .C1(_03779_),
    .X(_03780_));
 sky130_fd_sc_hd__o21a_1 _07844_ (.A1(\mem[69][12] ),
    .A2(_02405_),
    .B1(_02463_),
    .X(_03781_));
 sky130_fd_sc_hd__or3_1 _07845_ (.A(_02411_),
    .B(_02868_),
    .C(\mem[68][12] ),
    .X(_03782_));
 sky130_fd_sc_hd__o221a_1 _07846_ (.A1(\mem[70][12] ),
    .A2(_02407_),
    .B1(_02409_),
    .B2(\mem[71][12] ),
    .C1(_03782_),
    .X(_03783_));
 sky130_fd_sc_hd__a32o_1 _07847_ (.A1(_02439_),
    .A2(_03778_),
    .A3(_03780_),
    .B1(_03781_),
    .B2(_03783_),
    .X(_03784_));
 sky130_fd_sc_hd__or4_1 _07848_ (.A(_02420_),
    .B(_03774_),
    .C(_03777_),
    .D(_03784_),
    .X(_03785_));
 sky130_fd_sc_hd__mux4_1 _07849_ (.A0(\mem[96][12] ),
    .A1(\mem[97][12] ),
    .A2(\mem[98][12] ),
    .A3(\mem[99][12] ),
    .S0(_02645_),
    .S1(_02591_),
    .X(_03786_));
 sky130_fd_sc_hd__mux4_1 _07850_ (.A0(\mem[100][12] ),
    .A1(\mem[101][12] ),
    .A2(\mem[102][12] ),
    .A3(\mem[103][12] ),
    .S0(_02593_),
    .S1(_02594_),
    .X(_03787_));
 sky130_fd_sc_hd__a22o_1 _07851_ (.A1(_02651_),
    .A2(_03786_),
    .B1(_03787_),
    .B2(_02825_),
    .X(_03788_));
 sky130_fd_sc_hd__mux4_1 _07852_ (.A0(\mem[108][12] ),
    .A1(\mem[109][12] ),
    .A2(\mem[110][12] ),
    .A3(\mem[111][12] ),
    .S0(_02458_),
    .S1(_02461_),
    .X(_03789_));
 sky130_fd_sc_hd__mux4_1 _07853_ (.A0(\mem[104][12] ),
    .A1(\mem[105][12] ),
    .A2(\mem[106][12] ),
    .A3(\mem[107][12] ),
    .S0(_02501_),
    .S1(_02877_),
    .X(_03790_));
 sky130_fd_sc_hd__or2_1 _07854_ (.A(_02474_),
    .B(_03790_),
    .X(_03791_));
 sky130_fd_sc_hd__o211a_1 _07855_ (.A1(_02598_),
    .A2(_03789_),
    .B1(_03791_),
    .C1(_02478_),
    .X(_03792_));
 sky130_fd_sc_hd__or3_2 _07856_ (.A(_02421_),
    .B(_03788_),
    .C(_03792_),
    .X(_03793_));
 sky130_fd_sc_hd__mux4_1 _07857_ (.A0(\mem[124][12] ),
    .A1(\mem[125][12] ),
    .A2(\mem[126][12] ),
    .A3(\mem[127][12] ),
    .S0(_02671_),
    .S1(_02703_),
    .X(_03794_));
 sky130_fd_sc_hd__mux4_1 _07858_ (.A0(\mem[112][12] ),
    .A1(\mem[113][12] ),
    .A2(\mem[114][12] ),
    .A3(\mem[115][12] ),
    .S0(_02726_),
    .S1(_02618_),
    .X(_03795_));
 sky130_fd_sc_hd__mux4_1 _07859_ (.A0(\mem[116][12] ),
    .A1(\mem[117][12] ),
    .A2(\mem[118][12] ),
    .A3(\mem[119][12] ),
    .S0(_02985_),
    .S1(_02617_),
    .X(_03796_));
 sky130_fd_sc_hd__mux4_1 _07860_ (.A0(\mem[120][12] ),
    .A1(\mem[121][12] ),
    .A2(\mem[122][12] ),
    .A3(\mem[123][12] ),
    .S0(_02887_),
    .S1(_02499_),
    .X(_03797_));
 sky130_fd_sc_hd__o22a_1 _07861_ (.A1(_02885_),
    .A2(_03796_),
    .B1(_03797_),
    .B2(_02889_),
    .X(_03798_));
 sky130_fd_sc_hd__o221a_2 _07862_ (.A1(_02612_),
    .A2(_03794_),
    .B1(_03795_),
    .B2(_02884_),
    .C1(_03798_),
    .X(_03799_));
 sky130_fd_sc_hd__o21a_1 _07863_ (.A1(_02358_),
    .A2(_03799_),
    .B1(_02509_),
    .X(_03800_));
 sky130_fd_sc_hd__a32o_1 _07864_ (.A1(_02355_),
    .A2(_03771_),
    .A3(_03785_),
    .B1(_03793_),
    .B2(_03800_),
    .X(_03801_));
 sky130_fd_sc_hd__mux2_1 _07865_ (.A0(_03757_),
    .A1(_03801_),
    .S(_02634_),
    .X(_03802_));
 sky130_fd_sc_hd__clkbuf_1 _07866_ (.A(_03802_),
    .X(_00003_));
 sky130_fd_sc_hd__o21a_1 _07867_ (.A1(\mem[93][13] ),
    .A2(_02654_),
    .B1(_02641_),
    .X(_03803_));
 sky130_fd_sc_hd__or3_1 _07868_ (.A(_02646_),
    .B(_02489_),
    .C(\mem[92][13] ),
    .X(_03804_));
 sky130_fd_sc_hd__o221a_1 _07869_ (.A1(\mem[94][13] ),
    .A2(_02437_),
    .B1(_02644_),
    .B2(\mem[95][13] ),
    .C1(_03804_),
    .X(_03805_));
 sky130_fd_sc_hd__o21a_1 _07870_ (.A1(\mem[80][13] ),
    .A2(_02650_),
    .B1(_02596_),
    .X(_03806_));
 sky130_fd_sc_hd__or3b_1 _07871_ (.A(_02646_),
    .B(\mem[82][13] ),
    .C_N(_02492_),
    .X(_03807_));
 sky130_fd_sc_hd__o221a_1 _07872_ (.A1(\mem[81][13] ),
    .A2(_02654_),
    .B1(_03092_),
    .B2(\mem[83][13] ),
    .C1(_03807_),
    .X(_03808_));
 sky130_fd_sc_hd__a22o_1 _07873_ (.A1(_03803_),
    .A2(_03805_),
    .B1(_03806_),
    .B2(_03808_),
    .X(_03809_));
 sky130_fd_sc_hd__o21a_1 _07874_ (.A1(\mem[88][13] ),
    .A2(_02650_),
    .B1(_02662_),
    .X(_03810_));
 sky130_fd_sc_hd__o22a_1 _07875_ (.A1(\mem[89][13] ),
    .A2(_02640_),
    .B1(_02666_),
    .B2(\mem[91][13] ),
    .X(_03811_));
 sky130_fd_sc_hd__o211a_1 _07876_ (.A1(\mem[90][13] ),
    .A2(_02661_),
    .B1(_03810_),
    .C1(_03811_),
    .X(_03812_));
 sky130_fd_sc_hd__or3_1 _07877_ (.A(_02672_),
    .B(_02682_),
    .C(\mem[84][13] ),
    .X(_03813_));
 sky130_fd_sc_hd__o221a_1 _07878_ (.A1(\mem[86][13] ),
    .A2(_02643_),
    .B1(_02655_),
    .B2(\mem[87][13] ),
    .C1(_03813_),
    .X(_03814_));
 sky130_fd_sc_hd__o211a_1 _07879_ (.A1(\mem[85][13] ),
    .A2(_02669_),
    .B1(_03814_),
    .C1(_02677_),
    .X(_03815_));
 sky130_fd_sc_hd__nor4_4 _07880_ (.A(_02638_),
    .B(_03809_),
    .C(_03812_),
    .D(_03815_),
    .Y(_03816_));
 sky130_fd_sc_hd__or3_1 _07881_ (.A(_02681_),
    .B(_02682_),
    .C(\mem[76][13] ),
    .X(_03817_));
 sky130_fd_sc_hd__o221a_1 _07882_ (.A1(\mem[78][13] ),
    .A2(_02643_),
    .B1(_02655_),
    .B2(\mem[79][13] ),
    .C1(_03817_),
    .X(_03818_));
 sky130_fd_sc_hd__o211a_1 _07883_ (.A1(\mem[77][13] ),
    .A2(_02669_),
    .B1(_03818_),
    .C1(_02641_),
    .X(_03819_));
 sky130_fd_sc_hd__o21a_1 _07884_ (.A1(\mem[64][13] ),
    .A2(_02650_),
    .B1(_02652_),
    .X(_03820_));
 sky130_fd_sc_hd__o22a_1 _07885_ (.A1(\mem[65][13] ),
    .A2(_02640_),
    .B1(_02666_),
    .B2(\mem[67][13] ),
    .X(_03821_));
 sky130_fd_sc_hd__o211a_1 _07886_ (.A1(\mem[66][13] ),
    .A2(_02661_),
    .B1(_03820_),
    .C1(_03821_),
    .X(_03822_));
 sky130_fd_sc_hd__or2_1 _07887_ (.A(\mem[72][13] ),
    .B(_02649_),
    .X(_03823_));
 sky130_fd_sc_hd__or3b_1 _07888_ (.A(_02672_),
    .B(\mem[74][13] ),
    .C_N(_02682_),
    .X(_03824_));
 sky130_fd_sc_hd__o221a_1 _07889_ (.A1(\mem[73][13] ),
    .A2(_02654_),
    .B1(_02655_),
    .B2(\mem[75][13] ),
    .C1(_03824_),
    .X(_03825_));
 sky130_fd_sc_hd__o21a_1 _07890_ (.A1(\mem[69][13] ),
    .A2(_02669_),
    .B1(_02465_),
    .X(_03826_));
 sky130_fd_sc_hd__or3_1 _07891_ (.A(_02693_),
    .B(_02674_),
    .C(\mem[68][13] ),
    .X(_03827_));
 sky130_fd_sc_hd__o221a_1 _07892_ (.A1(\mem[70][13] ),
    .A2(_02643_),
    .B1(_02666_),
    .B2(\mem[71][13] ),
    .C1(_03827_),
    .X(_03828_));
 sky130_fd_sc_hd__a32o_1 _07893_ (.A1(_02662_),
    .A2(_03823_),
    .A3(_03825_),
    .B1(_03826_),
    .B2(_03828_),
    .X(_03829_));
 sky130_fd_sc_hd__nor4_2 _07894_ (.A(_02680_),
    .B(_03819_),
    .C(_03822_),
    .D(_03829_),
    .Y(_03830_));
 sky130_fd_sc_hd__mux4_1 _07895_ (.A0(\mem[124][13] ),
    .A1(\mem[125][13] ),
    .A2(\mem[126][13] ),
    .A3(\mem[127][13] ),
    .S0(_02711_),
    .S1(_02699_),
    .X(_03831_));
 sky130_fd_sc_hd__mux4_1 _07896_ (.A0(\mem[112][13] ),
    .A1(\mem[113][13] ),
    .A2(\mem[114][13] ),
    .A3(\mem[115][13] ),
    .S0(_02698_),
    .S1(_02699_),
    .X(_03832_));
 sky130_fd_sc_hd__mux4_1 _07897_ (.A0(\mem[116][13] ),
    .A1(\mem[117][13] ),
    .A2(\mem[118][13] ),
    .A3(\mem[119][13] ),
    .S0(_02681_),
    .S1(_02743_),
    .X(_03833_));
 sky130_fd_sc_hd__mux4_1 _07898_ (.A0(\mem[120][13] ),
    .A1(\mem[121][13] ),
    .A2(\mem[122][13] ),
    .A3(\mem[123][13] ),
    .S0(_02672_),
    .S1(_02704_),
    .X(_03834_));
 sky130_fd_sc_hd__o22a_1 _07899_ (.A1(_02702_),
    .A2(_03833_),
    .B1(_03834_),
    .B2(_02707_),
    .X(_03835_));
 sky130_fd_sc_hd__o221a_1 _07900_ (.A1(_02485_),
    .A2(_03831_),
    .B1(_03832_),
    .B2(_02496_),
    .C1(_03835_),
    .X(_03836_));
 sky130_fd_sc_hd__nor2_1 _07901_ (.A(_02638_),
    .B(_03836_),
    .Y(_03837_));
 sky130_fd_sc_hd__mux4_1 _07902_ (.A0(\mem[100][13] ),
    .A1(\mem[101][13] ),
    .A2(\mem[102][13] ),
    .A3(\mem[103][13] ),
    .S0(_02749_),
    .S1(_02712_),
    .X(_03838_));
 sky130_fd_sc_hd__mux4_1 _07903_ (.A0(\mem[96][13] ),
    .A1(\mem[97][13] ),
    .A2(\mem[98][13] ),
    .A3(\mem[99][13] ),
    .S0(_02711_),
    .S1(_02712_),
    .X(_03839_));
 sky130_fd_sc_hd__a22o_1 _07904_ (.A1(_02677_),
    .A2(_03838_),
    .B1(_03839_),
    .B2(_02652_),
    .X(_03840_));
 sky130_fd_sc_hd__mux4_1 _07905_ (.A0(\mem[108][13] ),
    .A1(\mem[109][13] ),
    .A2(\mem[110][13] ),
    .A3(\mem[111][13] ),
    .S0(_02711_),
    .S1(_02712_),
    .X(_03841_));
 sky130_fd_sc_hd__mux4_1 _07906_ (.A0(\mem[104][13] ),
    .A1(\mem[105][13] ),
    .A2(\mem[106][13] ),
    .A3(\mem[107][13] ),
    .S0(_02428_),
    .S1(_02674_),
    .X(_03842_));
 sky130_fd_sc_hd__or2_1 _07907_ (.A(_02718_),
    .B(_03842_),
    .X(_03843_));
 sky130_fd_sc_hd__o211a_1 _07908_ (.A1(_02716_),
    .A2(_03841_),
    .B1(_03843_),
    .C1(_02721_),
    .X(_03844_));
 sky130_fd_sc_hd__o31ai_2 _07909_ (.A1(_02680_),
    .A2(_03840_),
    .A3(_03844_),
    .B1(_02637_),
    .Y(_03845_));
 sky130_fd_sc_hd__o32a_1 _07910_ (.A1(_02637_),
    .A2(_03816_),
    .A3(_03830_),
    .B1(_03837_),
    .B2(_03845_),
    .X(_03846_));
 sky130_fd_sc_hd__or3_1 _07911_ (.A(_02726_),
    .B(_02673_),
    .C(\mem[28][13] ),
    .X(_03847_));
 sky130_fd_sc_hd__o221a_1 _07912_ (.A1(\mem[30][13] ),
    .A2(_02660_),
    .B1(_02665_),
    .B2(\mem[31][13] ),
    .C1(_03847_),
    .X(_03848_));
 sky130_fd_sc_hd__o211a_1 _07913_ (.A1(\mem[29][13] ),
    .A2(_02640_),
    .B1(_03848_),
    .C1(_02641_),
    .X(_03849_));
 sky130_fd_sc_hd__o21a_1 _07914_ (.A1(\mem[16][13] ),
    .A2(_02649_),
    .B1(_02651_),
    .X(_03850_));
 sky130_fd_sc_hd__o22a_1 _07915_ (.A1(\mem[17][13] ),
    .A2(_02406_),
    .B1(_02665_),
    .B2(\mem[19][13] ),
    .X(_03851_));
 sky130_fd_sc_hd__o211a_1 _07916_ (.A1(\mem[18][13] ),
    .A2(_02661_),
    .B1(_03850_),
    .C1(_03851_),
    .X(_03852_));
 sky130_fd_sc_hd__or2_1 _07917_ (.A(\mem[24][13] ),
    .B(_02649_),
    .X(_03853_));
 sky130_fd_sc_hd__or3b_1 _07918_ (.A(_02671_),
    .B(\mem[26][13] ),
    .C_N(_02673_),
    .X(_03854_));
 sky130_fd_sc_hd__o221a_1 _07919_ (.A1(\mem[25][13] ),
    .A2(_02639_),
    .B1(_02442_),
    .B2(\mem[27][13] ),
    .C1(_03854_),
    .X(_03855_));
 sky130_fd_sc_hd__o21a_1 _07920_ (.A1(\mem[21][13] ),
    .A2(_02737_),
    .B1(_02417_),
    .X(_03856_));
 sky130_fd_sc_hd__or3_1 _07921_ (.A(_02491_),
    .B(_02430_),
    .C(\mem[20][13] ),
    .X(_03857_));
 sky130_fd_sc_hd__o221a_1 _07922_ (.A1(\mem[22][13] ),
    .A2(_02660_),
    .B1(_02665_),
    .B2(\mem[23][13] ),
    .C1(_03857_),
    .X(_03858_));
 sky130_fd_sc_hd__a32o_1 _07923_ (.A1(_02662_),
    .A2(_03853_),
    .A3(_03855_),
    .B1(_03856_),
    .B2(_03858_),
    .X(_03859_));
 sky130_fd_sc_hd__or3_2 _07924_ (.A(_03849_),
    .B(_03852_),
    .C(_03859_),
    .X(_03860_));
 sky130_fd_sc_hd__mux4_1 _07925_ (.A0(\mem[8][13] ),
    .A1(\mem[9][13] ),
    .A2(\mem[10][13] ),
    .A3(\mem[11][13] ),
    .S0(_02646_),
    .S1(_02674_),
    .X(_03861_));
 sky130_fd_sc_hd__or2_1 _07926_ (.A(_02718_),
    .B(_03861_),
    .X(_03862_));
 sky130_fd_sc_hd__mux2_1 _07927_ (.A0(\mem[14][13] ),
    .A1(\mem[15][13] ),
    .S(_02749_),
    .X(_03863_));
 sky130_fd_sc_hd__mux2_1 _07928_ (.A0(\mem[12][13] ),
    .A1(\mem[13][13] ),
    .S(_02428_),
    .X(_03864_));
 sky130_fd_sc_hd__and2b_1 _07929_ (.A_N(_02747_),
    .B(_03864_),
    .X(_03865_));
 sky130_fd_sc_hd__a211o_1 _07930_ (.A1(_02748_),
    .A2(_03863_),
    .B1(_03865_),
    .C1(_02716_),
    .X(_03866_));
 sky130_fd_sc_hd__mux2_1 _07931_ (.A0(\mem[6][13] ),
    .A1(\mem[7][13] ),
    .S(_02749_),
    .X(_03867_));
 sky130_fd_sc_hd__mux2_1 _07932_ (.A0(\mem[4][13] ),
    .A1(\mem[5][13] ),
    .S(_02428_),
    .X(_03868_));
 sky130_fd_sc_hd__and2b_1 _07933_ (.A_N(_02712_),
    .B(_03868_),
    .X(_03869_));
 sky130_fd_sc_hd__a211o_1 _07934_ (.A1(_02748_),
    .A2(_03867_),
    .B1(_03869_),
    .C1(_02716_),
    .X(_03870_));
 sky130_fd_sc_hd__mux4_1 _07935_ (.A0(\mem[0][13] ),
    .A1(\mem[1][13] ),
    .A2(\mem[2][13] ),
    .A3(\mem[3][13] ),
    .S0(_02693_),
    .S1(_02704_),
    .X(_03871_));
 sky130_fd_sc_hd__o21ba_1 _07936_ (.A1(_02718_),
    .A2(_03871_),
    .B1_N(_02479_),
    .X(_03872_));
 sky130_fd_sc_hd__a32o_1 _07937_ (.A1(_02721_),
    .A2(_03862_),
    .A3(_03866_),
    .B1(_03870_),
    .B2(_03872_),
    .X(_03873_));
 sky130_fd_sc_hd__a221o_1 _07938_ (.A1(_02725_),
    .A2(_03860_),
    .B1(_03873_),
    .B2(_02761_),
    .C1(_02634_),
    .X(_03874_));
 sky130_fd_sc_hd__mux4_1 _07939_ (.A0(\mem[60][13] ),
    .A1(\mem[61][13] ),
    .A2(\mem[62][13] ),
    .A3(\mem[63][13] ),
    .S0(_02698_),
    .S1(_02699_),
    .X(_03875_));
 sky130_fd_sc_hd__mux4_1 _07940_ (.A0(\mem[48][13] ),
    .A1(\mem[49][13] ),
    .A2(\mem[50][13] ),
    .A3(\mem[51][13] ),
    .S0(_02698_),
    .S1(_02748_),
    .X(_03876_));
 sky130_fd_sc_hd__mux4_1 _07941_ (.A0(\mem[52][13] ),
    .A1(\mem[53][13] ),
    .A2(\mem[54][13] ),
    .A3(\mem[55][13] ),
    .S0(_02693_),
    .S1(_02747_),
    .X(_03877_));
 sky130_fd_sc_hd__mux4_1 _07942_ (.A0(\mem[56][13] ),
    .A1(\mem[57][13] ),
    .A2(\mem[58][13] ),
    .A3(\mem[59][13] ),
    .S0(_02693_),
    .S1(_02747_),
    .X(_03878_));
 sky130_fd_sc_hd__o22a_1 _07943_ (.A1(_02702_),
    .A2(_03877_),
    .B1(_03878_),
    .B2(_02707_),
    .X(_03879_));
 sky130_fd_sc_hd__o221a_1 _07944_ (.A1(_02485_),
    .A2(_03875_),
    .B1(_03876_),
    .B2(_02496_),
    .C1(_03879_),
    .X(_03880_));
 sky130_fd_sc_hd__mux4_1 _07945_ (.A0(\mem[36][13] ),
    .A1(\mem[37][13] ),
    .A2(\mem[38][13] ),
    .A3(\mem[39][13] ),
    .S0(_02656_),
    .S1(_02743_),
    .X(_03881_));
 sky130_fd_sc_hd__mux4_1 _07946_ (.A0(\mem[32][13] ),
    .A1(\mem[33][13] ),
    .A2(\mem[34][13] ),
    .A3(\mem[35][13] ),
    .S0(_02681_),
    .S1(_02704_),
    .X(_03882_));
 sky130_fd_sc_hd__a22o_1 _07947_ (.A1(_02677_),
    .A2(_03881_),
    .B1(_03882_),
    .B2(_02652_),
    .X(_03883_));
 sky130_fd_sc_hd__mux4_1 _07948_ (.A0(\mem[44][13] ),
    .A1(\mem[45][13] ),
    .A2(\mem[46][13] ),
    .A3(\mem[47][13] ),
    .S0(_02656_),
    .S1(_02743_),
    .X(_03884_));
 sky130_fd_sc_hd__mux4_1 _07949_ (.A0(\mem[40][13] ),
    .A1(\mem[41][13] ),
    .A2(\mem[42][13] ),
    .A3(\mem[43][13] ),
    .S0(_02645_),
    .S1(_02430_),
    .X(_03885_));
 sky130_fd_sc_hd__or2_1 _07950_ (.A(_02475_),
    .B(_03885_),
    .X(_03886_));
 sky130_fd_sc_hd__o211a_1 _07951_ (.A1(_02472_),
    .A2(_03884_),
    .B1(_03886_),
    .C1(_02721_),
    .X(_03887_));
 sky130_fd_sc_hd__or3_1 _07952_ (.A(_02680_),
    .B(_03883_),
    .C(_03887_),
    .X(_03888_));
 sky130_fd_sc_hd__o211a_1 _07953_ (.A1(_02638_),
    .A2(_03880_),
    .B1(_03888_),
    .C1(_02637_),
    .X(_03889_));
 sky130_fd_sc_hd__o2bb2a_1 _07954_ (.A1_N(_02635_),
    .A2_N(_03846_),
    .B1(_03874_),
    .B2(_03889_),
    .X(_00004_));
 sky130_fd_sc_hd__o21a_1 _07955_ (.A1(\mem[29][14] ),
    .A2(_02515_),
    .B1(_02516_),
    .X(_03890_));
 sky130_fd_sc_hd__or3_1 _07956_ (.A(_02520_),
    .B(_02521_),
    .C(\mem[28][14] ),
    .X(_03891_));
 sky130_fd_sc_hd__o221a_1 _07957_ (.A1(\mem[30][14] ),
    .A2(_02995_),
    .B1(_02519_),
    .B2(\mem[31][14] ),
    .C1(_03891_),
    .X(_03892_));
 sky130_fd_sc_hd__o21a_1 _07958_ (.A1(\mem[16][14] ),
    .A2(_02524_),
    .B1(_02525_),
    .X(_03893_));
 sky130_fd_sc_hd__or3b_1 _07959_ (.A(_02529_),
    .B(\mem[18][14] ),
    .C_N(_02530_),
    .X(_03894_));
 sky130_fd_sc_hd__o221a_1 _07960_ (.A1(\mem[17][14] ),
    .A2(_02899_),
    .B1(_02528_),
    .B2(\mem[19][14] ),
    .C1(_03894_),
    .X(_03895_));
 sky130_fd_sc_hd__a22o_1 _07961_ (.A1(_03890_),
    .A2(_03892_),
    .B1(_03893_),
    .B2(_03895_),
    .X(_03896_));
 sky130_fd_sc_hd__o21a_1 _07962_ (.A1(\mem[24][14] ),
    .A2(_02535_),
    .B1(_02536_),
    .X(_03897_));
 sky130_fd_sc_hd__o22a_1 _07963_ (.A1(\mem[25][14] ),
    .A2(_02538_),
    .B1(_02539_),
    .B2(\mem[27][14] ),
    .X(_03898_));
 sky130_fd_sc_hd__o211a_1 _07964_ (.A1(\mem[26][14] ),
    .A2(_02534_),
    .B1(_03897_),
    .C1(_03898_),
    .X(_03899_));
 sky130_fd_sc_hd__or3_1 _07965_ (.A(_02545_),
    .B(_02546_),
    .C(\mem[20][14] ),
    .X(_03900_));
 sky130_fd_sc_hd__o221a_1 _07966_ (.A1(\mem[22][14] ),
    .A2(_02543_),
    .B1(_02544_),
    .B2(\mem[23][14] ),
    .C1(_03900_),
    .X(_03901_));
 sky130_fd_sc_hd__o211a_1 _07967_ (.A1(\mem[21][14] ),
    .A2(_02542_),
    .B1(_03901_),
    .C1(_02549_),
    .X(_03902_));
 sky130_fd_sc_hd__or4_2 _07968_ (.A(_02993_),
    .B(_03896_),
    .C(_03899_),
    .D(_03902_),
    .X(_03903_));
 sky130_fd_sc_hd__or3_1 _07969_ (.A(_02432_),
    .B(_02433_),
    .C(\mem[12][14] ),
    .X(_03904_));
 sky130_fd_sc_hd__o221a_1 _07970_ (.A1(\mem[14][14] ),
    .A2(_02554_),
    .B1(_03009_),
    .B2(\mem[15][14] ),
    .C1(_03904_),
    .X(_03905_));
 sky130_fd_sc_hd__o211a_1 _07971_ (.A1(\mem[13][14] ),
    .A2(_02553_),
    .B1(_03905_),
    .C1(_02559_),
    .X(_03906_));
 sky130_fd_sc_hd__o21a_1 _07972_ (.A1(\mem[0][14] ),
    .A2(_02562_),
    .B1(_03013_),
    .X(_03907_));
 sky130_fd_sc_hd__o22a_1 _07973_ (.A1(\mem[1][14] ),
    .A2(_02565_),
    .B1(_02914_),
    .B2(\mem[3][14] ),
    .X(_03908_));
 sky130_fd_sc_hd__o211a_1 _07974_ (.A1(\mem[2][14] ),
    .A2(_02561_),
    .B1(_03907_),
    .C1(_03908_),
    .X(_03909_));
 sky130_fd_sc_hd__or2_1 _07975_ (.A(\mem[8][14] ),
    .B(_02917_),
    .X(_03910_));
 sky130_fd_sc_hd__or3b_1 _07976_ (.A(_02574_),
    .B(\mem[10][14] ),
    .C_N(_02575_),
    .X(_03911_));
 sky130_fd_sc_hd__o221a_1 _07977_ (.A1(\mem[9][14] ),
    .A2(_02572_),
    .B1(_02573_),
    .B2(\mem[11][14] ),
    .C1(_03911_),
    .X(_03912_));
 sky130_fd_sc_hd__o21a_1 _07978_ (.A1(\mem[5][14] ),
    .A2(_02578_),
    .B1(_02579_),
    .X(_03913_));
 sky130_fd_sc_hd__or3_1 _07979_ (.A(_02583_),
    .B(_02584_),
    .C(\mem[4][14] ),
    .X(_03914_));
 sky130_fd_sc_hd__o221a_1 _07980_ (.A1(\mem[6][14] ),
    .A2(_02581_),
    .B1(_02582_),
    .B2(\mem[7][14] ),
    .C1(_03914_),
    .X(_03915_));
 sky130_fd_sc_hd__a32o_1 _07981_ (.A1(_02569_),
    .A2(_03910_),
    .A3(_03912_),
    .B1(_03913_),
    .B2(_03915_),
    .X(_03916_));
 sky130_fd_sc_hd__or4_1 _07982_ (.A(_02552_),
    .B(_03906_),
    .C(_03909_),
    .D(_03916_),
    .X(_03917_));
 sky130_fd_sc_hd__mux4_1 _07983_ (.A0(\mem[32][14] ),
    .A1(\mem[33][14] ),
    .A2(\mem[34][14] ),
    .A3(\mem[35][14] ),
    .S0(_02590_),
    .S1(_02926_),
    .X(_03918_));
 sky130_fd_sc_hd__mux4_1 _07984_ (.A0(\mem[36][14] ),
    .A1(\mem[37][14] ),
    .A2(\mem[38][14] ),
    .A3(\mem[39][14] ),
    .S0(_02928_),
    .S1(_02929_),
    .X(_03919_));
 sky130_fd_sc_hd__a22o_1 _07985_ (.A1(_02456_),
    .A2(_03918_),
    .B1(_03919_),
    .B2(_02465_),
    .X(_03920_));
 sky130_fd_sc_hd__mux4_1 _07986_ (.A0(\mem[44][14] ),
    .A1(\mem[45][14] ),
    .A2(\mem[46][14] ),
    .A3(\mem[47][14] ),
    .S0(_02600_),
    .S1(_02601_),
    .X(_03921_));
 sky130_fd_sc_hd__mux4_1 _07987_ (.A0(\mem[40][14] ),
    .A1(\mem[41][14] ),
    .A2(\mem[42][14] ),
    .A3(\mem[43][14] ),
    .S0(_02604_),
    .S1(_02605_),
    .X(_03922_));
 sky130_fd_sc_hd__or2_1 _07988_ (.A(_02603_),
    .B(_03922_),
    .X(_03923_));
 sky130_fd_sc_hd__o211a_1 _07989_ (.A1(_02599_),
    .A2(_03921_),
    .B1(_03923_),
    .C1(_02608_),
    .X(_03924_));
 sky130_fd_sc_hd__or3_4 _07990_ (.A(_02589_),
    .B(_03920_),
    .C(_03924_),
    .X(_03925_));
 sky130_fd_sc_hd__mux4_1 _07991_ (.A0(\mem[60][14] ),
    .A1(\mem[61][14] ),
    .A2(\mem[62][14] ),
    .A3(\mem[63][14] ),
    .S0(_02613_),
    .S1(_02614_),
    .X(_03926_));
 sky130_fd_sc_hd__mux4_1 _07992_ (.A0(\mem[48][14] ),
    .A1(\mem[49][14] ),
    .A2(\mem[50][14] ),
    .A3(\mem[51][14] ),
    .S0(_02616_),
    .S1(_02746_),
    .X(_03927_));
 sky130_fd_sc_hd__mux4_1 _07993_ (.A0(\mem[52][14] ),
    .A1(\mem[53][14] ),
    .A2(\mem[54][14] ),
    .A3(\mem[55][14] ),
    .S0(_02622_),
    .S1(_02623_),
    .X(_03928_));
 sky130_fd_sc_hd__mux4_1 _07994_ (.A0(\mem[56][14] ),
    .A1(\mem[57][14] ),
    .A2(\mem[58][14] ),
    .A3(\mem[59][14] ),
    .S0(_02625_),
    .S1(_02626_),
    .X(_03929_));
 sky130_fd_sc_hd__o22a_1 _07995_ (.A1(_02621_),
    .A2(_03928_),
    .B1(_03929_),
    .B2(_02628_),
    .X(_03930_));
 sky130_fd_sc_hd__o221a_1 _07996_ (.A1(_03033_),
    .A2(_03926_),
    .B1(_03927_),
    .B2(_02620_),
    .C1(_03930_),
    .X(_03931_));
 sky130_fd_sc_hd__o21a_1 _07997_ (.A1(_02611_),
    .A2(_03931_),
    .B1(_02631_),
    .X(_03932_));
 sky130_fd_sc_hd__a32o_1 _07998_ (.A1(_02513_),
    .A2(_03903_),
    .A3(_03917_),
    .B1(_03925_),
    .B2(_03932_),
    .X(_03933_));
 sky130_fd_sc_hd__o21a_1 _07999_ (.A1(\mem[93][14] ),
    .A2(_03042_),
    .B1(_02365_),
    .X(_03934_));
 sky130_fd_sc_hd__or3_1 _08000_ (.A(_02466_),
    .B(_02459_),
    .C(\mem[92][14] ),
    .X(_03935_));
 sky130_fd_sc_hd__o221a_1 _08001_ (.A1(\mem[94][14] ),
    .A2(_02518_),
    .B1(_02400_),
    .B2(\mem[95][14] ),
    .C1(_03935_),
    .X(_03936_));
 sky130_fd_sc_hd__o21a_1 _08002_ (.A1(\mem[80][14] ),
    .A2(_02812_),
    .B1(_02454_),
    .X(_03937_));
 sky130_fd_sc_hd__or3b_1 _08003_ (.A(_02670_),
    .B(\mem[82][14] ),
    .C_N(_02375_),
    .X(_03938_));
 sky130_fd_sc_hd__o221a_1 _08004_ (.A1(\mem[81][14] ),
    .A2(_02404_),
    .B1(_02424_),
    .B2(\mem[83][14] ),
    .C1(_03938_),
    .X(_03939_));
 sky130_fd_sc_hd__a22o_1 _08005_ (.A1(_03934_),
    .A2(_03936_),
    .B1(_03937_),
    .B2(_03939_),
    .X(_03940_));
 sky130_fd_sc_hd__o21a_1 _08006_ (.A1(\mem[88][14] ),
    .A2(_02380_),
    .B1(_02396_),
    .X(_03941_));
 sky130_fd_sc_hd__o22a_1 _08007_ (.A1(\mem[89][14] ),
    .A2(_02363_),
    .B1(_03231_),
    .B2(\mem[91][14] ),
    .X(_03942_));
 sky130_fd_sc_hd__o211a_1 _08008_ (.A1(\mem[90][14] ),
    .A2(_02660_),
    .B1(_03941_),
    .C1(_03942_),
    .X(_03943_));
 sky130_fd_sc_hd__or3_1 _08009_ (.A(_02486_),
    .B(_03224_),
    .C(\mem[84][14] ),
    .X(_03944_));
 sky130_fd_sc_hd__o221a_1 _08010_ (.A1(\mem[86][14] ),
    .A2(_02956_),
    .B1(_02664_),
    .B2(\mem[87][14] ),
    .C1(_03944_),
    .X(_03945_));
 sky130_fd_sc_hd__o211a_1 _08011_ (.A1(\mem[85][14] ),
    .A2(_02955_),
    .B1(_03945_),
    .C1(_02464_),
    .X(_03946_));
 sky130_fd_sc_hd__or4_2 _08012_ (.A(_02514_),
    .B(_03940_),
    .C(_03943_),
    .D(_03946_),
    .X(_03947_));
 sky130_fd_sc_hd__or3_1 _08013_ (.A(_02556_),
    .B(_02389_),
    .C(\mem[76][14] ),
    .X(_03948_));
 sky130_fd_sc_hd__o221a_1 _08014_ (.A1(\mem[78][14] ),
    .A2(_02370_),
    .B1(_02555_),
    .B2(\mem[79][14] ),
    .C1(_03948_),
    .X(_03949_));
 sky130_fd_sc_hd__o211a_1 _08015_ (.A1(\mem[77][14] ),
    .A2(_02639_),
    .B1(_03949_),
    .C1(_02422_),
    .X(_03950_));
 sky130_fd_sc_hd__o21a_1 _08016_ (.A1(\mem[64][14] ),
    .A2(_02395_),
    .B1(_02563_),
    .X(_03951_));
 sky130_fd_sc_hd__o22a_1 _08017_ (.A1(\mem[65][14] ),
    .A2(_02399_),
    .B1(_02401_),
    .B2(\mem[67][14] ),
    .X(_03952_));
 sky130_fd_sc_hd__o211a_1 _08018_ (.A1(\mem[66][14] ),
    .A2(_02394_),
    .B1(_03951_),
    .C1(_03952_),
    .X(_03953_));
 sky130_fd_sc_hd__or2_1 _08019_ (.A(\mem[72][14] ),
    .B(_02379_),
    .X(_03954_));
 sky130_fd_sc_hd__or3b_1 _08020_ (.A(_02802_),
    .B(\mem[74][14] ),
    .C_N(_02803_),
    .X(_03955_));
 sky130_fd_sc_hd__o221a_1 _08021_ (.A1(\mem[73][14] ),
    .A2(_02385_),
    .B1(_02801_),
    .B2(\mem[75][14] ),
    .C1(_03955_),
    .X(_03956_));
 sky130_fd_sc_hd__o21a_1 _08022_ (.A1(\mem[69][14] ),
    .A2(_02405_),
    .B1(_02463_),
    .X(_03957_));
 sky130_fd_sc_hd__or3_1 _08023_ (.A(_02411_),
    .B(_02868_),
    .C(\mem[68][14] ),
    .X(_03958_));
 sky130_fd_sc_hd__o221a_1 _08024_ (.A1(\mem[70][14] ),
    .A2(_02407_),
    .B1(_02409_),
    .B2(\mem[71][14] ),
    .C1(_03958_),
    .X(_03959_));
 sky130_fd_sc_hd__a32o_1 _08025_ (.A1(_02439_),
    .A2(_03954_),
    .A3(_03956_),
    .B1(_03957_),
    .B2(_03959_),
    .X(_03960_));
 sky130_fd_sc_hd__or4_1 _08026_ (.A(_02420_),
    .B(_03950_),
    .C(_03953_),
    .D(_03960_),
    .X(_03961_));
 sky130_fd_sc_hd__mux4_1 _08027_ (.A0(\mem[96][14] ),
    .A1(\mem[97][14] ),
    .A2(\mem[98][14] ),
    .A3(\mem[99][14] ),
    .S0(_02645_),
    .S1(_02430_),
    .X(_03962_));
 sky130_fd_sc_hd__mux4_1 _08028_ (.A0(\mem[100][14] ),
    .A1(\mem[101][14] ),
    .A2(\mem[102][14] ),
    .A3(\mem[103][14] ),
    .S0(_02467_),
    .S1(_02468_),
    .X(_03963_));
 sky130_fd_sc_hd__a22o_1 _08029_ (.A1(_02651_),
    .A2(_03962_),
    .B1(_03963_),
    .B2(_02825_),
    .X(_03964_));
 sky130_fd_sc_hd__mux4_1 _08030_ (.A0(\mem[108][14] ),
    .A1(\mem[109][14] ),
    .A2(\mem[110][14] ),
    .A3(\mem[111][14] ),
    .S0(_02458_),
    .S1(_02461_),
    .X(_03965_));
 sky130_fd_sc_hd__mux4_1 _08031_ (.A0(\mem[104][14] ),
    .A1(\mem[105][14] ),
    .A2(\mem[106][14] ),
    .A3(\mem[107][14] ),
    .S0(_02501_),
    .S1(_02877_),
    .X(_03966_));
 sky130_fd_sc_hd__or2_1 _08032_ (.A(_02474_),
    .B(_03966_),
    .X(_03967_));
 sky130_fd_sc_hd__o211a_1 _08033_ (.A1(_02598_),
    .A2(_03965_),
    .B1(_03967_),
    .C1(_02478_),
    .X(_03968_));
 sky130_fd_sc_hd__or3_2 _08034_ (.A(_02421_),
    .B(_03964_),
    .C(_03968_),
    .X(_03969_));
 sky130_fd_sc_hd__mux4_1 _08035_ (.A0(\mem[124][14] ),
    .A1(\mem[125][14] ),
    .A2(\mem[126][14] ),
    .A3(\mem[127][14] ),
    .S0(_02671_),
    .S1(_02703_),
    .X(_03970_));
 sky130_fd_sc_hd__mux4_1 _08036_ (.A0(\mem[112][14] ),
    .A1(\mem[113][14] ),
    .A2(\mem[114][14] ),
    .A3(\mem[115][14] ),
    .S0(_02726_),
    .S1(_02618_),
    .X(_03971_));
 sky130_fd_sc_hd__mux4_1 _08037_ (.A0(\mem[116][14] ),
    .A1(\mem[117][14] ),
    .A2(\mem[118][14] ),
    .A3(\mem[119][14] ),
    .S0(_02985_),
    .S1(_02617_),
    .X(_03972_));
 sky130_fd_sc_hd__mux4_1 _08038_ (.A0(\mem[120][14] ),
    .A1(\mem[121][14] ),
    .A2(\mem[122][14] ),
    .A3(\mem[123][14] ),
    .S0(_02887_),
    .S1(_02499_),
    .X(_03973_));
 sky130_fd_sc_hd__o22a_1 _08039_ (.A1(_02885_),
    .A2(_03972_),
    .B1(_03973_),
    .B2(_02889_),
    .X(_03974_));
 sky130_fd_sc_hd__o221a_2 _08040_ (.A1(_02612_),
    .A2(_03970_),
    .B1(_03971_),
    .B2(_02884_),
    .C1(_03974_),
    .X(_03975_));
 sky130_fd_sc_hd__o21a_1 _08041_ (.A1(_02358_),
    .A2(_03975_),
    .B1(_02509_),
    .X(_03976_));
 sky130_fd_sc_hd__a32o_1 _08042_ (.A1(_02355_),
    .A2(_03947_),
    .A3(_03961_),
    .B1(_03969_),
    .B2(_03976_),
    .X(_03977_));
 sky130_fd_sc_hd__mux2_1 _08043_ (.A0(_03933_),
    .A1(_03977_),
    .S(_02634_),
    .X(_03978_));
 sky130_fd_sc_hd__clkbuf_1 _08044_ (.A(_03978_),
    .X(_00005_));
 sky130_fd_sc_hd__o21a_1 _08045_ (.A1(\mem[29][15] ),
    .A2(_02515_),
    .B1(_02516_),
    .X(_03979_));
 sky130_fd_sc_hd__or3_1 _08046_ (.A(_02520_),
    .B(_02521_),
    .C(\mem[28][15] ),
    .X(_03980_));
 sky130_fd_sc_hd__o221a_1 _08047_ (.A1(\mem[30][15] ),
    .A2(_02995_),
    .B1(_02519_),
    .B2(\mem[31][15] ),
    .C1(_03980_),
    .X(_03981_));
 sky130_fd_sc_hd__o21a_1 _08048_ (.A1(\mem[16][15] ),
    .A2(_02524_),
    .B1(_02525_),
    .X(_03982_));
 sky130_fd_sc_hd__or3b_1 _08049_ (.A(_02529_),
    .B(\mem[18][15] ),
    .C_N(_02530_),
    .X(_03983_));
 sky130_fd_sc_hd__o221a_1 _08050_ (.A1(\mem[17][15] ),
    .A2(_02527_),
    .B1(_02528_),
    .B2(\mem[19][15] ),
    .C1(_03983_),
    .X(_03984_));
 sky130_fd_sc_hd__a22o_1 _08051_ (.A1(_03979_),
    .A2(_03981_),
    .B1(_03982_),
    .B2(_03984_),
    .X(_03985_));
 sky130_fd_sc_hd__o21a_1 _08052_ (.A1(\mem[24][15] ),
    .A2(_02535_),
    .B1(_02536_),
    .X(_03986_));
 sky130_fd_sc_hd__o22a_1 _08053_ (.A1(\mem[25][15] ),
    .A2(_02538_),
    .B1(_02539_),
    .B2(\mem[27][15] ),
    .X(_03987_));
 sky130_fd_sc_hd__o211a_1 _08054_ (.A1(\mem[26][15] ),
    .A2(_02534_),
    .B1(_03986_),
    .C1(_03987_),
    .X(_03988_));
 sky130_fd_sc_hd__or3_1 _08055_ (.A(_02545_),
    .B(_02546_),
    .C(\mem[20][15] ),
    .X(_03989_));
 sky130_fd_sc_hd__o221a_1 _08056_ (.A1(\mem[22][15] ),
    .A2(_02543_),
    .B1(_02544_),
    .B2(\mem[23][15] ),
    .C1(_03989_),
    .X(_03990_));
 sky130_fd_sc_hd__o211a_1 _08057_ (.A1(\mem[21][15] ),
    .A2(_02542_),
    .B1(_03990_),
    .C1(_02549_),
    .X(_03991_));
 sky130_fd_sc_hd__or4_2 _08058_ (.A(_02993_),
    .B(_03985_),
    .C(_03988_),
    .D(_03991_),
    .X(_03992_));
 sky130_fd_sc_hd__or3_1 _08059_ (.A(_02432_),
    .B(_02433_),
    .C(\mem[12][15] ),
    .X(_03993_));
 sky130_fd_sc_hd__o221a_1 _08060_ (.A1(\mem[14][15] ),
    .A2(_02554_),
    .B1(_03009_),
    .B2(\mem[15][15] ),
    .C1(_03993_),
    .X(_03994_));
 sky130_fd_sc_hd__o211a_1 _08061_ (.A1(\mem[13][15] ),
    .A2(_02553_),
    .B1(_03994_),
    .C1(_02559_),
    .X(_03995_));
 sky130_fd_sc_hd__o21a_1 _08062_ (.A1(\mem[0][15] ),
    .A2(_02562_),
    .B1(_03013_),
    .X(_03996_));
 sky130_fd_sc_hd__o22a_1 _08063_ (.A1(\mem[1][15] ),
    .A2(_02565_),
    .B1(_02566_),
    .B2(\mem[3][15] ),
    .X(_03997_));
 sky130_fd_sc_hd__o211a_1 _08064_ (.A1(\mem[2][15] ),
    .A2(_02561_),
    .B1(_03996_),
    .C1(_03997_),
    .X(_03998_));
 sky130_fd_sc_hd__or2_1 _08065_ (.A(\mem[8][15] ),
    .B(_02570_),
    .X(_03999_));
 sky130_fd_sc_hd__or3b_1 _08066_ (.A(_02574_),
    .B(\mem[10][15] ),
    .C_N(_02575_),
    .X(_04000_));
 sky130_fd_sc_hd__o221a_1 _08067_ (.A1(\mem[9][15] ),
    .A2(_02572_),
    .B1(_02573_),
    .B2(\mem[11][15] ),
    .C1(_04000_),
    .X(_04001_));
 sky130_fd_sc_hd__o21a_1 _08068_ (.A1(\mem[5][15] ),
    .A2(_02578_),
    .B1(_02579_),
    .X(_04002_));
 sky130_fd_sc_hd__or3_1 _08069_ (.A(_02583_),
    .B(_02584_),
    .C(\mem[4][15] ),
    .X(_04003_));
 sky130_fd_sc_hd__o221a_1 _08070_ (.A1(\mem[6][15] ),
    .A2(_02581_),
    .B1(_02582_),
    .B2(\mem[7][15] ),
    .C1(_04003_),
    .X(_04004_));
 sky130_fd_sc_hd__a32o_2 _08071_ (.A1(_02569_),
    .A2(_03999_),
    .A3(_04001_),
    .B1(_04002_),
    .B2(_04004_),
    .X(_04005_));
 sky130_fd_sc_hd__or4_1 _08072_ (.A(_02552_),
    .B(_03995_),
    .C(_03998_),
    .D(_04005_),
    .X(_04006_));
 sky130_fd_sc_hd__mux4_1 _08073_ (.A0(\mem[32][15] ),
    .A1(\mem[33][15] ),
    .A2(\mem[34][15] ),
    .A3(\mem[35][15] ),
    .S0(_02590_),
    .S1(_02591_),
    .X(_04007_));
 sky130_fd_sc_hd__mux4_1 _08074_ (.A0(\mem[36][15] ),
    .A1(\mem[37][15] ),
    .A2(\mem[38][15] ),
    .A3(\mem[39][15] ),
    .S0(_02593_),
    .S1(_02594_),
    .X(_04008_));
 sky130_fd_sc_hd__a22o_1 _08075_ (.A1(_02456_),
    .A2(_04007_),
    .B1(_04008_),
    .B2(_02465_),
    .X(_04009_));
 sky130_fd_sc_hd__mux4_1 _08076_ (.A0(\mem[44][15] ),
    .A1(\mem[45][15] ),
    .A2(\mem[46][15] ),
    .A3(\mem[47][15] ),
    .S0(_02600_),
    .S1(_02601_),
    .X(_04010_));
 sky130_fd_sc_hd__mux4_1 _08077_ (.A0(\mem[40][15] ),
    .A1(\mem[41][15] ),
    .A2(\mem[42][15] ),
    .A3(\mem[43][15] ),
    .S0(_02604_),
    .S1(_02605_),
    .X(_04011_));
 sky130_fd_sc_hd__or2_1 _08078_ (.A(_02603_),
    .B(_04011_),
    .X(_04012_));
 sky130_fd_sc_hd__o211a_1 _08079_ (.A1(_02599_),
    .A2(_04010_),
    .B1(_04012_),
    .C1(_02608_),
    .X(_04013_));
 sky130_fd_sc_hd__or3_2 _08080_ (.A(_02589_),
    .B(_04009_),
    .C(_04013_),
    .X(_04014_));
 sky130_fd_sc_hd__mux4_1 _08081_ (.A0(\mem[60][15] ),
    .A1(\mem[61][15] ),
    .A2(\mem[62][15] ),
    .A3(\mem[63][15] ),
    .S0(_02613_),
    .S1(_02614_),
    .X(_04015_));
 sky130_fd_sc_hd__mux4_1 _08082_ (.A0(\mem[48][15] ),
    .A1(\mem[49][15] ),
    .A2(\mem[50][15] ),
    .A3(\mem[51][15] ),
    .S0(_02616_),
    .S1(_02746_),
    .X(_04016_));
 sky130_fd_sc_hd__mux4_1 _08083_ (.A0(\mem[52][15] ),
    .A1(\mem[53][15] ),
    .A2(\mem[54][15] ),
    .A3(\mem[55][15] ),
    .S0(_02622_),
    .S1(_02623_),
    .X(_04017_));
 sky130_fd_sc_hd__mux4_1 _08084_ (.A0(\mem[56][15] ),
    .A1(\mem[57][15] ),
    .A2(\mem[58][15] ),
    .A3(\mem[59][15] ),
    .S0(_02625_),
    .S1(_02626_),
    .X(_04018_));
 sky130_fd_sc_hd__o22a_1 _08085_ (.A1(_02621_),
    .A2(_04017_),
    .B1(_04018_),
    .B2(_02628_),
    .X(_04019_));
 sky130_fd_sc_hd__o221a_1 _08086_ (.A1(_03033_),
    .A2(_04015_),
    .B1(_04016_),
    .B2(_02620_),
    .C1(_04019_),
    .X(_04020_));
 sky130_fd_sc_hd__o21a_1 _08087_ (.A1(_02611_),
    .A2(_04020_),
    .B1(_02631_),
    .X(_04021_));
 sky130_fd_sc_hd__a32o_1 _08088_ (.A1(_02513_),
    .A2(_03992_),
    .A3(_04006_),
    .B1(_04014_),
    .B2(_04021_),
    .X(_04022_));
 sky130_fd_sc_hd__o21a_1 _08089_ (.A1(\mem[93][15] ),
    .A2(_03042_),
    .B1(_02365_),
    .X(_04023_));
 sky130_fd_sc_hd__or3_1 _08090_ (.A(_02466_),
    .B(_02459_),
    .C(\mem[92][15] ),
    .X(_04024_));
 sky130_fd_sc_hd__o221a_1 _08091_ (.A1(\mem[94][15] ),
    .A2(_02369_),
    .B1(_02400_),
    .B2(\mem[95][15] ),
    .C1(_04024_),
    .X(_04025_));
 sky130_fd_sc_hd__o21a_1 _08092_ (.A1(\mem[80][15] ),
    .A2(_02812_),
    .B1(_02454_),
    .X(_04026_));
 sky130_fd_sc_hd__or3b_1 _08093_ (.A(_02670_),
    .B(\mem[82][15] ),
    .C_N(_02375_),
    .X(_04027_));
 sky130_fd_sc_hd__o221a_1 _08094_ (.A1(\mem[81][15] ),
    .A2(_02404_),
    .B1(_02424_),
    .B2(\mem[83][15] ),
    .C1(_04027_),
    .X(_04028_));
 sky130_fd_sc_hd__a22o_1 _08095_ (.A1(_04023_),
    .A2(_04025_),
    .B1(_04026_),
    .B2(_04028_),
    .X(_04029_));
 sky130_fd_sc_hd__o21a_1 _08096_ (.A1(\mem[88][15] ),
    .A2(_02380_),
    .B1(_02396_),
    .X(_04030_));
 sky130_fd_sc_hd__o22a_1 _08097_ (.A1(\mem[89][15] ),
    .A2(_02363_),
    .B1(_03231_),
    .B2(\mem[91][15] ),
    .X(_04031_));
 sky130_fd_sc_hd__o211a_1 _08098_ (.A1(\mem[90][15] ),
    .A2(_02660_),
    .B1(_04030_),
    .C1(_04031_),
    .X(_04032_));
 sky130_fd_sc_hd__or3_1 _08099_ (.A(_02486_),
    .B(_03224_),
    .C(\mem[84][15] ),
    .X(_04033_));
 sky130_fd_sc_hd__o221a_1 _08100_ (.A1(\mem[86][15] ),
    .A2(_02956_),
    .B1(_02664_),
    .B2(\mem[87][15] ),
    .C1(_04033_),
    .X(_04034_));
 sky130_fd_sc_hd__o211a_1 _08101_ (.A1(\mem[85][15] ),
    .A2(_02955_),
    .B1(_04034_),
    .C1(_02464_),
    .X(_04035_));
 sky130_fd_sc_hd__or4_2 _08102_ (.A(_02357_),
    .B(_04029_),
    .C(_04032_),
    .D(_04035_),
    .X(_04036_));
 sky130_fd_sc_hd__or3_1 _08103_ (.A(_02387_),
    .B(_02389_),
    .C(\mem[76][15] ),
    .X(_04037_));
 sky130_fd_sc_hd__o221a_1 _08104_ (.A1(\mem[78][15] ),
    .A2(_02370_),
    .B1(_02386_),
    .B2(\mem[79][15] ),
    .C1(_04037_),
    .X(_04038_));
 sky130_fd_sc_hd__o211a_1 _08105_ (.A1(\mem[77][15] ),
    .A2(_02639_),
    .B1(_04038_),
    .C1(_02422_),
    .X(_04039_));
 sky130_fd_sc_hd__o21a_1 _08106_ (.A1(\mem[64][15] ),
    .A2(_02395_),
    .B1(_02383_),
    .X(_04040_));
 sky130_fd_sc_hd__o22a_1 _08107_ (.A1(\mem[65][15] ),
    .A2(_02399_),
    .B1(_02401_),
    .B2(\mem[67][15] ),
    .X(_04041_));
 sky130_fd_sc_hd__o211a_1 _08108_ (.A1(\mem[66][15] ),
    .A2(_02394_),
    .B1(_04040_),
    .C1(_04041_),
    .X(_04042_));
 sky130_fd_sc_hd__or2_1 _08109_ (.A(\mem[72][15] ),
    .B(_02379_),
    .X(_04043_));
 sky130_fd_sc_hd__or3b_1 _08110_ (.A(_02802_),
    .B(\mem[74][15] ),
    .C_N(_02803_),
    .X(_04044_));
 sky130_fd_sc_hd__o221a_1 _08111_ (.A1(\mem[73][15] ),
    .A2(_02385_),
    .B1(_02801_),
    .B2(\mem[75][15] ),
    .C1(_04044_),
    .X(_04045_));
 sky130_fd_sc_hd__o21a_1 _08112_ (.A1(\mem[69][15] ),
    .A2(_02405_),
    .B1(_02463_),
    .X(_04046_));
 sky130_fd_sc_hd__or3_1 _08113_ (.A(_02411_),
    .B(_02868_),
    .C(\mem[68][15] ),
    .X(_04047_));
 sky130_fd_sc_hd__o221a_1 _08114_ (.A1(\mem[70][15] ),
    .A2(_02407_),
    .B1(_02409_),
    .B2(\mem[71][15] ),
    .C1(_04047_),
    .X(_04048_));
 sky130_fd_sc_hd__a32o_1 _08115_ (.A1(_02439_),
    .A2(_04043_),
    .A3(_04045_),
    .B1(_04046_),
    .B2(_04048_),
    .X(_04049_));
 sky130_fd_sc_hd__or4_1 _08116_ (.A(_02420_),
    .B(_04039_),
    .C(_04042_),
    .D(_04049_),
    .X(_04050_));
 sky130_fd_sc_hd__mux4_1 _08117_ (.A0(\mem[100][15] ),
    .A1(\mem[101][15] ),
    .A2(\mem[102][15] ),
    .A3(\mem[103][15] ),
    .S0(_02645_),
    .S1(_02430_),
    .X(_04051_));
 sky130_fd_sc_hd__mux4_1 _08118_ (.A0(\mem[96][15] ),
    .A1(\mem[97][15] ),
    .A2(\mem[98][15] ),
    .A3(\mem[99][15] ),
    .S0(_02467_),
    .S1(_02468_),
    .X(_04052_));
 sky130_fd_sc_hd__a22o_1 _08119_ (.A1(_02450_),
    .A2(_04051_),
    .B1(_04052_),
    .B2(_02456_),
    .X(_04053_));
 sky130_fd_sc_hd__mux4_1 _08120_ (.A0(\mem[108][15] ),
    .A1(\mem[109][15] ),
    .A2(\mem[110][15] ),
    .A3(\mem[111][15] ),
    .S0(_02458_),
    .S1(_02461_),
    .X(_04054_));
 sky130_fd_sc_hd__mux4_1 _08121_ (.A0(\mem[104][15] ),
    .A1(\mem[105][15] ),
    .A2(\mem[106][15] ),
    .A3(\mem[107][15] ),
    .S0(_02501_),
    .S1(_02877_),
    .X(_04055_));
 sky130_fd_sc_hd__or2_1 _08122_ (.A(_02474_),
    .B(_04055_),
    .X(_04056_));
 sky130_fd_sc_hd__o211a_1 _08123_ (.A1(_02598_),
    .A2(_04054_),
    .B1(_04056_),
    .C1(_02478_),
    .X(_04057_));
 sky130_fd_sc_hd__or3_2 _08124_ (.A(_02421_),
    .B(_04053_),
    .C(_04057_),
    .X(_04058_));
 sky130_fd_sc_hd__buf_8 _08125_ (.A(_02483_),
    .X(_04059_));
 sky130_fd_sc_hd__mux4_1 _08126_ (.A0(\mem[124][15] ),
    .A1(\mem[125][15] ),
    .A2(\mem[126][15] ),
    .A3(\mem[127][15] ),
    .S0(_02671_),
    .S1(_02703_),
    .X(_04060_));
 sky130_fd_sc_hd__mux4_1 _08127_ (.A0(\mem[112][15] ),
    .A1(\mem[113][15] ),
    .A2(\mem[114][15] ),
    .A3(\mem[115][15] ),
    .S0(_02726_),
    .S1(_02489_),
    .X(_04061_));
 sky130_fd_sc_hd__mux4_1 _08128_ (.A0(\mem[116][15] ),
    .A1(\mem[117][15] ),
    .A2(\mem[118][15] ),
    .A3(\mem[119][15] ),
    .S0(_02985_),
    .S1(_02617_),
    .X(_04062_));
 sky130_fd_sc_hd__mux4_1 _08129_ (.A0(\mem[120][15] ),
    .A1(\mem[121][15] ),
    .A2(\mem[122][15] ),
    .A3(\mem[123][15] ),
    .S0(_02887_),
    .S1(_02499_),
    .X(_04063_));
 sky130_fd_sc_hd__o22a_1 _08130_ (.A1(_02885_),
    .A2(_04062_),
    .B1(_04063_),
    .B2(_02889_),
    .X(_04064_));
 sky130_fd_sc_hd__o221a_2 _08131_ (.A1(_04059_),
    .A2(_04060_),
    .B1(_04061_),
    .B2(_02884_),
    .C1(_04064_),
    .X(_04065_));
 sky130_fd_sc_hd__o21a_1 _08132_ (.A1(_02358_),
    .A2(_04065_),
    .B1(_02509_),
    .X(_04066_));
 sky130_fd_sc_hd__a32o_1 _08133_ (.A1(_02355_),
    .A2(_04036_),
    .A3(_04050_),
    .B1(_04058_),
    .B2(_04066_),
    .X(_04067_));
 sky130_fd_sc_hd__mux2_1 _08134_ (.A0(_04022_),
    .A1(_04067_),
    .S(_02634_),
    .X(_04068_));
 sky130_fd_sc_hd__clkbuf_1 _08135_ (.A(_04068_),
    .X(_00006_));
 sky130_fd_sc_hd__buf_8 _08136_ (.A(net8),
    .X(_04069_));
 sky130_fd_sc_hd__buf_6 _08137_ (.A(_04069_),
    .X(_04070_));
 sky130_fd_sc_hd__or2_1 _08138_ (.A(_02495_),
    .B(_02639_),
    .X(_04071_));
 sky130_fd_sc_hd__buf_12 _08139_ (.A(_04071_),
    .X(_04072_));
 sky130_fd_sc_hd__nand2_1 _08140_ (.A(net5),
    .B(net6),
    .Y(_04073_));
 sky130_fd_sc_hd__or2b_1 _08141_ (.A(net7),
    .B_N(net24),
    .X(_04074_));
 sky130_fd_sc_hd__or2_4 _08142_ (.A(_04073_),
    .B(_04074_),
    .X(_04075_));
 sky130_fd_sc_hd__buf_6 _08143_ (.A(_04075_),
    .X(_04076_));
 sky130_fd_sc_hd__nor2_4 _08144_ (.A(_04072_),
    .B(_04076_),
    .Y(_04077_));
 sky130_fd_sc_hd__clkbuf_4 _08145_ (.A(_04077_),
    .X(_04078_));
 sky130_fd_sc_hd__mux2_1 _08146_ (.A0(net2082),
    .A1(_04070_),
    .S(_04078_),
    .X(_04079_));
 sky130_fd_sc_hd__clkbuf_1 _08147_ (.A(_04079_),
    .X(_01505_));
 sky130_fd_sc_hd__buf_6 _08148_ (.A(net15),
    .X(_04080_));
 sky130_fd_sc_hd__buf_4 _08149_ (.A(_04080_),
    .X(_04081_));
 sky130_fd_sc_hd__mux2_1 _08150_ (.A0(net2064),
    .A1(_04081_),
    .S(_04078_),
    .X(_04082_));
 sky130_fd_sc_hd__clkbuf_1 _08151_ (.A(_04082_),
    .X(_01506_));
 sky130_fd_sc_hd__clkbuf_16 _08152_ (.A(net16),
    .X(_04083_));
 sky130_fd_sc_hd__buf_6 _08153_ (.A(_04083_),
    .X(_04084_));
 sky130_fd_sc_hd__mux2_1 _08154_ (.A0(net2084),
    .A1(_04084_),
    .S(_04078_),
    .X(_04085_));
 sky130_fd_sc_hd__clkbuf_1 _08155_ (.A(_04085_),
    .X(_01507_));
 sky130_fd_sc_hd__buf_8 _08156_ (.A(net17),
    .X(_04086_));
 sky130_fd_sc_hd__buf_6 _08157_ (.A(_04086_),
    .X(_04087_));
 sky130_fd_sc_hd__mux2_1 _08158_ (.A0(net2085),
    .A1(_04087_),
    .S(_04078_),
    .X(_04088_));
 sky130_fd_sc_hd__clkbuf_1 _08159_ (.A(_04088_),
    .X(_01508_));
 sky130_fd_sc_hd__buf_8 _08160_ (.A(net18),
    .X(_04089_));
 sky130_fd_sc_hd__buf_6 _08161_ (.A(_04089_),
    .X(_04090_));
 sky130_fd_sc_hd__mux2_1 _08162_ (.A0(net2088),
    .A1(_04090_),
    .S(_04078_),
    .X(_04091_));
 sky130_fd_sc_hd__clkbuf_1 _08163_ (.A(_04091_),
    .X(_01509_));
 sky130_fd_sc_hd__buf_6 _08164_ (.A(net19),
    .X(_04092_));
 sky130_fd_sc_hd__buf_4 _08165_ (.A(_04092_),
    .X(_04093_));
 sky130_fd_sc_hd__mux2_1 _08166_ (.A0(net2070),
    .A1(_04093_),
    .S(_04078_),
    .X(_04094_));
 sky130_fd_sc_hd__clkbuf_1 _08167_ (.A(_04094_),
    .X(_01510_));
 sky130_fd_sc_hd__buf_6 _08168_ (.A(net20),
    .X(_04095_));
 sky130_fd_sc_hd__buf_6 _08169_ (.A(_04095_),
    .X(_04096_));
 sky130_fd_sc_hd__mux2_1 _08170_ (.A0(net2077),
    .A1(_04096_),
    .S(_04078_),
    .X(_04097_));
 sky130_fd_sc_hd__clkbuf_1 _08171_ (.A(_04097_),
    .X(_01511_));
 sky130_fd_sc_hd__buf_8 _08172_ (.A(net21),
    .X(_04098_));
 sky130_fd_sc_hd__buf_6 _08173_ (.A(_04098_),
    .X(_04099_));
 sky130_fd_sc_hd__mux2_1 _08174_ (.A0(net2086),
    .A1(_04099_),
    .S(_04078_),
    .X(_04100_));
 sky130_fd_sc_hd__clkbuf_1 _08175_ (.A(_04100_),
    .X(_01512_));
 sky130_fd_sc_hd__buf_6 _08176_ (.A(net22),
    .X(_04101_));
 sky130_fd_sc_hd__buf_6 _08177_ (.A(_04101_),
    .X(_04102_));
 sky130_fd_sc_hd__mux2_1 _08178_ (.A0(net2081),
    .A1(_04102_),
    .S(_04078_),
    .X(_04103_));
 sky130_fd_sc_hd__clkbuf_1 _08179_ (.A(_04103_),
    .X(_01513_));
 sky130_fd_sc_hd__buf_8 _08180_ (.A(net23),
    .X(_04104_));
 sky130_fd_sc_hd__buf_6 _08181_ (.A(_04104_),
    .X(_04105_));
 sky130_fd_sc_hd__mux2_1 _08182_ (.A0(net2063),
    .A1(_04105_),
    .S(_04078_),
    .X(_04106_));
 sky130_fd_sc_hd__clkbuf_1 _08183_ (.A(_04106_),
    .X(_01514_));
 sky130_fd_sc_hd__buf_6 _08184_ (.A(net9),
    .X(_04107_));
 sky130_fd_sc_hd__buf_6 _08185_ (.A(_04107_),
    .X(_04108_));
 sky130_fd_sc_hd__mux2_1 _08186_ (.A0(net238),
    .A1(_04108_),
    .S(_04077_),
    .X(_04109_));
 sky130_fd_sc_hd__clkbuf_1 _08187_ (.A(_04109_),
    .X(_01515_));
 sky130_fd_sc_hd__buf_4 _08188_ (.A(net10),
    .X(_04110_));
 sky130_fd_sc_hd__buf_6 _08189_ (.A(_04110_),
    .X(_04111_));
 sky130_fd_sc_hd__mux2_1 _08190_ (.A0(net692),
    .A1(_04111_),
    .S(_04077_),
    .X(_04112_));
 sky130_fd_sc_hd__clkbuf_1 _08191_ (.A(_04112_),
    .X(_01516_));
 sky130_fd_sc_hd__buf_6 _08192_ (.A(net11),
    .X(_04113_));
 sky130_fd_sc_hd__buf_6 _08193_ (.A(_04113_),
    .X(_04114_));
 sky130_fd_sc_hd__mux2_1 _08194_ (.A0(net2054),
    .A1(_04114_),
    .S(_04077_),
    .X(_04115_));
 sky130_fd_sc_hd__clkbuf_1 _08195_ (.A(_04115_),
    .X(_01517_));
 sky130_fd_sc_hd__buf_6 _08196_ (.A(net12),
    .X(_04116_));
 sky130_fd_sc_hd__buf_6 _08197_ (.A(_04116_),
    .X(_04117_));
 sky130_fd_sc_hd__mux2_1 _08198_ (.A0(net2035),
    .A1(_04117_),
    .S(_04077_),
    .X(_04118_));
 sky130_fd_sc_hd__clkbuf_1 _08199_ (.A(_04118_),
    .X(_01518_));
 sky130_fd_sc_hd__buf_8 _08200_ (.A(net13),
    .X(_04119_));
 sky130_fd_sc_hd__buf_6 _08201_ (.A(_04119_),
    .X(_04120_));
 sky130_fd_sc_hd__mux2_1 _08202_ (.A0(net2060),
    .A1(_04120_),
    .S(_04077_),
    .X(_04121_));
 sky130_fd_sc_hd__clkbuf_1 _08203_ (.A(_04121_),
    .X(_01519_));
 sky130_fd_sc_hd__buf_8 _08204_ (.A(net14),
    .X(_04122_));
 sky130_fd_sc_hd__buf_6 _08205_ (.A(_04122_),
    .X(_04123_));
 sky130_fd_sc_hd__mux2_1 _08206_ (.A0(net1919),
    .A1(_04123_),
    .S(_04077_),
    .X(_04124_));
 sky130_fd_sc_hd__clkbuf_1 _08207_ (.A(_04124_),
    .X(_01520_));
 sky130_fd_sc_hd__buf_12 _08208_ (.A(_04069_),
    .X(_04125_));
 sky130_fd_sc_hd__or2_1 _08209_ (.A(_02505_),
    .B(_02404_),
    .X(_04126_));
 sky130_fd_sc_hd__buf_12 _08210_ (.A(_04126_),
    .X(_04127_));
 sky130_fd_sc_hd__nand2_1 _08211_ (.A(net7),
    .B(net24),
    .Y(_04128_));
 sky130_fd_sc_hd__or3_2 _08212_ (.A(_02357_),
    .B(net6),
    .C(_04128_),
    .X(_04129_));
 sky130_fd_sc_hd__or2_1 _08213_ (.A(_04127_),
    .B(_04129_),
    .X(_04130_));
 sky130_fd_sc_hd__clkbuf_4 _08214_ (.A(_04130_),
    .X(_04131_));
 sky130_fd_sc_hd__buf_4 _08215_ (.A(_04131_),
    .X(_04132_));
 sky130_fd_sc_hd__mux2_1 _08216_ (.A0(_04125_),
    .A1(net1196),
    .S(_04132_),
    .X(_04133_));
 sky130_fd_sc_hd__clkbuf_1 _08217_ (.A(_04133_),
    .X(_01521_));
 sky130_fd_sc_hd__buf_8 _08218_ (.A(_04080_),
    .X(_04134_));
 sky130_fd_sc_hd__mux2_1 _08219_ (.A0(_04134_),
    .A1(net1891),
    .S(_04132_),
    .X(_04135_));
 sky130_fd_sc_hd__clkbuf_1 _08220_ (.A(_04135_),
    .X(_01522_));
 sky130_fd_sc_hd__buf_12 _08221_ (.A(_04083_),
    .X(_04136_));
 sky130_fd_sc_hd__mux2_1 _08222_ (.A0(_04136_),
    .A1(net1797),
    .S(_04132_),
    .X(_04137_));
 sky130_fd_sc_hd__clkbuf_1 _08223_ (.A(_04137_),
    .X(_01523_));
 sky130_fd_sc_hd__buf_12 _08224_ (.A(_04086_),
    .X(_04138_));
 sky130_fd_sc_hd__mux2_1 _08225_ (.A0(_04138_),
    .A1(net1822),
    .S(_04132_),
    .X(_04139_));
 sky130_fd_sc_hd__clkbuf_1 _08226_ (.A(_04139_),
    .X(_01524_));
 sky130_fd_sc_hd__buf_12 _08227_ (.A(_04089_),
    .X(_04140_));
 sky130_fd_sc_hd__mux2_1 _08228_ (.A0(_04140_),
    .A1(net1548),
    .S(_04132_),
    .X(_04141_));
 sky130_fd_sc_hd__clkbuf_1 _08229_ (.A(_04141_),
    .X(_01525_));
 sky130_fd_sc_hd__clkbuf_16 _08230_ (.A(_04092_),
    .X(_04142_));
 sky130_fd_sc_hd__mux2_1 _08231_ (.A0(_04142_),
    .A1(net1791),
    .S(_04132_),
    .X(_04143_));
 sky130_fd_sc_hd__clkbuf_1 _08232_ (.A(_04143_),
    .X(_01526_));
 sky130_fd_sc_hd__buf_12 _08233_ (.A(_04095_),
    .X(_04144_));
 sky130_fd_sc_hd__mux2_1 _08234_ (.A0(_04144_),
    .A1(net1750),
    .S(_04132_),
    .X(_04145_));
 sky130_fd_sc_hd__clkbuf_1 _08235_ (.A(_04145_),
    .X(_01527_));
 sky130_fd_sc_hd__buf_12 _08236_ (.A(_04098_),
    .X(_04146_));
 sky130_fd_sc_hd__mux2_1 _08237_ (.A0(_04146_),
    .A1(net910),
    .S(_04132_),
    .X(_04147_));
 sky130_fd_sc_hd__clkbuf_1 _08238_ (.A(_04147_),
    .X(_01528_));
 sky130_fd_sc_hd__buf_12 _08239_ (.A(_04101_),
    .X(_04148_));
 sky130_fd_sc_hd__mux2_1 _08240_ (.A0(_04148_),
    .A1(net1469),
    .S(_04132_),
    .X(_04149_));
 sky130_fd_sc_hd__clkbuf_1 _08241_ (.A(_04149_),
    .X(_01529_));
 sky130_fd_sc_hd__buf_12 _08242_ (.A(_04104_),
    .X(_04150_));
 sky130_fd_sc_hd__mux2_1 _08243_ (.A0(_04150_),
    .A1(net1543),
    .S(_04132_),
    .X(_04151_));
 sky130_fd_sc_hd__clkbuf_1 _08244_ (.A(_04151_),
    .X(_01530_));
 sky130_fd_sc_hd__buf_12 _08245_ (.A(_04107_),
    .X(_04152_));
 sky130_fd_sc_hd__mux2_1 _08246_ (.A0(_04152_),
    .A1(net1161),
    .S(_04131_),
    .X(_04153_));
 sky130_fd_sc_hd__clkbuf_1 _08247_ (.A(_04153_),
    .X(_01531_));
 sky130_fd_sc_hd__buf_12 _08248_ (.A(_04110_),
    .X(_04154_));
 sky130_fd_sc_hd__mux2_1 _08249_ (.A0(_04154_),
    .A1(net1488),
    .S(_04131_),
    .X(_04155_));
 sky130_fd_sc_hd__clkbuf_1 _08250_ (.A(_04155_),
    .X(_01532_));
 sky130_fd_sc_hd__buf_12 _08251_ (.A(_04113_),
    .X(_04156_));
 sky130_fd_sc_hd__mux2_1 _08252_ (.A0(_04156_),
    .A1(net1495),
    .S(_04131_),
    .X(_04157_));
 sky130_fd_sc_hd__clkbuf_1 _08253_ (.A(_04157_),
    .X(_01533_));
 sky130_fd_sc_hd__clkbuf_16 _08254_ (.A(_04116_),
    .X(_04158_));
 sky130_fd_sc_hd__mux2_1 _08255_ (.A0(_04158_),
    .A1(net975),
    .S(_04131_),
    .X(_04159_));
 sky130_fd_sc_hd__clkbuf_1 _08256_ (.A(_04159_),
    .X(_01534_));
 sky130_fd_sc_hd__buf_12 _08257_ (.A(_04119_),
    .X(_04160_));
 sky130_fd_sc_hd__mux2_1 _08258_ (.A0(_04160_),
    .A1(net1824),
    .S(_04131_),
    .X(_04161_));
 sky130_fd_sc_hd__clkbuf_1 _08259_ (.A(_04161_),
    .X(_01535_));
 sky130_fd_sc_hd__buf_12 _08260_ (.A(_04122_),
    .X(_04162_));
 sky130_fd_sc_hd__mux2_1 _08261_ (.A0(_04162_),
    .A1(net1749),
    .S(_04131_),
    .X(_04163_));
 sky130_fd_sc_hd__clkbuf_1 _08262_ (.A(_04163_),
    .X(_01536_));
 sky130_fd_sc_hd__or3_1 _08263_ (.A(_02707_),
    .B(_03092_),
    .C(_04075_),
    .X(_04164_));
 sky130_fd_sc_hd__clkbuf_4 _08264_ (.A(_04164_),
    .X(_04165_));
 sky130_fd_sc_hd__buf_4 _08265_ (.A(_04165_),
    .X(_04166_));
 sky130_fd_sc_hd__mux2_1 _08266_ (.A0(_04125_),
    .A1(net1062),
    .S(_04166_),
    .X(_04167_));
 sky130_fd_sc_hd__clkbuf_1 _08267_ (.A(_04167_),
    .X(_01537_));
 sky130_fd_sc_hd__mux2_1 _08268_ (.A0(_04134_),
    .A1(net979),
    .S(_04166_),
    .X(_04168_));
 sky130_fd_sc_hd__clkbuf_1 _08269_ (.A(_04168_),
    .X(_01538_));
 sky130_fd_sc_hd__mux2_1 _08270_ (.A0(_04136_),
    .A1(net1671),
    .S(_04166_),
    .X(_04169_));
 sky130_fd_sc_hd__clkbuf_1 _08271_ (.A(_04169_),
    .X(_01539_));
 sky130_fd_sc_hd__mux2_1 _08272_ (.A0(_04138_),
    .A1(net1189),
    .S(_04166_),
    .X(_04170_));
 sky130_fd_sc_hd__clkbuf_1 _08273_ (.A(_04170_),
    .X(_01540_));
 sky130_fd_sc_hd__mux2_1 _08274_ (.A0(_04140_),
    .A1(net1102),
    .S(_04166_),
    .X(_04171_));
 sky130_fd_sc_hd__clkbuf_1 _08275_ (.A(_04171_),
    .X(_01541_));
 sky130_fd_sc_hd__mux2_1 _08276_ (.A0(_04142_),
    .A1(net1371),
    .S(_04166_),
    .X(_04172_));
 sky130_fd_sc_hd__clkbuf_1 _08277_ (.A(_04172_),
    .X(_01542_));
 sky130_fd_sc_hd__mux2_1 _08278_ (.A0(_04144_),
    .A1(net518),
    .S(_04166_),
    .X(_04173_));
 sky130_fd_sc_hd__clkbuf_1 _08279_ (.A(_04173_),
    .X(_01543_));
 sky130_fd_sc_hd__mux2_1 _08280_ (.A0(_04146_),
    .A1(net1706),
    .S(_04166_),
    .X(_04174_));
 sky130_fd_sc_hd__clkbuf_1 _08281_ (.A(_04174_),
    .X(_01544_));
 sky130_fd_sc_hd__mux2_1 _08282_ (.A0(_04148_),
    .A1(net1391),
    .S(_04166_),
    .X(_04175_));
 sky130_fd_sc_hd__clkbuf_1 _08283_ (.A(_04175_),
    .X(_01545_));
 sky130_fd_sc_hd__mux2_1 _08284_ (.A0(_04150_),
    .A1(net885),
    .S(_04166_),
    .X(_04176_));
 sky130_fd_sc_hd__clkbuf_1 _08285_ (.A(_04176_),
    .X(_01546_));
 sky130_fd_sc_hd__mux2_1 _08286_ (.A0(_04152_),
    .A1(net1687),
    .S(_04165_),
    .X(_04177_));
 sky130_fd_sc_hd__clkbuf_1 _08287_ (.A(_04177_),
    .X(_01547_));
 sky130_fd_sc_hd__mux2_1 _08288_ (.A0(_04154_),
    .A1(net1082),
    .S(_04165_),
    .X(_04178_));
 sky130_fd_sc_hd__clkbuf_1 _08289_ (.A(_04178_),
    .X(_01548_));
 sky130_fd_sc_hd__mux2_1 _08290_ (.A0(_04156_),
    .A1(net508),
    .S(_04165_),
    .X(_04179_));
 sky130_fd_sc_hd__clkbuf_1 _08291_ (.A(_04179_),
    .X(_01549_));
 sky130_fd_sc_hd__mux2_1 _08292_ (.A0(_04158_),
    .A1(net1319),
    .S(_04165_),
    .X(_04180_));
 sky130_fd_sc_hd__clkbuf_1 _08293_ (.A(_04180_),
    .X(_01550_));
 sky130_fd_sc_hd__mux2_1 _08294_ (.A0(_04160_),
    .A1(net1424),
    .S(_04165_),
    .X(_04181_));
 sky130_fd_sc_hd__clkbuf_1 _08295_ (.A(_04181_),
    .X(_01551_));
 sky130_fd_sc_hd__mux2_1 _08296_ (.A0(_04162_),
    .A1(net1227),
    .S(_04165_),
    .X(_04182_));
 sky130_fd_sc_hd__clkbuf_1 _08297_ (.A(_04182_),
    .X(_01552_));
 sky130_fd_sc_hd__or2_1 _08298_ (.A(_02497_),
    .B(_02404_),
    .X(_04183_));
 sky130_fd_sc_hd__buf_12 _08299_ (.A(_04183_),
    .X(_04184_));
 sky130_fd_sc_hd__or3_4 _08300_ (.A(_02420_),
    .B(net6),
    .C(_04128_),
    .X(_04185_));
 sky130_fd_sc_hd__buf_8 _08301_ (.A(_04185_),
    .X(_04186_));
 sky130_fd_sc_hd__nor2_4 _08302_ (.A(_04184_),
    .B(_04186_),
    .Y(_04187_));
 sky130_fd_sc_hd__buf_4 _08303_ (.A(_04187_),
    .X(_04188_));
 sky130_fd_sc_hd__mux2_1 _08304_ (.A0(net1998),
    .A1(_04070_),
    .S(_04188_),
    .X(_04189_));
 sky130_fd_sc_hd__clkbuf_1 _08305_ (.A(_04189_),
    .X(_01553_));
 sky130_fd_sc_hd__mux2_1 _08306_ (.A0(net2072),
    .A1(_04081_),
    .S(_04188_),
    .X(_04190_));
 sky130_fd_sc_hd__clkbuf_1 _08307_ (.A(_04190_),
    .X(_01554_));
 sky130_fd_sc_hd__mux2_1 _08308_ (.A0(net1553),
    .A1(_04084_),
    .S(_04188_),
    .X(_04191_));
 sky130_fd_sc_hd__clkbuf_1 _08309_ (.A(_04191_),
    .X(_01555_));
 sky130_fd_sc_hd__mux2_1 _08310_ (.A0(net2040),
    .A1(_04087_),
    .S(_04188_),
    .X(_04192_));
 sky130_fd_sc_hd__clkbuf_1 _08311_ (.A(_04192_),
    .X(_01556_));
 sky130_fd_sc_hd__mux2_1 _08312_ (.A0(net1678),
    .A1(_04090_),
    .S(_04188_),
    .X(_04193_));
 sky130_fd_sc_hd__clkbuf_1 _08313_ (.A(_04193_),
    .X(_01557_));
 sky130_fd_sc_hd__mux2_1 _08314_ (.A0(net532),
    .A1(_04093_),
    .S(_04188_),
    .X(_04194_));
 sky130_fd_sc_hd__clkbuf_1 _08315_ (.A(_04194_),
    .X(_01558_));
 sky130_fd_sc_hd__mux2_1 _08316_ (.A0(net1047),
    .A1(_04096_),
    .S(_04188_),
    .X(_04195_));
 sky130_fd_sc_hd__clkbuf_1 _08317_ (.A(_04195_),
    .X(_01559_));
 sky130_fd_sc_hd__mux2_1 _08318_ (.A0(net1937),
    .A1(_04099_),
    .S(_04188_),
    .X(_04196_));
 sky130_fd_sc_hd__clkbuf_1 _08319_ (.A(_04196_),
    .X(_01560_));
 sky130_fd_sc_hd__mux2_1 _08320_ (.A0(net1874),
    .A1(_04102_),
    .S(_04188_),
    .X(_04197_));
 sky130_fd_sc_hd__clkbuf_1 _08321_ (.A(_04197_),
    .X(_01561_));
 sky130_fd_sc_hd__mux2_1 _08322_ (.A0(net1944),
    .A1(_04105_),
    .S(_04188_),
    .X(_04198_));
 sky130_fd_sc_hd__clkbuf_1 _08323_ (.A(_04198_),
    .X(_01562_));
 sky130_fd_sc_hd__mux2_1 _08324_ (.A0(net1662),
    .A1(_04108_),
    .S(_04187_),
    .X(_04199_));
 sky130_fd_sc_hd__clkbuf_1 _08325_ (.A(_04199_),
    .X(_01563_));
 sky130_fd_sc_hd__mux2_1 _08326_ (.A0(net1207),
    .A1(_04111_),
    .S(_04187_),
    .X(_04200_));
 sky130_fd_sc_hd__clkbuf_1 _08327_ (.A(_04200_),
    .X(_01564_));
 sky130_fd_sc_hd__mux2_1 _08328_ (.A0(net630),
    .A1(_04114_),
    .S(_04187_),
    .X(_04201_));
 sky130_fd_sc_hd__clkbuf_1 _08329_ (.A(_04201_),
    .X(_01565_));
 sky130_fd_sc_hd__mux2_1 _08330_ (.A0(net1435),
    .A1(_04117_),
    .S(_04187_),
    .X(_04202_));
 sky130_fd_sc_hd__clkbuf_1 _08331_ (.A(_04202_),
    .X(_01566_));
 sky130_fd_sc_hd__mux2_1 _08332_ (.A0(net1003),
    .A1(_04120_),
    .S(_04187_),
    .X(_04203_));
 sky130_fd_sc_hd__clkbuf_1 _08333_ (.A(_04203_),
    .X(_01567_));
 sky130_fd_sc_hd__mux2_1 _08334_ (.A0(net466),
    .A1(_04123_),
    .S(_04187_),
    .X(_04204_));
 sky130_fd_sc_hd__clkbuf_1 _08335_ (.A(_04204_),
    .X(_01568_));
 sky130_fd_sc_hd__or3_1 _08336_ (.A(_04059_),
    .B(_03092_),
    .C(_04185_),
    .X(_04205_));
 sky130_fd_sc_hd__buf_2 _08337_ (.A(_04205_),
    .X(_04206_));
 sky130_fd_sc_hd__buf_4 _08338_ (.A(_04206_),
    .X(_04207_));
 sky130_fd_sc_hd__mux2_1 _08339_ (.A0(_04125_),
    .A1(net1779),
    .S(_04207_),
    .X(_04208_));
 sky130_fd_sc_hd__clkbuf_1 _08340_ (.A(_04208_),
    .X(_01569_));
 sky130_fd_sc_hd__mux2_1 _08341_ (.A0(_04134_),
    .A1(net1607),
    .S(_04207_),
    .X(_04209_));
 sky130_fd_sc_hd__clkbuf_1 _08342_ (.A(_04209_),
    .X(_01570_));
 sky130_fd_sc_hd__mux2_1 _08343_ (.A0(_04136_),
    .A1(net1537),
    .S(_04207_),
    .X(_04210_));
 sky130_fd_sc_hd__clkbuf_1 _08344_ (.A(_04210_),
    .X(_01571_));
 sky130_fd_sc_hd__mux2_1 _08345_ (.A0(_04138_),
    .A1(net1914),
    .S(_04207_),
    .X(_04211_));
 sky130_fd_sc_hd__clkbuf_1 _08346_ (.A(_04211_),
    .X(_01572_));
 sky130_fd_sc_hd__mux2_1 _08347_ (.A0(_04140_),
    .A1(net1188),
    .S(_04207_),
    .X(_04212_));
 sky130_fd_sc_hd__clkbuf_1 _08348_ (.A(_04212_),
    .X(_01573_));
 sky130_fd_sc_hd__mux2_1 _08349_ (.A0(_04142_),
    .A1(net1213),
    .S(_04207_),
    .X(_04213_));
 sky130_fd_sc_hd__clkbuf_1 _08350_ (.A(_04213_),
    .X(_01574_));
 sky130_fd_sc_hd__mux2_1 _08351_ (.A0(_04144_),
    .A1(net1317),
    .S(_04207_),
    .X(_04214_));
 sky130_fd_sc_hd__clkbuf_1 _08352_ (.A(_04214_),
    .X(_01575_));
 sky130_fd_sc_hd__mux2_1 _08353_ (.A0(_04146_),
    .A1(net1335),
    .S(_04207_),
    .X(_04215_));
 sky130_fd_sc_hd__clkbuf_1 _08354_ (.A(_04215_),
    .X(_01576_));
 sky130_fd_sc_hd__mux2_1 _08355_ (.A0(_04148_),
    .A1(net1855),
    .S(_04207_),
    .X(_04216_));
 sky130_fd_sc_hd__clkbuf_1 _08356_ (.A(_04216_),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_1 _08357_ (.A0(_04150_),
    .A1(net1612),
    .S(_04207_),
    .X(_04217_));
 sky130_fd_sc_hd__clkbuf_1 _08358_ (.A(_04217_),
    .X(_01578_));
 sky130_fd_sc_hd__mux2_1 _08359_ (.A0(_04152_),
    .A1(net1534),
    .S(_04206_),
    .X(_04218_));
 sky130_fd_sc_hd__clkbuf_1 _08360_ (.A(_04218_),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_1 _08361_ (.A0(_04154_),
    .A1(net1975),
    .S(_04206_),
    .X(_04219_));
 sky130_fd_sc_hd__clkbuf_1 _08362_ (.A(_04219_),
    .X(_01580_));
 sky130_fd_sc_hd__mux2_1 _08363_ (.A0(_04156_),
    .A1(net1995),
    .S(_04206_),
    .X(_04220_));
 sky130_fd_sc_hd__clkbuf_1 _08364_ (.A(_04220_),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _08365_ (.A0(_04158_),
    .A1(net1759),
    .S(_04206_),
    .X(_04221_));
 sky130_fd_sc_hd__clkbuf_1 _08366_ (.A(_04221_),
    .X(_01582_));
 sky130_fd_sc_hd__mux2_1 _08367_ (.A0(_04160_),
    .A1(net1783),
    .S(_04206_),
    .X(_04222_));
 sky130_fd_sc_hd__clkbuf_1 _08368_ (.A(_04222_),
    .X(_01583_));
 sky130_fd_sc_hd__mux2_1 _08369_ (.A0(_04162_),
    .A1(net1531),
    .S(_04206_),
    .X(_04223_));
 sky130_fd_sc_hd__clkbuf_1 _08370_ (.A(_04223_),
    .X(_01584_));
 sky130_fd_sc_hd__or2_1 _08371_ (.A(_02495_),
    .B(_02400_),
    .X(_04224_));
 sky130_fd_sc_hd__buf_12 _08372_ (.A(_04224_),
    .X(_04225_));
 sky130_fd_sc_hd__or3_4 _08373_ (.A(_02357_),
    .B(net6),
    .C(_04074_),
    .X(_04226_));
 sky130_fd_sc_hd__buf_12 _08374_ (.A(_04226_),
    .X(_04227_));
 sky130_fd_sc_hd__nor2_4 _08375_ (.A(_04225_),
    .B(_04227_),
    .Y(_04228_));
 sky130_fd_sc_hd__buf_4 _08376_ (.A(_04228_),
    .X(_04229_));
 sky130_fd_sc_hd__mux2_1 _08377_ (.A0(net1653),
    .A1(_04070_),
    .S(_04229_),
    .X(_04230_));
 sky130_fd_sc_hd__clkbuf_1 _08378_ (.A(_04230_),
    .X(_01585_));
 sky130_fd_sc_hd__mux2_1 _08379_ (.A0(net779),
    .A1(_04081_),
    .S(_04229_),
    .X(_04231_));
 sky130_fd_sc_hd__clkbuf_1 _08380_ (.A(_04231_),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _08381_ (.A0(net1940),
    .A1(_04084_),
    .S(_04229_),
    .X(_04232_));
 sky130_fd_sc_hd__clkbuf_1 _08382_ (.A(_04232_),
    .X(_01587_));
 sky130_fd_sc_hd__mux2_1 _08383_ (.A0(net1628),
    .A1(_04087_),
    .S(_04229_),
    .X(_04233_));
 sky130_fd_sc_hd__clkbuf_1 _08384_ (.A(_04233_),
    .X(_01588_));
 sky130_fd_sc_hd__mux2_1 _08385_ (.A0(net1826),
    .A1(_04090_),
    .S(_04229_),
    .X(_04234_));
 sky130_fd_sc_hd__clkbuf_1 _08386_ (.A(_04234_),
    .X(_01589_));
 sky130_fd_sc_hd__mux2_1 _08387_ (.A0(net316),
    .A1(_04093_),
    .S(_04229_),
    .X(_04235_));
 sky130_fd_sc_hd__clkbuf_1 _08388_ (.A(_04235_),
    .X(_01590_));
 sky130_fd_sc_hd__mux2_1 _08389_ (.A0(net1305),
    .A1(_04096_),
    .S(_04229_),
    .X(_04236_));
 sky130_fd_sc_hd__clkbuf_1 _08390_ (.A(_04236_),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_1 _08391_ (.A0(net587),
    .A1(_04099_),
    .S(_04229_),
    .X(_04237_));
 sky130_fd_sc_hd__clkbuf_1 _08392_ (.A(_04237_),
    .X(_01592_));
 sky130_fd_sc_hd__mux2_1 _08393_ (.A0(net1856),
    .A1(_04102_),
    .S(_04229_),
    .X(_04238_));
 sky130_fd_sc_hd__clkbuf_1 _08394_ (.A(_04238_),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _08395_ (.A0(net871),
    .A1(_04105_),
    .S(_04229_),
    .X(_04239_));
 sky130_fd_sc_hd__clkbuf_1 _08396_ (.A(_04239_),
    .X(_01594_));
 sky130_fd_sc_hd__mux2_1 _08397_ (.A0(net832),
    .A1(_04108_),
    .S(_04228_),
    .X(_04240_));
 sky130_fd_sc_hd__clkbuf_1 _08398_ (.A(_04240_),
    .X(_01595_));
 sky130_fd_sc_hd__mux2_1 _08399_ (.A0(net1452),
    .A1(_04111_),
    .S(_04228_),
    .X(_04241_));
 sky130_fd_sc_hd__clkbuf_1 _08400_ (.A(_04241_),
    .X(_01596_));
 sky130_fd_sc_hd__mux2_1 _08401_ (.A0(net1836),
    .A1(_04114_),
    .S(_04228_),
    .X(_04242_));
 sky130_fd_sc_hd__clkbuf_1 _08402_ (.A(_04242_),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _08403_ (.A0(net279),
    .A1(_04117_),
    .S(_04228_),
    .X(_04243_));
 sky130_fd_sc_hd__clkbuf_1 _08404_ (.A(_04243_),
    .X(_01598_));
 sky130_fd_sc_hd__mux2_1 _08405_ (.A0(net909),
    .A1(_04120_),
    .S(_04228_),
    .X(_04244_));
 sky130_fd_sc_hd__clkbuf_1 _08406_ (.A(_04244_),
    .X(_01599_));
 sky130_fd_sc_hd__mux2_1 _08407_ (.A0(net1318),
    .A1(_04123_),
    .S(_04228_),
    .X(_04245_));
 sky130_fd_sc_hd__clkbuf_1 _08408_ (.A(_04245_),
    .X(_01600_));
 sky130_fd_sc_hd__or3_4 _08409_ (.A(_02420_),
    .B(_02355_),
    .C(_04074_),
    .X(_04246_));
 sky130_fd_sc_hd__or3_1 _08410_ (.A(_02702_),
    .B(_03092_),
    .C(_04246_),
    .X(_04247_));
 sky130_fd_sc_hd__clkbuf_4 _08411_ (.A(_04247_),
    .X(_04248_));
 sky130_fd_sc_hd__clkbuf_8 _08412_ (.A(_04248_),
    .X(_04249_));
 sky130_fd_sc_hd__mux2_1 _08413_ (.A0(_04125_),
    .A1(net1511),
    .S(_04249_),
    .X(_04250_));
 sky130_fd_sc_hd__clkbuf_1 _08414_ (.A(_04250_),
    .X(_01601_));
 sky130_fd_sc_hd__mux2_1 _08415_ (.A0(_04134_),
    .A1(net1234),
    .S(_04249_),
    .X(_04251_));
 sky130_fd_sc_hd__clkbuf_1 _08416_ (.A(_04251_),
    .X(_01602_));
 sky130_fd_sc_hd__mux2_1 _08417_ (.A0(_04136_),
    .A1(net2048),
    .S(_04249_),
    .X(_04252_));
 sky130_fd_sc_hd__clkbuf_1 _08418_ (.A(_04252_),
    .X(_01603_));
 sky130_fd_sc_hd__mux2_1 _08419_ (.A0(_04138_),
    .A1(net1184),
    .S(_04249_),
    .X(_04253_));
 sky130_fd_sc_hd__clkbuf_1 _08420_ (.A(_04253_),
    .X(_01604_));
 sky130_fd_sc_hd__mux2_1 _08421_ (.A0(_04140_),
    .A1(net666),
    .S(_04249_),
    .X(_04254_));
 sky130_fd_sc_hd__clkbuf_1 _08422_ (.A(_04254_),
    .X(_01605_));
 sky130_fd_sc_hd__mux2_1 _08423_ (.A0(_04142_),
    .A1(net977),
    .S(_04249_),
    .X(_04255_));
 sky130_fd_sc_hd__clkbuf_1 _08424_ (.A(_04255_),
    .X(_01606_));
 sky130_fd_sc_hd__mux2_1 _08425_ (.A0(_04144_),
    .A1(net275),
    .S(_04249_),
    .X(_04256_));
 sky130_fd_sc_hd__clkbuf_1 _08426_ (.A(_04256_),
    .X(_01607_));
 sky130_fd_sc_hd__mux2_1 _08427_ (.A0(_04146_),
    .A1(net1898),
    .S(_04249_),
    .X(_04257_));
 sky130_fd_sc_hd__clkbuf_1 _08428_ (.A(_04257_),
    .X(_01608_));
 sky130_fd_sc_hd__mux2_1 _08429_ (.A0(_04148_),
    .A1(net1902),
    .S(_04249_),
    .X(_04258_));
 sky130_fd_sc_hd__clkbuf_1 _08430_ (.A(_04258_),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _08431_ (.A0(_04150_),
    .A1(net817),
    .S(_04249_),
    .X(_04259_));
 sky130_fd_sc_hd__clkbuf_1 _08432_ (.A(_04259_),
    .X(_01610_));
 sky130_fd_sc_hd__mux2_1 _08433_ (.A0(_04152_),
    .A1(net2000),
    .S(_04248_),
    .X(_04260_));
 sky130_fd_sc_hd__clkbuf_1 _08434_ (.A(_04260_),
    .X(_01611_));
 sky130_fd_sc_hd__mux2_1 _08435_ (.A0(_04154_),
    .A1(net1403),
    .S(_04248_),
    .X(_04261_));
 sky130_fd_sc_hd__clkbuf_1 _08436_ (.A(_04261_),
    .X(_01612_));
 sky130_fd_sc_hd__mux2_1 _08437_ (.A0(_04156_),
    .A1(net1512),
    .S(_04248_),
    .X(_04262_));
 sky130_fd_sc_hd__clkbuf_1 _08438_ (.A(_04262_),
    .X(_01613_));
 sky130_fd_sc_hd__mux2_1 _08439_ (.A0(_04158_),
    .A1(net1221),
    .S(_04248_),
    .X(_04263_));
 sky130_fd_sc_hd__clkbuf_1 _08440_ (.A(_04263_),
    .X(_01614_));
 sky130_fd_sc_hd__mux2_1 _08441_ (.A0(_04160_),
    .A1(net1587),
    .S(_04248_),
    .X(_04264_));
 sky130_fd_sc_hd__clkbuf_1 _08442_ (.A(_04264_),
    .X(_01615_));
 sky130_fd_sc_hd__mux2_1 _08443_ (.A0(_04162_),
    .A1(net739),
    .S(_04248_),
    .X(_04265_));
 sky130_fd_sc_hd__clkbuf_1 _08444_ (.A(_04265_),
    .X(_01616_));
 sky130_fd_sc_hd__or3_1 _08445_ (.A(_04059_),
    .B(_02654_),
    .C(_04226_),
    .X(_04266_));
 sky130_fd_sc_hd__clkbuf_4 _08446_ (.A(_04266_),
    .X(_04267_));
 sky130_fd_sc_hd__buf_4 _08447_ (.A(_04267_),
    .X(_04268_));
 sky130_fd_sc_hd__mux2_1 _08448_ (.A0(_04125_),
    .A1(net1611),
    .S(_04268_),
    .X(_04269_));
 sky130_fd_sc_hd__clkbuf_1 _08449_ (.A(_04269_),
    .X(_01617_));
 sky130_fd_sc_hd__mux2_1 _08450_ (.A0(_04134_),
    .A1(net1400),
    .S(_04268_),
    .X(_04270_));
 sky130_fd_sc_hd__clkbuf_1 _08451_ (.A(_04270_),
    .X(_01618_));
 sky130_fd_sc_hd__mux2_1 _08452_ (.A0(_04136_),
    .A1(net1732),
    .S(_04268_),
    .X(_04271_));
 sky130_fd_sc_hd__clkbuf_1 _08453_ (.A(_04271_),
    .X(_01619_));
 sky130_fd_sc_hd__mux2_1 _08454_ (.A0(_04138_),
    .A1(net1434),
    .S(_04268_),
    .X(_04272_));
 sky130_fd_sc_hd__clkbuf_1 _08455_ (.A(_04272_),
    .X(_01620_));
 sky130_fd_sc_hd__mux2_1 _08456_ (.A0(_04140_),
    .A1(net1510),
    .S(_04268_),
    .X(_04273_));
 sky130_fd_sc_hd__clkbuf_1 _08457_ (.A(_04273_),
    .X(_01621_));
 sky130_fd_sc_hd__mux2_1 _08458_ (.A0(_04142_),
    .A1(net1163),
    .S(_04268_),
    .X(_04274_));
 sky130_fd_sc_hd__clkbuf_1 _08459_ (.A(_04274_),
    .X(_01622_));
 sky130_fd_sc_hd__mux2_1 _08460_ (.A0(_04144_),
    .A1(net824),
    .S(_04268_),
    .X(_04275_));
 sky130_fd_sc_hd__clkbuf_1 _08461_ (.A(_04275_),
    .X(_01623_));
 sky130_fd_sc_hd__mux2_1 _08462_ (.A0(_04146_),
    .A1(net2002),
    .S(_04268_),
    .X(_04276_));
 sky130_fd_sc_hd__clkbuf_1 _08463_ (.A(_04276_),
    .X(_01624_));
 sky130_fd_sc_hd__mux2_1 _08464_ (.A0(_04148_),
    .A1(net1571),
    .S(_04268_),
    .X(_04277_));
 sky130_fd_sc_hd__clkbuf_1 _08465_ (.A(_04277_),
    .X(_01625_));
 sky130_fd_sc_hd__mux2_1 _08466_ (.A0(_04150_),
    .A1(net1380),
    .S(_04268_),
    .X(_04278_));
 sky130_fd_sc_hd__clkbuf_1 _08467_ (.A(_04278_),
    .X(_01626_));
 sky130_fd_sc_hd__mux2_1 _08468_ (.A0(_04152_),
    .A1(net1843),
    .S(_04267_),
    .X(_04279_));
 sky130_fd_sc_hd__clkbuf_1 _08469_ (.A(_04279_),
    .X(_01627_));
 sky130_fd_sc_hd__mux2_1 _08470_ (.A0(_04154_),
    .A1(net2030),
    .S(_04267_),
    .X(_04280_));
 sky130_fd_sc_hd__clkbuf_1 _08471_ (.A(_04280_),
    .X(_01628_));
 sky130_fd_sc_hd__mux2_1 _08472_ (.A0(_04156_),
    .A1(net2059),
    .S(_04267_),
    .X(_04281_));
 sky130_fd_sc_hd__clkbuf_1 _08473_ (.A(_04281_),
    .X(_01629_));
 sky130_fd_sc_hd__mux2_1 _08474_ (.A0(_04158_),
    .A1(net1621),
    .S(_04267_),
    .X(_04282_));
 sky130_fd_sc_hd__clkbuf_1 _08475_ (.A(_04282_),
    .X(_01630_));
 sky130_fd_sc_hd__mux2_1 _08476_ (.A0(_04160_),
    .A1(net1990),
    .S(_04267_),
    .X(_04283_));
 sky130_fd_sc_hd__clkbuf_1 _08477_ (.A(_04283_),
    .X(_01631_));
 sky130_fd_sc_hd__mux2_1 _08478_ (.A0(_04162_),
    .A1(net2043),
    .S(_04267_),
    .X(_04284_));
 sky130_fd_sc_hd__clkbuf_1 _08479_ (.A(_04284_),
    .X(_01632_));
 sky130_fd_sc_hd__or3_4 _08480_ (.A(net5),
    .B(_02355_),
    .C(_04128_),
    .X(_04285_));
 sky130_fd_sc_hd__buf_6 _08481_ (.A(_04285_),
    .X(_04286_));
 sky130_fd_sc_hd__or2_1 _08482_ (.A(_04225_),
    .B(_04286_),
    .X(_04287_));
 sky130_fd_sc_hd__clkbuf_4 _08483_ (.A(_04287_),
    .X(_04288_));
 sky130_fd_sc_hd__clkbuf_8 _08484_ (.A(_04288_),
    .X(_04289_));
 sky130_fd_sc_hd__mux2_1 _08485_ (.A0(_04125_),
    .A1(net1423),
    .S(_04289_),
    .X(_04290_));
 sky130_fd_sc_hd__clkbuf_1 _08486_ (.A(_04290_),
    .X(_01633_));
 sky130_fd_sc_hd__mux2_1 _08487_ (.A0(_04134_),
    .A1(net940),
    .S(_04289_),
    .X(_04291_));
 sky130_fd_sc_hd__clkbuf_1 _08488_ (.A(_04291_),
    .X(_01634_));
 sky130_fd_sc_hd__mux2_1 _08489_ (.A0(_04136_),
    .A1(net1059),
    .S(_04289_),
    .X(_04292_));
 sky130_fd_sc_hd__clkbuf_1 _08490_ (.A(_04292_),
    .X(_01635_));
 sky130_fd_sc_hd__mux2_1 _08491_ (.A0(_04138_),
    .A1(net1090),
    .S(_04289_),
    .X(_04293_));
 sky130_fd_sc_hd__clkbuf_1 _08492_ (.A(_04293_),
    .X(_01636_));
 sky130_fd_sc_hd__mux2_1 _08493_ (.A0(_04140_),
    .A1(net715),
    .S(_04289_),
    .X(_04294_));
 sky130_fd_sc_hd__clkbuf_1 _08494_ (.A(_04294_),
    .X(_01637_));
 sky130_fd_sc_hd__mux2_1 _08495_ (.A0(_04142_),
    .A1(net1383),
    .S(_04289_),
    .X(_04295_));
 sky130_fd_sc_hd__clkbuf_1 _08496_ (.A(_04295_),
    .X(_01638_));
 sky130_fd_sc_hd__mux2_1 _08497_ (.A0(_04144_),
    .A1(net551),
    .S(_04289_),
    .X(_04296_));
 sky130_fd_sc_hd__clkbuf_1 _08498_ (.A(_04296_),
    .X(_01639_));
 sky130_fd_sc_hd__mux2_1 _08499_ (.A0(_04146_),
    .A1(net1541),
    .S(_04289_),
    .X(_04297_));
 sky130_fd_sc_hd__clkbuf_1 _08500_ (.A(_04297_),
    .X(_01640_));
 sky130_fd_sc_hd__mux2_1 _08501_ (.A0(_04148_),
    .A1(net517),
    .S(_04289_),
    .X(_04298_));
 sky130_fd_sc_hd__clkbuf_1 _08502_ (.A(_04298_),
    .X(_01641_));
 sky130_fd_sc_hd__mux2_1 _08503_ (.A0(_04150_),
    .A1(net913),
    .S(_04289_),
    .X(_04299_));
 sky130_fd_sc_hd__clkbuf_1 _08504_ (.A(_04299_),
    .X(_01642_));
 sky130_fd_sc_hd__mux2_1 _08505_ (.A0(_04152_),
    .A1(net917),
    .S(_04288_),
    .X(_04300_));
 sky130_fd_sc_hd__clkbuf_1 _08506_ (.A(_04300_),
    .X(_01643_));
 sky130_fd_sc_hd__mux2_1 _08507_ (.A0(_04154_),
    .A1(net1589),
    .S(_04288_),
    .X(_04301_));
 sky130_fd_sc_hd__clkbuf_1 _08508_ (.A(_04301_),
    .X(_01644_));
 sky130_fd_sc_hd__mux2_1 _08509_ (.A0(_04156_),
    .A1(net1513),
    .S(_04288_),
    .X(_04302_));
 sky130_fd_sc_hd__clkbuf_1 _08510_ (.A(_04302_),
    .X(_01645_));
 sky130_fd_sc_hd__mux2_1 _08511_ (.A0(_04158_),
    .A1(net1795),
    .S(_04288_),
    .X(_04303_));
 sky130_fd_sc_hd__clkbuf_1 _08512_ (.A(_04303_),
    .X(_01646_));
 sky130_fd_sc_hd__mux2_1 _08513_ (.A0(_04160_),
    .A1(net1595),
    .S(_04288_),
    .X(_04304_));
 sky130_fd_sc_hd__clkbuf_1 _08514_ (.A(_04304_),
    .X(_01647_));
 sky130_fd_sc_hd__mux2_1 _08515_ (.A0(_04162_),
    .A1(net690),
    .S(_04288_),
    .X(_04305_));
 sky130_fd_sc_hd__clkbuf_1 _08516_ (.A(_04305_),
    .X(_01648_));
 sky130_fd_sc_hd__or3_1 _08517_ (.A(_04059_),
    .B(_02654_),
    .C(_04285_),
    .X(_04306_));
 sky130_fd_sc_hd__clkbuf_4 _08518_ (.A(_04306_),
    .X(_04307_));
 sky130_fd_sc_hd__buf_4 _08519_ (.A(_04307_),
    .X(_04308_));
 sky130_fd_sc_hd__mux2_1 _08520_ (.A0(_04125_),
    .A1(net523),
    .S(_04308_),
    .X(_04309_));
 sky130_fd_sc_hd__clkbuf_1 _08521_ (.A(_04309_),
    .X(_01649_));
 sky130_fd_sc_hd__mux2_1 _08522_ (.A0(_04134_),
    .A1(net945),
    .S(_04308_),
    .X(_04310_));
 sky130_fd_sc_hd__clkbuf_1 _08523_ (.A(_04310_),
    .X(_01650_));
 sky130_fd_sc_hd__mux2_1 _08524_ (.A0(_04136_),
    .A1(net1220),
    .S(_04308_),
    .X(_04311_));
 sky130_fd_sc_hd__clkbuf_1 _08525_ (.A(_04311_),
    .X(_01651_));
 sky130_fd_sc_hd__mux2_1 _08526_ (.A0(_04138_),
    .A1(net1052),
    .S(_04308_),
    .X(_04312_));
 sky130_fd_sc_hd__clkbuf_1 _08527_ (.A(_04312_),
    .X(_01652_));
 sky130_fd_sc_hd__mux2_1 _08528_ (.A0(_04140_),
    .A1(net447),
    .S(_04308_),
    .X(_04313_));
 sky130_fd_sc_hd__clkbuf_1 _08529_ (.A(_04313_),
    .X(_01653_));
 sky130_fd_sc_hd__mux2_1 _08530_ (.A0(_04142_),
    .A1(net482),
    .S(_04308_),
    .X(_04314_));
 sky130_fd_sc_hd__clkbuf_1 _08531_ (.A(_04314_),
    .X(_01654_));
 sky130_fd_sc_hd__mux2_1 _08532_ (.A0(_04144_),
    .A1(net1396),
    .S(_04308_),
    .X(_04315_));
 sky130_fd_sc_hd__clkbuf_1 _08533_ (.A(_04315_),
    .X(_01655_));
 sky130_fd_sc_hd__mux2_1 _08534_ (.A0(_04146_),
    .A1(net713),
    .S(_04308_),
    .X(_04316_));
 sky130_fd_sc_hd__clkbuf_1 _08535_ (.A(_04316_),
    .X(_01656_));
 sky130_fd_sc_hd__mux2_1 _08536_ (.A0(_04148_),
    .A1(net561),
    .S(_04308_),
    .X(_04317_));
 sky130_fd_sc_hd__clkbuf_1 _08537_ (.A(_04317_),
    .X(_01657_));
 sky130_fd_sc_hd__mux2_1 _08538_ (.A0(_04150_),
    .A1(net1853),
    .S(_04308_),
    .X(_04318_));
 sky130_fd_sc_hd__clkbuf_1 _08539_ (.A(_04318_),
    .X(_01658_));
 sky130_fd_sc_hd__mux2_1 _08540_ (.A0(_04152_),
    .A1(net1794),
    .S(_04307_),
    .X(_04319_));
 sky130_fd_sc_hd__clkbuf_1 _08541_ (.A(_04319_),
    .X(_01659_));
 sky130_fd_sc_hd__mux2_1 _08542_ (.A0(_04154_),
    .A1(net1179),
    .S(_04307_),
    .X(_04320_));
 sky130_fd_sc_hd__clkbuf_1 _08543_ (.A(_04320_),
    .X(_01660_));
 sky130_fd_sc_hd__mux2_1 _08544_ (.A0(_04156_),
    .A1(net1676),
    .S(_04307_),
    .X(_04321_));
 sky130_fd_sc_hd__clkbuf_1 _08545_ (.A(_04321_),
    .X(_01661_));
 sky130_fd_sc_hd__mux2_1 _08546_ (.A0(_04158_),
    .A1(net1451),
    .S(_04307_),
    .X(_04322_));
 sky130_fd_sc_hd__clkbuf_1 _08547_ (.A(_04322_),
    .X(_01662_));
 sky130_fd_sc_hd__mux2_1 _08548_ (.A0(_04160_),
    .A1(net227),
    .S(_04307_),
    .X(_04323_));
 sky130_fd_sc_hd__clkbuf_1 _08549_ (.A(_04323_),
    .X(_01663_));
 sky130_fd_sc_hd__mux2_1 _08550_ (.A0(_04162_),
    .A1(net807),
    .S(_04307_),
    .X(_04324_));
 sky130_fd_sc_hd__clkbuf_1 _08551_ (.A(_04324_),
    .X(_01664_));
 sky130_fd_sc_hd__or2_4 _08552_ (.A(_04073_),
    .B(_04128_),
    .X(_04325_));
 sky130_fd_sc_hd__or3_1 _08553_ (.A(_02702_),
    .B(_03092_),
    .C(_04325_),
    .X(_04326_));
 sky130_fd_sc_hd__clkbuf_4 _08554_ (.A(_04326_),
    .X(_04327_));
 sky130_fd_sc_hd__buf_4 _08555_ (.A(_04327_),
    .X(_04328_));
 sky130_fd_sc_hd__mux2_1 _08556_ (.A0(_04125_),
    .A1(net1053),
    .S(_04328_),
    .X(_04329_));
 sky130_fd_sc_hd__clkbuf_1 _08557_ (.A(_04329_),
    .X(_01665_));
 sky130_fd_sc_hd__mux2_1 _08558_ (.A0(_04134_),
    .A1(net563),
    .S(_04328_),
    .X(_04330_));
 sky130_fd_sc_hd__clkbuf_1 _08559_ (.A(_04330_),
    .X(_01666_));
 sky130_fd_sc_hd__mux2_1 _08560_ (.A0(_04136_),
    .A1(net1151),
    .S(_04328_),
    .X(_04331_));
 sky130_fd_sc_hd__clkbuf_1 _08561_ (.A(_04331_),
    .X(_01667_));
 sky130_fd_sc_hd__mux2_1 _08562_ (.A0(_04138_),
    .A1(net1369),
    .S(_04328_),
    .X(_04332_));
 sky130_fd_sc_hd__clkbuf_1 _08563_ (.A(_04332_),
    .X(_01668_));
 sky130_fd_sc_hd__mux2_1 _08564_ (.A0(_04140_),
    .A1(net1841),
    .S(_04328_),
    .X(_04333_));
 sky130_fd_sc_hd__clkbuf_1 _08565_ (.A(_04333_),
    .X(_01669_));
 sky130_fd_sc_hd__mux2_1 _08566_ (.A0(_04142_),
    .A1(net763),
    .S(_04328_),
    .X(_04334_));
 sky130_fd_sc_hd__clkbuf_1 _08567_ (.A(_04334_),
    .X(_01670_));
 sky130_fd_sc_hd__mux2_1 _08568_ (.A0(_04144_),
    .A1(net1605),
    .S(_04328_),
    .X(_04335_));
 sky130_fd_sc_hd__clkbuf_1 _08569_ (.A(_04335_),
    .X(_01671_));
 sky130_fd_sc_hd__mux2_1 _08570_ (.A0(_04146_),
    .A1(net1185),
    .S(_04328_),
    .X(_04336_));
 sky130_fd_sc_hd__clkbuf_1 _08571_ (.A(_04336_),
    .X(_01672_));
 sky130_fd_sc_hd__mux2_1 _08572_ (.A0(_04148_),
    .A1(net1116),
    .S(_04328_),
    .X(_04337_));
 sky130_fd_sc_hd__clkbuf_1 _08573_ (.A(_04337_),
    .X(_01673_));
 sky130_fd_sc_hd__mux2_1 _08574_ (.A0(_04150_),
    .A1(net1263),
    .S(_04328_),
    .X(_04338_));
 sky130_fd_sc_hd__clkbuf_1 _08575_ (.A(_04338_),
    .X(_01674_));
 sky130_fd_sc_hd__mux2_1 _08576_ (.A0(_04152_),
    .A1(net519),
    .S(_04327_),
    .X(_04339_));
 sky130_fd_sc_hd__clkbuf_1 _08577_ (.A(_04339_),
    .X(_01675_));
 sky130_fd_sc_hd__mux2_1 _08578_ (.A0(_04154_),
    .A1(net246),
    .S(_04327_),
    .X(_04340_));
 sky130_fd_sc_hd__clkbuf_1 _08579_ (.A(_04340_),
    .X(_01676_));
 sky130_fd_sc_hd__mux2_1 _08580_ (.A0(_04156_),
    .A1(net1684),
    .S(_04327_),
    .X(_04341_));
 sky130_fd_sc_hd__clkbuf_1 _08581_ (.A(_04341_),
    .X(_01677_));
 sky130_fd_sc_hd__mux2_1 _08582_ (.A0(_04158_),
    .A1(net744),
    .S(_04327_),
    .X(_04342_));
 sky130_fd_sc_hd__clkbuf_1 _08583_ (.A(_04342_),
    .X(_01678_));
 sky130_fd_sc_hd__mux2_1 _08584_ (.A0(_04160_),
    .A1(net1344),
    .S(_04327_),
    .X(_04343_));
 sky130_fd_sc_hd__clkbuf_1 _08585_ (.A(_04343_),
    .X(_01679_));
 sky130_fd_sc_hd__mux2_1 _08586_ (.A0(_04162_),
    .A1(net322),
    .S(_04327_),
    .X(_04344_));
 sky130_fd_sc_hd__clkbuf_1 _08587_ (.A(_04344_),
    .X(_01680_));
 sky130_fd_sc_hd__or3_1 _08588_ (.A(_04059_),
    .B(_03092_),
    .C(_04325_),
    .X(_04345_));
 sky130_fd_sc_hd__clkbuf_4 _08589_ (.A(_04345_),
    .X(_04346_));
 sky130_fd_sc_hd__buf_4 _08590_ (.A(_04346_),
    .X(_04347_));
 sky130_fd_sc_hd__mux2_1 _08591_ (.A0(_04125_),
    .A1(net837),
    .S(_04347_),
    .X(_04348_));
 sky130_fd_sc_hd__clkbuf_1 _08592_ (.A(_04348_),
    .X(_01681_));
 sky130_fd_sc_hd__mux2_1 _08593_ (.A0(_04134_),
    .A1(net1255),
    .S(_04347_),
    .X(_04349_));
 sky130_fd_sc_hd__clkbuf_1 _08594_ (.A(_04349_),
    .X(_01682_));
 sky130_fd_sc_hd__mux2_1 _08595_ (.A0(_04136_),
    .A1(net1009),
    .S(_04347_),
    .X(_04350_));
 sky130_fd_sc_hd__clkbuf_1 _08596_ (.A(_04350_),
    .X(_01683_));
 sky130_fd_sc_hd__mux2_1 _08597_ (.A0(_04138_),
    .A1(net1021),
    .S(_04347_),
    .X(_04351_));
 sky130_fd_sc_hd__clkbuf_1 _08598_ (.A(_04351_),
    .X(_01684_));
 sky130_fd_sc_hd__mux2_1 _08599_ (.A0(_04140_),
    .A1(net789),
    .S(_04347_),
    .X(_04352_));
 sky130_fd_sc_hd__clkbuf_1 _08600_ (.A(_04352_),
    .X(_01685_));
 sky130_fd_sc_hd__mux2_1 _08601_ (.A0(_04142_),
    .A1(net1478),
    .S(_04347_),
    .X(_04353_));
 sky130_fd_sc_hd__clkbuf_1 _08602_ (.A(_04353_),
    .X(_01686_));
 sky130_fd_sc_hd__mux2_1 _08603_ (.A0(_04144_),
    .A1(net605),
    .S(_04347_),
    .X(_04354_));
 sky130_fd_sc_hd__clkbuf_1 _08604_ (.A(_04354_),
    .X(_01687_));
 sky130_fd_sc_hd__mux2_1 _08605_ (.A0(_04146_),
    .A1(net633),
    .S(_04347_),
    .X(_04355_));
 sky130_fd_sc_hd__clkbuf_1 _08606_ (.A(_04355_),
    .X(_01688_));
 sky130_fd_sc_hd__mux2_1 _08607_ (.A0(_04148_),
    .A1(net778),
    .S(_04347_),
    .X(_04356_));
 sky130_fd_sc_hd__clkbuf_1 _08608_ (.A(_04356_),
    .X(_01689_));
 sky130_fd_sc_hd__mux2_1 _08609_ (.A0(_04150_),
    .A1(net924),
    .S(_04347_),
    .X(_04357_));
 sky130_fd_sc_hd__clkbuf_1 _08610_ (.A(_04357_),
    .X(_01690_));
 sky130_fd_sc_hd__mux2_1 _08611_ (.A0(_04152_),
    .A1(net1376),
    .S(_04346_),
    .X(_04358_));
 sky130_fd_sc_hd__clkbuf_1 _08612_ (.A(_04358_),
    .X(_01691_));
 sky130_fd_sc_hd__mux2_1 _08613_ (.A0(_04154_),
    .A1(net1539),
    .S(_04346_),
    .X(_04359_));
 sky130_fd_sc_hd__clkbuf_1 _08614_ (.A(_04359_),
    .X(_01692_));
 sky130_fd_sc_hd__mux2_1 _08615_ (.A0(_04156_),
    .A1(net1031),
    .S(_04346_),
    .X(_04360_));
 sky130_fd_sc_hd__clkbuf_1 _08616_ (.A(_04360_),
    .X(_01693_));
 sky130_fd_sc_hd__mux2_1 _08617_ (.A0(_04158_),
    .A1(net1203),
    .S(_04346_),
    .X(_04361_));
 sky130_fd_sc_hd__clkbuf_1 _08618_ (.A(_04361_),
    .X(_01694_));
 sky130_fd_sc_hd__mux2_1 _08619_ (.A0(_04160_),
    .A1(net1370),
    .S(_04346_),
    .X(_04362_));
 sky130_fd_sc_hd__clkbuf_1 _08620_ (.A(_04362_),
    .X(_01695_));
 sky130_fd_sc_hd__mux2_1 _08621_ (.A0(_04162_),
    .A1(net307),
    .S(_04346_),
    .X(_04363_));
 sky130_fd_sc_hd__clkbuf_1 _08622_ (.A(_04363_),
    .X(_01696_));
 sky130_fd_sc_hd__or3_1 _08623_ (.A(_02645_),
    .B(_02617_),
    .C(_02483_),
    .X(_04364_));
 sky130_fd_sc_hd__buf_12 _08624_ (.A(_04364_),
    .X(_04365_));
 sky130_fd_sc_hd__or3_1 _08625_ (.A(net5),
    .B(net6),
    .C(_04074_),
    .X(_04366_));
 sky130_fd_sc_hd__clkbuf_4 _08626_ (.A(_04366_),
    .X(_04367_));
 sky130_fd_sc_hd__buf_12 _08627_ (.A(_04367_),
    .X(_04368_));
 sky130_fd_sc_hd__nor2_4 _08628_ (.A(_04365_),
    .B(_04368_),
    .Y(_04369_));
 sky130_fd_sc_hd__buf_4 _08629_ (.A(_04369_),
    .X(_04370_));
 sky130_fd_sc_hd__mux2_1 _08630_ (.A0(net1819),
    .A1(_04070_),
    .S(_04370_),
    .X(_04371_));
 sky130_fd_sc_hd__clkbuf_1 _08631_ (.A(_04371_),
    .X(_01697_));
 sky130_fd_sc_hd__mux2_1 _08632_ (.A0(net293),
    .A1(_04081_),
    .S(_04370_),
    .X(_04372_));
 sky130_fd_sc_hd__clkbuf_1 _08633_ (.A(_04372_),
    .X(_01698_));
 sky130_fd_sc_hd__mux2_1 _08634_ (.A0(net197),
    .A1(_04084_),
    .S(_04370_),
    .X(_04373_));
 sky130_fd_sc_hd__clkbuf_1 _08635_ (.A(_04373_),
    .X(_01699_));
 sky130_fd_sc_hd__mux2_1 _08636_ (.A0(net152),
    .A1(_04087_),
    .S(_04370_),
    .X(_04374_));
 sky130_fd_sc_hd__clkbuf_1 _08637_ (.A(_04374_),
    .X(_01700_));
 sky130_fd_sc_hd__mux2_1 _08638_ (.A0(net100),
    .A1(_04090_),
    .S(_04370_),
    .X(_04375_));
 sky130_fd_sc_hd__clkbuf_1 _08639_ (.A(_04375_),
    .X(_01701_));
 sky130_fd_sc_hd__mux2_1 _08640_ (.A0(net44),
    .A1(_04093_),
    .S(_04370_),
    .X(_04376_));
 sky130_fd_sc_hd__clkbuf_1 _08641_ (.A(_04376_),
    .X(_01702_));
 sky130_fd_sc_hd__mux2_1 _08642_ (.A0(net92),
    .A1(_04096_),
    .S(_04370_),
    .X(_04377_));
 sky130_fd_sc_hd__clkbuf_1 _08643_ (.A(_04377_),
    .X(_01703_));
 sky130_fd_sc_hd__mux2_1 _08644_ (.A0(net399),
    .A1(_04099_),
    .S(_04370_),
    .X(_04378_));
 sky130_fd_sc_hd__clkbuf_1 _08645_ (.A(_04378_),
    .X(_01704_));
 sky130_fd_sc_hd__mux2_1 _08646_ (.A0(net60),
    .A1(_04102_),
    .S(_04370_),
    .X(_04379_));
 sky130_fd_sc_hd__clkbuf_1 _08647_ (.A(_04379_),
    .X(_01705_));
 sky130_fd_sc_hd__mux2_1 _08648_ (.A0(net140),
    .A1(_04105_),
    .S(_04370_),
    .X(_04380_));
 sky130_fd_sc_hd__clkbuf_1 _08649_ (.A(_04380_),
    .X(_01706_));
 sky130_fd_sc_hd__mux2_1 _08650_ (.A0(net124),
    .A1(_04108_),
    .S(_04369_),
    .X(_04381_));
 sky130_fd_sc_hd__clkbuf_1 _08651_ (.A(_04381_),
    .X(_01707_));
 sky130_fd_sc_hd__mux2_1 _08652_ (.A0(net134),
    .A1(_04111_),
    .S(_04369_),
    .X(_04382_));
 sky130_fd_sc_hd__clkbuf_1 _08653_ (.A(_04382_),
    .X(_01708_));
 sky130_fd_sc_hd__mux2_1 _08654_ (.A0(net73),
    .A1(_04114_),
    .S(_04369_),
    .X(_04383_));
 sky130_fd_sc_hd__clkbuf_1 _08655_ (.A(_04383_),
    .X(_01709_));
 sky130_fd_sc_hd__mux2_1 _08656_ (.A0(net42),
    .A1(_04117_),
    .S(_04369_),
    .X(_04384_));
 sky130_fd_sc_hd__clkbuf_1 _08657_ (.A(_04384_),
    .X(_01710_));
 sky130_fd_sc_hd__mux2_1 _08658_ (.A0(net1114),
    .A1(_04120_),
    .S(_04369_),
    .X(_04385_));
 sky130_fd_sc_hd__clkbuf_1 _08659_ (.A(_04385_),
    .X(_01711_));
 sky130_fd_sc_hd__mux2_1 _08660_ (.A0(net324),
    .A1(_04123_),
    .S(_04369_),
    .X(_04386_));
 sky130_fd_sc_hd__clkbuf_1 _08661_ (.A(_04386_),
    .X(_01712_));
 sky130_fd_sc_hd__or3_1 _08662_ (.A(_04059_),
    .B(_02654_),
    .C(_04367_),
    .X(_04387_));
 sky130_fd_sc_hd__clkbuf_4 _08663_ (.A(_04387_),
    .X(_04388_));
 sky130_fd_sc_hd__buf_4 _08664_ (.A(_04388_),
    .X(_04389_));
 sky130_fd_sc_hd__mux2_1 _08665_ (.A0(_04125_),
    .A1(net1348),
    .S(_04389_),
    .X(_04390_));
 sky130_fd_sc_hd__clkbuf_1 _08666_ (.A(_04390_),
    .X(_01713_));
 sky130_fd_sc_hd__mux2_1 _08667_ (.A0(_04134_),
    .A1(net554),
    .S(_04389_),
    .X(_04391_));
 sky130_fd_sc_hd__clkbuf_1 _08668_ (.A(_04391_),
    .X(_01714_));
 sky130_fd_sc_hd__mux2_1 _08669_ (.A0(_04136_),
    .A1(net1487),
    .S(_04389_),
    .X(_04392_));
 sky130_fd_sc_hd__clkbuf_1 _08670_ (.A(_04392_),
    .X(_01715_));
 sky130_fd_sc_hd__mux2_1 _08671_ (.A0(_04138_),
    .A1(net1325),
    .S(_04389_),
    .X(_04393_));
 sky130_fd_sc_hd__clkbuf_1 _08672_ (.A(_04393_),
    .X(_01716_));
 sky130_fd_sc_hd__mux2_1 _08673_ (.A0(_04140_),
    .A1(net1644),
    .S(_04389_),
    .X(_04394_));
 sky130_fd_sc_hd__clkbuf_1 _08674_ (.A(_04394_),
    .X(_01717_));
 sky130_fd_sc_hd__mux2_1 _08675_ (.A0(_04142_),
    .A1(net1025),
    .S(_04389_),
    .X(_04395_));
 sky130_fd_sc_hd__clkbuf_1 _08676_ (.A(_04395_),
    .X(_01718_));
 sky130_fd_sc_hd__mux2_1 _08677_ (.A0(_04144_),
    .A1(net1311),
    .S(_04389_),
    .X(_04396_));
 sky130_fd_sc_hd__clkbuf_1 _08678_ (.A(_04396_),
    .X(_01719_));
 sky130_fd_sc_hd__mux2_1 _08679_ (.A0(_04146_),
    .A1(net1682),
    .S(_04389_),
    .X(_04397_));
 sky130_fd_sc_hd__clkbuf_1 _08680_ (.A(_04397_),
    .X(_01720_));
 sky130_fd_sc_hd__mux2_1 _08681_ (.A0(_04148_),
    .A1(net1518),
    .S(_04389_),
    .X(_04398_));
 sky130_fd_sc_hd__clkbuf_1 _08682_ (.A(_04398_),
    .X(_01721_));
 sky130_fd_sc_hd__mux2_1 _08683_ (.A0(_04150_),
    .A1(net1104),
    .S(_04389_),
    .X(_04399_));
 sky130_fd_sc_hd__clkbuf_1 _08684_ (.A(_04399_),
    .X(_01722_));
 sky130_fd_sc_hd__mux2_1 _08685_ (.A0(_04152_),
    .A1(net1880),
    .S(_04388_),
    .X(_04400_));
 sky130_fd_sc_hd__clkbuf_1 _08686_ (.A(_04400_),
    .X(_01723_));
 sky130_fd_sc_hd__mux2_1 _08687_ (.A0(_04154_),
    .A1(net1960),
    .S(_04388_),
    .X(_04401_));
 sky130_fd_sc_hd__clkbuf_1 _08688_ (.A(_04401_),
    .X(_01724_));
 sky130_fd_sc_hd__mux2_1 _08689_ (.A0(_04156_),
    .A1(net952),
    .S(_04388_),
    .X(_04402_));
 sky130_fd_sc_hd__clkbuf_1 _08690_ (.A(_04402_),
    .X(_01725_));
 sky130_fd_sc_hd__mux2_1 _08691_ (.A0(_04158_),
    .A1(net1790),
    .S(_04388_),
    .X(_04403_));
 sky130_fd_sc_hd__clkbuf_1 _08692_ (.A(_04403_),
    .X(_01726_));
 sky130_fd_sc_hd__mux2_1 _08693_ (.A0(_04160_),
    .A1(net1871),
    .S(_04388_),
    .X(_04404_));
 sky130_fd_sc_hd__clkbuf_1 _08694_ (.A(_04404_),
    .X(_01727_));
 sky130_fd_sc_hd__mux2_1 _08695_ (.A0(_04162_),
    .A1(net1593),
    .S(_04388_),
    .X(_04405_));
 sky130_fd_sc_hd__clkbuf_1 _08696_ (.A(_04405_),
    .X(_01728_));
 sky130_fd_sc_hd__buf_6 _08697_ (.A(_04069_),
    .X(_04406_));
 sky130_fd_sc_hd__and3b_1 _08698_ (.A_N(_02749_),
    .B(_02674_),
    .C(_02422_),
    .X(_04407_));
 sky130_fd_sc_hd__buf_12 _08699_ (.A(_04407_),
    .X(_04408_));
 sky130_fd_sc_hd__nand2b_4 _08700_ (.A_N(_04367_),
    .B(_04408_),
    .Y(_04409_));
 sky130_fd_sc_hd__buf_4 _08701_ (.A(_04409_),
    .X(_04410_));
 sky130_fd_sc_hd__mux2_1 _08702_ (.A0(_04406_),
    .A1(net1588),
    .S(_04410_),
    .X(_04411_));
 sky130_fd_sc_hd__clkbuf_1 _08703_ (.A(_04411_),
    .X(_01729_));
 sky130_fd_sc_hd__buf_6 _08704_ (.A(_04080_),
    .X(_04412_));
 sky130_fd_sc_hd__mux2_1 _08705_ (.A0(_04412_),
    .A1(net1308),
    .S(_04410_),
    .X(_04413_));
 sky130_fd_sc_hd__clkbuf_1 _08706_ (.A(_04413_),
    .X(_01730_));
 sky130_fd_sc_hd__buf_6 _08707_ (.A(_04083_),
    .X(_04414_));
 sky130_fd_sc_hd__mux2_1 _08708_ (.A0(_04414_),
    .A1(net1776),
    .S(_04410_),
    .X(_04415_));
 sky130_fd_sc_hd__clkbuf_1 _08709_ (.A(_04415_),
    .X(_01731_));
 sky130_fd_sc_hd__buf_6 _08710_ (.A(_04086_),
    .X(_04416_));
 sky130_fd_sc_hd__mux2_1 _08711_ (.A0(_04416_),
    .A1(net1834),
    .S(_04410_),
    .X(_04417_));
 sky130_fd_sc_hd__clkbuf_1 _08712_ (.A(_04417_),
    .X(_01732_));
 sky130_fd_sc_hd__buf_8 _08713_ (.A(_04089_),
    .X(_04418_));
 sky130_fd_sc_hd__mux2_1 _08714_ (.A0(_04418_),
    .A1(net1951),
    .S(_04410_),
    .X(_04419_));
 sky130_fd_sc_hd__clkbuf_1 _08715_ (.A(_04419_),
    .X(_01733_));
 sky130_fd_sc_hd__buf_6 _08716_ (.A(_04092_),
    .X(_04420_));
 sky130_fd_sc_hd__mux2_1 _08717_ (.A0(_04420_),
    .A1(net333),
    .S(_04410_),
    .X(_04421_));
 sky130_fd_sc_hd__clkbuf_1 _08718_ (.A(_04421_),
    .X(_01734_));
 sky130_fd_sc_hd__buf_8 _08719_ (.A(_04095_),
    .X(_04422_));
 sky130_fd_sc_hd__mux2_1 _08720_ (.A0(_04422_),
    .A1(net1406),
    .S(_04410_),
    .X(_04423_));
 sky130_fd_sc_hd__clkbuf_1 _08721_ (.A(_04423_),
    .X(_01735_));
 sky130_fd_sc_hd__buf_8 _08722_ (.A(_04098_),
    .X(_04424_));
 sky130_fd_sc_hd__mux2_1 _08723_ (.A0(_04424_),
    .A1(net1616),
    .S(_04410_),
    .X(_04425_));
 sky130_fd_sc_hd__clkbuf_1 _08724_ (.A(_04425_),
    .X(_01736_));
 sky130_fd_sc_hd__buf_8 _08725_ (.A(_04101_),
    .X(_04426_));
 sky130_fd_sc_hd__mux2_1 _08726_ (.A0(_04426_),
    .A1(net1637),
    .S(_04410_),
    .X(_04427_));
 sky130_fd_sc_hd__clkbuf_1 _08727_ (.A(_04427_),
    .X(_01737_));
 sky130_fd_sc_hd__buf_8 _08728_ (.A(_04104_),
    .X(_04428_));
 sky130_fd_sc_hd__mux2_1 _08729_ (.A0(_04428_),
    .A1(net1629),
    .S(_04410_),
    .X(_04429_));
 sky130_fd_sc_hd__clkbuf_1 _08730_ (.A(_04429_),
    .X(_01738_));
 sky130_fd_sc_hd__buf_8 _08731_ (.A(_04107_),
    .X(_04430_));
 sky130_fd_sc_hd__mux2_1 _08732_ (.A0(_04430_),
    .A1(net1385),
    .S(_04409_),
    .X(_04431_));
 sky130_fd_sc_hd__clkbuf_1 _08733_ (.A(_04431_),
    .X(_01739_));
 sky130_fd_sc_hd__buf_8 _08734_ (.A(_04110_),
    .X(_04432_));
 sky130_fd_sc_hd__mux2_1 _08735_ (.A0(_04432_),
    .A1(net1827),
    .S(_04409_),
    .X(_04433_));
 sky130_fd_sc_hd__clkbuf_1 _08736_ (.A(_04433_),
    .X(_01740_));
 sky130_fd_sc_hd__buf_8 _08737_ (.A(_04113_),
    .X(_04434_));
 sky130_fd_sc_hd__mux2_1 _08738_ (.A0(_04434_),
    .A1(net1564),
    .S(_04409_),
    .X(_04435_));
 sky130_fd_sc_hd__clkbuf_1 _08739_ (.A(_04435_),
    .X(_01741_));
 sky130_fd_sc_hd__buf_6 _08740_ (.A(_04116_),
    .X(_04436_));
 sky130_fd_sc_hd__mux2_1 _08741_ (.A0(_04436_),
    .A1(net1367),
    .S(_04409_),
    .X(_04437_));
 sky130_fd_sc_hd__clkbuf_1 _08742_ (.A(_04437_),
    .X(_01742_));
 sky130_fd_sc_hd__buf_8 _08743_ (.A(_04119_),
    .X(_04438_));
 sky130_fd_sc_hd__mux2_1 _08744_ (.A0(_04438_),
    .A1(net1740),
    .S(_04409_),
    .X(_04439_));
 sky130_fd_sc_hd__clkbuf_1 _08745_ (.A(_04439_),
    .X(_01743_));
 sky130_fd_sc_hd__buf_8 _08746_ (.A(_04122_),
    .X(_04440_));
 sky130_fd_sc_hd__mux2_1 _08747_ (.A0(_04440_),
    .A1(net1948),
    .S(_04409_),
    .X(_04441_));
 sky130_fd_sc_hd__clkbuf_1 _08748_ (.A(_04441_),
    .X(_01744_));
 sky130_fd_sc_hd__nor3_4 _08749_ (.A(_02485_),
    .B(_02666_),
    .C(_04367_),
    .Y(_04442_));
 sky130_fd_sc_hd__buf_4 _08750_ (.A(_04442_),
    .X(_04443_));
 sky130_fd_sc_hd__mux2_1 _08751_ (.A0(net2001),
    .A1(_04070_),
    .S(_04443_),
    .X(_04444_));
 sky130_fd_sc_hd__clkbuf_1 _08752_ (.A(_04444_),
    .X(_01745_));
 sky130_fd_sc_hd__mux2_1 _08753_ (.A0(net660),
    .A1(_04081_),
    .S(_04443_),
    .X(_04445_));
 sky130_fd_sc_hd__clkbuf_1 _08754_ (.A(_04445_),
    .X(_01746_));
 sky130_fd_sc_hd__mux2_1 _08755_ (.A0(net1230),
    .A1(_04084_),
    .S(_04443_),
    .X(_04446_));
 sky130_fd_sc_hd__clkbuf_1 _08756_ (.A(_04446_),
    .X(_01747_));
 sky130_fd_sc_hd__mux2_1 _08757_ (.A0(net1444),
    .A1(_04087_),
    .S(_04443_),
    .X(_04447_));
 sky130_fd_sc_hd__clkbuf_1 _08758_ (.A(_04447_),
    .X(_01748_));
 sky130_fd_sc_hd__mux2_1 _08759_ (.A0(net1010),
    .A1(_04090_),
    .S(_04443_),
    .X(_04448_));
 sky130_fd_sc_hd__clkbuf_1 _08760_ (.A(_04448_),
    .X(_01749_));
 sky130_fd_sc_hd__mux2_1 _08761_ (.A0(net527),
    .A1(_04093_),
    .S(_04443_),
    .X(_04449_));
 sky130_fd_sc_hd__clkbuf_1 _08762_ (.A(_04449_),
    .X(_01750_));
 sky130_fd_sc_hd__mux2_1 _08763_ (.A0(net1079),
    .A1(_04096_),
    .S(_04443_),
    .X(_04450_));
 sky130_fd_sc_hd__clkbuf_1 _08764_ (.A(_04450_),
    .X(_01751_));
 sky130_fd_sc_hd__mux2_1 _08765_ (.A0(net897),
    .A1(_04099_),
    .S(_04443_),
    .X(_04451_));
 sky130_fd_sc_hd__clkbuf_1 _08766_ (.A(_04451_),
    .X(_01752_));
 sky130_fd_sc_hd__mux2_1 _08767_ (.A0(net1771),
    .A1(_04102_),
    .S(_04443_),
    .X(_04452_));
 sky130_fd_sc_hd__clkbuf_1 _08768_ (.A(_04452_),
    .X(_01753_));
 sky130_fd_sc_hd__mux2_1 _08769_ (.A0(net810),
    .A1(_04105_),
    .S(_04443_),
    .X(_04453_));
 sky130_fd_sc_hd__clkbuf_1 _08770_ (.A(_04453_),
    .X(_01754_));
 sky130_fd_sc_hd__mux2_1 _08771_ (.A0(net224),
    .A1(_04108_),
    .S(_04442_),
    .X(_04454_));
 sky130_fd_sc_hd__clkbuf_1 _08772_ (.A(_04454_),
    .X(_01755_));
 sky130_fd_sc_hd__mux2_1 _08773_ (.A0(net803),
    .A1(_04111_),
    .S(_04442_),
    .X(_04455_));
 sky130_fd_sc_hd__clkbuf_1 _08774_ (.A(_04455_),
    .X(_01756_));
 sky130_fd_sc_hd__mux2_1 _08775_ (.A0(net830),
    .A1(_04114_),
    .S(_04442_),
    .X(_04456_));
 sky130_fd_sc_hd__clkbuf_1 _08776_ (.A(_04456_),
    .X(_01757_));
 sky130_fd_sc_hd__mux2_1 _08777_ (.A0(net56),
    .A1(_04117_),
    .S(_04442_),
    .X(_04457_));
 sky130_fd_sc_hd__clkbuf_1 _08778_ (.A(_04457_),
    .X(_01758_));
 sky130_fd_sc_hd__mux2_1 _08779_ (.A0(net1291),
    .A1(_04120_),
    .S(_04442_),
    .X(_04458_));
 sky130_fd_sc_hd__clkbuf_1 _08780_ (.A(_04458_),
    .X(_01759_));
 sky130_fd_sc_hd__mux2_1 _08781_ (.A0(net1164),
    .A1(_04123_),
    .S(_04442_),
    .X(_04459_));
 sky130_fd_sc_hd__clkbuf_1 _08782_ (.A(_04459_),
    .X(_01760_));
 sky130_fd_sc_hd__or3_1 _08783_ (.A(_02656_),
    .B(_02492_),
    .C(_02495_),
    .X(_04460_));
 sky130_fd_sc_hd__buf_12 _08784_ (.A(_04460_),
    .X(_04461_));
 sky130_fd_sc_hd__nor2_4 _08785_ (.A(_04227_),
    .B(_04461_),
    .Y(_04462_));
 sky130_fd_sc_hd__buf_4 _08786_ (.A(_04462_),
    .X(_04463_));
 sky130_fd_sc_hd__mux2_1 _08787_ (.A0(net1094),
    .A1(_04070_),
    .S(_04463_),
    .X(_04464_));
 sky130_fd_sc_hd__clkbuf_1 _08788_ (.A(_04464_),
    .X(_01761_));
 sky130_fd_sc_hd__mux2_1 _08789_ (.A0(net1330),
    .A1(_04081_),
    .S(_04463_),
    .X(_04465_));
 sky130_fd_sc_hd__clkbuf_1 _08790_ (.A(_04465_),
    .X(_01762_));
 sky130_fd_sc_hd__mux2_1 _08791_ (.A0(net670),
    .A1(_04084_),
    .S(_04463_),
    .X(_04466_));
 sky130_fd_sc_hd__clkbuf_1 _08792_ (.A(_04466_),
    .X(_01763_));
 sky130_fd_sc_hd__mux2_1 _08793_ (.A0(net1219),
    .A1(_04087_),
    .S(_04463_),
    .X(_04467_));
 sky130_fd_sc_hd__clkbuf_1 _08794_ (.A(_04467_),
    .X(_01764_));
 sky130_fd_sc_hd__mux2_1 _08795_ (.A0(net271),
    .A1(_04090_),
    .S(_04463_),
    .X(_04468_));
 sky130_fd_sc_hd__clkbuf_1 _08796_ (.A(_04468_),
    .X(_01765_));
 sky130_fd_sc_hd__mux2_1 _08797_ (.A0(net987),
    .A1(_04093_),
    .S(_04463_),
    .X(_04469_));
 sky130_fd_sc_hd__clkbuf_1 _08798_ (.A(_04469_),
    .X(_01766_));
 sky130_fd_sc_hd__mux2_1 _08799_ (.A0(net1398),
    .A1(_04096_),
    .S(_04463_),
    .X(_04470_));
 sky130_fd_sc_hd__clkbuf_1 _08800_ (.A(_04470_),
    .X(_01767_));
 sky130_fd_sc_hd__mux2_1 _08801_ (.A0(net680),
    .A1(_04099_),
    .S(_04463_),
    .X(_04471_));
 sky130_fd_sc_hd__clkbuf_1 _08802_ (.A(_04471_),
    .X(_01768_));
 sky130_fd_sc_hd__mux2_1 _08803_ (.A0(net1015),
    .A1(_04102_),
    .S(_04463_),
    .X(_04472_));
 sky130_fd_sc_hd__clkbuf_1 _08804_ (.A(_04472_),
    .X(_01769_));
 sky130_fd_sc_hd__mux2_1 _08805_ (.A0(net1022),
    .A1(_04105_),
    .S(_04463_),
    .X(_04473_));
 sky130_fd_sc_hd__clkbuf_1 _08806_ (.A(_04473_),
    .X(_01770_));
 sky130_fd_sc_hd__mux2_1 _08807_ (.A0(net468),
    .A1(_04108_),
    .S(_04462_),
    .X(_04474_));
 sky130_fd_sc_hd__clkbuf_1 _08808_ (.A(_04474_),
    .X(_01771_));
 sky130_fd_sc_hd__mux2_1 _08809_ (.A0(net655),
    .A1(_04111_),
    .S(_04462_),
    .X(_04475_));
 sky130_fd_sc_hd__clkbuf_1 _08810_ (.A(_04475_),
    .X(_01772_));
 sky130_fd_sc_hd__mux2_1 _08811_ (.A0(net1186),
    .A1(_04114_),
    .S(_04462_),
    .X(_04476_));
 sky130_fd_sc_hd__clkbuf_1 _08812_ (.A(_04476_),
    .X(_01773_));
 sky130_fd_sc_hd__mux2_1 _08813_ (.A0(net1138),
    .A1(_04117_),
    .S(_04462_),
    .X(_04477_));
 sky130_fd_sc_hd__clkbuf_1 _08814_ (.A(_04477_),
    .X(_01774_));
 sky130_fd_sc_hd__mux2_1 _08815_ (.A0(net961),
    .A1(_04120_),
    .S(_04462_),
    .X(_04478_));
 sky130_fd_sc_hd__clkbuf_1 _08816_ (.A(_04478_),
    .X(_01775_));
 sky130_fd_sc_hd__mux2_1 _08817_ (.A0(net1438),
    .A1(_04123_),
    .S(_04462_),
    .X(_04479_));
 sky130_fd_sc_hd__clkbuf_1 _08818_ (.A(_04479_),
    .X(_01776_));
 sky130_fd_sc_hd__nor2_4 _08819_ (.A(_04072_),
    .B(_04227_),
    .Y(_04480_));
 sky130_fd_sc_hd__clkbuf_8 _08820_ (.A(_04480_),
    .X(_04481_));
 sky130_fd_sc_hd__mux2_1 _08821_ (.A0(net1355),
    .A1(_04070_),
    .S(_04481_),
    .X(_04482_));
 sky130_fd_sc_hd__clkbuf_1 _08822_ (.A(_04482_),
    .X(_01777_));
 sky130_fd_sc_hd__mux2_1 _08823_ (.A0(net852),
    .A1(_04081_),
    .S(_04481_),
    .X(_04483_));
 sky130_fd_sc_hd__clkbuf_1 _08824_ (.A(_04483_),
    .X(_01778_));
 sky130_fd_sc_hd__mux2_1 _08825_ (.A0(net1029),
    .A1(_04084_),
    .S(_04481_),
    .X(_04484_));
 sky130_fd_sc_hd__clkbuf_1 _08826_ (.A(_04484_),
    .X(_01779_));
 sky130_fd_sc_hd__mux2_1 _08827_ (.A0(net1182),
    .A1(_04087_),
    .S(_04481_),
    .X(_04485_));
 sky130_fd_sc_hd__clkbuf_1 _08828_ (.A(_04485_),
    .X(_01780_));
 sky130_fd_sc_hd__mux2_1 _08829_ (.A0(net1645),
    .A1(_04090_),
    .S(_04481_),
    .X(_04486_));
 sky130_fd_sc_hd__clkbuf_1 _08830_ (.A(_04486_),
    .X(_01781_));
 sky130_fd_sc_hd__mux2_1 _08831_ (.A0(net1498),
    .A1(_04093_),
    .S(_04481_),
    .X(_04487_));
 sky130_fd_sc_hd__clkbuf_1 _08832_ (.A(_04487_),
    .X(_01782_));
 sky130_fd_sc_hd__mux2_1 _08833_ (.A0(net654),
    .A1(_04096_),
    .S(_04481_),
    .X(_04488_));
 sky130_fd_sc_hd__clkbuf_1 _08834_ (.A(_04488_),
    .X(_01783_));
 sky130_fd_sc_hd__mux2_1 _08835_ (.A0(net1049),
    .A1(_04099_),
    .S(_04481_),
    .X(_04489_));
 sky130_fd_sc_hd__clkbuf_1 _08836_ (.A(_04489_),
    .X(_01784_));
 sky130_fd_sc_hd__mux2_1 _08837_ (.A0(net535),
    .A1(_04102_),
    .S(_04481_),
    .X(_04490_));
 sky130_fd_sc_hd__clkbuf_1 _08838_ (.A(_04490_),
    .X(_01785_));
 sky130_fd_sc_hd__mux2_1 _08839_ (.A0(net1649),
    .A1(_04105_),
    .S(_04481_),
    .X(_04491_));
 sky130_fd_sc_hd__clkbuf_1 _08840_ (.A(_04491_),
    .X(_01786_));
 sky130_fd_sc_hd__mux2_1 _08841_ (.A0(net306),
    .A1(_04108_),
    .S(_04480_),
    .X(_04492_));
 sky130_fd_sc_hd__clkbuf_1 _08842_ (.A(_04492_),
    .X(_01787_));
 sky130_fd_sc_hd__mux2_1 _08843_ (.A0(net1173),
    .A1(_04111_),
    .S(_04480_),
    .X(_04493_));
 sky130_fd_sc_hd__clkbuf_1 _08844_ (.A(_04493_),
    .X(_01788_));
 sky130_fd_sc_hd__mux2_1 _08845_ (.A0(net936),
    .A1(_04114_),
    .S(_04480_),
    .X(_04494_));
 sky130_fd_sc_hd__clkbuf_1 _08846_ (.A(_04494_),
    .X(_01789_));
 sky130_fd_sc_hd__mux2_1 _08847_ (.A0(net1735),
    .A1(_04117_),
    .S(_04480_),
    .X(_04495_));
 sky130_fd_sc_hd__clkbuf_1 _08848_ (.A(_04495_),
    .X(_01790_));
 sky130_fd_sc_hd__mux2_1 _08849_ (.A0(net2011),
    .A1(_04120_),
    .S(_04480_),
    .X(_04496_));
 sky130_fd_sc_hd__clkbuf_1 _08850_ (.A(_04496_),
    .X(_01791_));
 sky130_fd_sc_hd__mux2_1 _08851_ (.A0(net873),
    .A1(_04123_),
    .S(_04480_),
    .X(_04497_));
 sky130_fd_sc_hd__clkbuf_1 _08852_ (.A(_04497_),
    .X(_01792_));
 sky130_fd_sc_hd__buf_6 _08853_ (.A(net8),
    .X(_04498_));
 sky130_fd_sc_hd__clkbuf_4 _08854_ (.A(_04498_),
    .X(_04499_));
 sky130_fd_sc_hd__or3b_1 _08855_ (.A(_02495_),
    .B(_02681_),
    .C_N(_02682_),
    .X(_04500_));
 sky130_fd_sc_hd__buf_12 _08856_ (.A(_04500_),
    .X(_04501_));
 sky130_fd_sc_hd__nor2_4 _08857_ (.A(_04227_),
    .B(_04501_),
    .Y(_04502_));
 sky130_fd_sc_hd__buf_4 _08858_ (.A(_04502_),
    .X(_04503_));
 sky130_fd_sc_hd__mux2_1 _08859_ (.A0(net460),
    .A1(_04499_),
    .S(_04503_),
    .X(_04504_));
 sky130_fd_sc_hd__clkbuf_1 _08860_ (.A(_04504_),
    .X(_01793_));
 sky130_fd_sc_hd__buf_4 _08861_ (.A(net15),
    .X(_04505_));
 sky130_fd_sc_hd__clkbuf_4 _08862_ (.A(_04505_),
    .X(_04506_));
 sky130_fd_sc_hd__mux2_1 _08863_ (.A0(net902),
    .A1(_04506_),
    .S(_04503_),
    .X(_04507_));
 sky130_fd_sc_hd__clkbuf_1 _08864_ (.A(_04507_),
    .X(_01794_));
 sky130_fd_sc_hd__buf_6 _08865_ (.A(net16),
    .X(_04508_));
 sky130_fd_sc_hd__buf_4 _08866_ (.A(_04508_),
    .X(_04509_));
 sky130_fd_sc_hd__mux2_1 _08867_ (.A0(net828),
    .A1(_04509_),
    .S(_04503_),
    .X(_04510_));
 sky130_fd_sc_hd__clkbuf_1 _08868_ (.A(_04510_),
    .X(_01795_));
 sky130_fd_sc_hd__buf_6 _08869_ (.A(net17),
    .X(_04511_));
 sky130_fd_sc_hd__clkbuf_4 _08870_ (.A(_04511_),
    .X(_04512_));
 sky130_fd_sc_hd__mux2_1 _08871_ (.A0(net1058),
    .A1(_04512_),
    .S(_04503_),
    .X(_04513_));
 sky130_fd_sc_hd__clkbuf_1 _08872_ (.A(_04513_),
    .X(_01796_));
 sky130_fd_sc_hd__buf_6 _08873_ (.A(net18),
    .X(_04514_));
 sky130_fd_sc_hd__clkbuf_4 _08874_ (.A(_04514_),
    .X(_04515_));
 sky130_fd_sc_hd__mux2_1 _08875_ (.A0(net1569),
    .A1(_04515_),
    .S(_04503_),
    .X(_04516_));
 sky130_fd_sc_hd__clkbuf_1 _08876_ (.A(_04516_),
    .X(_01797_));
 sky130_fd_sc_hd__clkbuf_8 _08877_ (.A(net19),
    .X(_04517_));
 sky130_fd_sc_hd__clkbuf_4 _08878_ (.A(_04517_),
    .X(_04518_));
 sky130_fd_sc_hd__mux2_1 _08879_ (.A0(net433),
    .A1(_04518_),
    .S(_04503_),
    .X(_04519_));
 sky130_fd_sc_hd__clkbuf_1 _08880_ (.A(_04519_),
    .X(_01798_));
 sky130_fd_sc_hd__buf_6 _08881_ (.A(net20),
    .X(_04520_));
 sky130_fd_sc_hd__clkbuf_4 _08882_ (.A(_04520_),
    .X(_04521_));
 sky130_fd_sc_hd__mux2_1 _08883_ (.A0(net2022),
    .A1(_04521_),
    .S(_04503_),
    .X(_04522_));
 sky130_fd_sc_hd__clkbuf_1 _08884_ (.A(_04522_),
    .X(_01799_));
 sky130_fd_sc_hd__buf_6 _08885_ (.A(net21),
    .X(_04523_));
 sky130_fd_sc_hd__clkbuf_4 _08886_ (.A(_04523_),
    .X(_04524_));
 sky130_fd_sc_hd__mux2_1 _08887_ (.A0(net1110),
    .A1(_04524_),
    .S(_04503_),
    .X(_04525_));
 sky130_fd_sc_hd__clkbuf_1 _08888_ (.A(_04525_),
    .X(_01800_));
 sky130_fd_sc_hd__buf_6 _08889_ (.A(net22),
    .X(_04526_));
 sky130_fd_sc_hd__clkbuf_4 _08890_ (.A(_04526_),
    .X(_04527_));
 sky130_fd_sc_hd__mux2_1 _08891_ (.A0(net1780),
    .A1(_04527_),
    .S(_04503_),
    .X(_04528_));
 sky130_fd_sc_hd__clkbuf_1 _08892_ (.A(_04528_),
    .X(_01801_));
 sky130_fd_sc_hd__buf_6 _08893_ (.A(net23),
    .X(_04529_));
 sky130_fd_sc_hd__buf_4 _08894_ (.A(_04529_),
    .X(_04530_));
 sky130_fd_sc_hd__mux2_1 _08895_ (.A0(net441),
    .A1(_04530_),
    .S(_04503_),
    .X(_04531_));
 sky130_fd_sc_hd__clkbuf_1 _08896_ (.A(_04531_),
    .X(_01802_));
 sky130_fd_sc_hd__buf_8 _08897_ (.A(net9),
    .X(_04532_));
 sky130_fd_sc_hd__buf_4 _08898_ (.A(_04532_),
    .X(_04533_));
 sky130_fd_sc_hd__mux2_1 _08899_ (.A0(net74),
    .A1(_04533_),
    .S(_04502_),
    .X(_04534_));
 sky130_fd_sc_hd__clkbuf_1 _08900_ (.A(_04534_),
    .X(_01803_));
 sky130_fd_sc_hd__buf_6 _08901_ (.A(net10),
    .X(_04535_));
 sky130_fd_sc_hd__buf_4 _08902_ (.A(_04535_),
    .X(_04536_));
 sky130_fd_sc_hd__mux2_1 _08903_ (.A0(net882),
    .A1(_04536_),
    .S(_04502_),
    .X(_04537_));
 sky130_fd_sc_hd__clkbuf_1 _08904_ (.A(_04537_),
    .X(_01804_));
 sky130_fd_sc_hd__buf_6 _08905_ (.A(net11),
    .X(_04538_));
 sky130_fd_sc_hd__buf_4 _08906_ (.A(_04538_),
    .X(_04539_));
 sky130_fd_sc_hd__mux2_1 _08907_ (.A0(net485),
    .A1(_04539_),
    .S(_04502_),
    .X(_04540_));
 sky130_fd_sc_hd__clkbuf_1 _08908_ (.A(_04540_),
    .X(_01805_));
 sky130_fd_sc_hd__clkbuf_8 _08909_ (.A(net12),
    .X(_04541_));
 sky130_fd_sc_hd__clkbuf_4 _08910_ (.A(_04541_),
    .X(_04542_));
 sky130_fd_sc_hd__mux2_1 _08911_ (.A0(net490),
    .A1(_04542_),
    .S(_04502_),
    .X(_04543_));
 sky130_fd_sc_hd__clkbuf_1 _08912_ (.A(_04543_),
    .X(_01806_));
 sky130_fd_sc_hd__buf_6 _08913_ (.A(net13),
    .X(_04544_));
 sky130_fd_sc_hd__buf_4 _08914_ (.A(_04544_),
    .X(_04545_));
 sky130_fd_sc_hd__mux2_1 _08915_ (.A0(net651),
    .A1(_04545_),
    .S(_04502_),
    .X(_04546_));
 sky130_fd_sc_hd__clkbuf_1 _08916_ (.A(_04546_),
    .X(_01807_));
 sky130_fd_sc_hd__buf_6 _08917_ (.A(net14),
    .X(_04547_));
 sky130_fd_sc_hd__buf_4 _08918_ (.A(_04547_),
    .X(_04548_));
 sky130_fd_sc_hd__mux2_1 _08919_ (.A0(net705),
    .A1(_04548_),
    .S(_04502_),
    .X(_04549_));
 sky130_fd_sc_hd__clkbuf_1 _08920_ (.A(_04549_),
    .X(_01808_));
 sky130_fd_sc_hd__nor2_4 _08921_ (.A(_04072_),
    .B(_04368_),
    .Y(_04550_));
 sky130_fd_sc_hd__buf_4 _08922_ (.A(_04550_),
    .X(_04551_));
 sky130_fd_sc_hd__mux2_1 _08923_ (.A0(net989),
    .A1(_04499_),
    .S(_04551_),
    .X(_04552_));
 sky130_fd_sc_hd__clkbuf_1 _08924_ (.A(_04552_),
    .X(_01809_));
 sky130_fd_sc_hd__mux2_1 _08925_ (.A0(net956),
    .A1(_04506_),
    .S(_04551_),
    .X(_04553_));
 sky130_fd_sc_hd__clkbuf_1 _08926_ (.A(_04553_),
    .X(_01810_));
 sky130_fd_sc_hd__mux2_1 _08927_ (.A0(net787),
    .A1(_04509_),
    .S(_04551_),
    .X(_04554_));
 sky130_fd_sc_hd__clkbuf_1 _08928_ (.A(_04554_),
    .X(_01811_));
 sky130_fd_sc_hd__mux2_1 _08929_ (.A0(net932),
    .A1(_04512_),
    .S(_04551_),
    .X(_04555_));
 sky130_fd_sc_hd__clkbuf_1 _08930_ (.A(_04555_),
    .X(_01812_));
 sky130_fd_sc_hd__mux2_1 _08931_ (.A0(net1601),
    .A1(_04515_),
    .S(_04551_),
    .X(_04556_));
 sky130_fd_sc_hd__clkbuf_1 _08932_ (.A(_04556_),
    .X(_01813_));
 sky130_fd_sc_hd__mux2_1 _08933_ (.A0(net556),
    .A1(_04518_),
    .S(_04551_),
    .X(_04557_));
 sky130_fd_sc_hd__clkbuf_1 _08934_ (.A(_04557_),
    .X(_01814_));
 sky130_fd_sc_hd__mux2_1 _08935_ (.A0(net470),
    .A1(_04521_),
    .S(_04551_),
    .X(_04558_));
 sky130_fd_sc_hd__clkbuf_1 _08936_ (.A(_04558_),
    .X(_01815_));
 sky130_fd_sc_hd__mux2_1 _08937_ (.A0(net1623),
    .A1(_04524_),
    .S(_04551_),
    .X(_04559_));
 sky130_fd_sc_hd__clkbuf_1 _08938_ (.A(_04559_),
    .X(_01816_));
 sky130_fd_sc_hd__mux2_1 _08939_ (.A0(net1097),
    .A1(_04527_),
    .S(_04551_),
    .X(_04560_));
 sky130_fd_sc_hd__clkbuf_1 _08940_ (.A(_04560_),
    .X(_01817_));
 sky130_fd_sc_hd__mux2_1 _08941_ (.A0(net998),
    .A1(_04530_),
    .S(_04551_),
    .X(_04561_));
 sky130_fd_sc_hd__clkbuf_1 _08942_ (.A(_04561_),
    .X(_01818_));
 sky130_fd_sc_hd__mux2_1 _08943_ (.A0(net357),
    .A1(_04533_),
    .S(_04550_),
    .X(_04562_));
 sky130_fd_sc_hd__clkbuf_1 _08944_ (.A(_04562_),
    .X(_01819_));
 sky130_fd_sc_hd__mux2_1 _08945_ (.A0(net452),
    .A1(_04536_),
    .S(_04550_),
    .X(_04563_));
 sky130_fd_sc_hd__clkbuf_1 _08946_ (.A(_04563_),
    .X(_01820_));
 sky130_fd_sc_hd__mux2_1 _08947_ (.A0(net1573),
    .A1(_04539_),
    .S(_04550_),
    .X(_04564_));
 sky130_fd_sc_hd__clkbuf_1 _08948_ (.A(_04564_),
    .X(_01821_));
 sky130_fd_sc_hd__mux2_1 _08949_ (.A0(net377),
    .A1(_04542_),
    .S(_04550_),
    .X(_04565_));
 sky130_fd_sc_hd__clkbuf_1 _08950_ (.A(_04565_),
    .X(_01822_));
 sky130_fd_sc_hd__mux2_1 _08951_ (.A0(net901),
    .A1(_04545_),
    .S(_04550_),
    .X(_04566_));
 sky130_fd_sc_hd__clkbuf_1 _08952_ (.A(_04566_),
    .X(_01823_));
 sky130_fd_sc_hd__mux2_1 _08953_ (.A0(net1265),
    .A1(_04548_),
    .S(_04550_),
    .X(_04567_));
 sky130_fd_sc_hd__clkbuf_1 _08954_ (.A(_04567_),
    .X(_01824_));
 sky130_fd_sc_hd__or3_1 _08955_ (.A(_02656_),
    .B(_02492_),
    .C(_02497_),
    .X(_04568_));
 sky130_fd_sc_hd__buf_12 _08956_ (.A(_04568_),
    .X(_04569_));
 sky130_fd_sc_hd__nor2_8 _08957_ (.A(_04227_),
    .B(_04569_),
    .Y(_04570_));
 sky130_fd_sc_hd__buf_4 _08958_ (.A(_04570_),
    .X(_04571_));
 sky130_fd_sc_hd__mux2_1 _08959_ (.A0(net336),
    .A1(_04499_),
    .S(_04571_),
    .X(_04572_));
 sky130_fd_sc_hd__clkbuf_1 _08960_ (.A(_04572_),
    .X(_01825_));
 sky130_fd_sc_hd__mux2_1 _08961_ (.A0(net101),
    .A1(_04506_),
    .S(_04571_),
    .X(_04573_));
 sky130_fd_sc_hd__clkbuf_1 _08962_ (.A(_04573_),
    .X(_01826_));
 sky130_fd_sc_hd__mux2_1 _08963_ (.A0(net59),
    .A1(_04509_),
    .S(_04571_),
    .X(_04574_));
 sky130_fd_sc_hd__clkbuf_1 _08964_ (.A(_04574_),
    .X(_01827_));
 sky130_fd_sc_hd__mux2_1 _08965_ (.A0(net185),
    .A1(_04512_),
    .S(_04571_),
    .X(_04575_));
 sky130_fd_sc_hd__clkbuf_1 _08966_ (.A(_04575_),
    .X(_01828_));
 sky130_fd_sc_hd__mux2_1 _08967_ (.A0(net106),
    .A1(_04515_),
    .S(_04571_),
    .X(_04576_));
 sky130_fd_sc_hd__clkbuf_1 _08968_ (.A(_04576_),
    .X(_01829_));
 sky130_fd_sc_hd__mux2_1 _08969_ (.A0(net1719),
    .A1(_04518_),
    .S(_04571_),
    .X(_04577_));
 sky130_fd_sc_hd__clkbuf_1 _08970_ (.A(_04577_),
    .X(_01830_));
 sky130_fd_sc_hd__mux2_1 _08971_ (.A0(net135),
    .A1(_04521_),
    .S(_04571_),
    .X(_04578_));
 sky130_fd_sc_hd__clkbuf_1 _08972_ (.A(_04578_),
    .X(_01831_));
 sky130_fd_sc_hd__mux2_1 _08973_ (.A0(net126),
    .A1(_04524_),
    .S(_04571_),
    .X(_04579_));
 sky130_fd_sc_hd__clkbuf_1 _08974_ (.A(_04579_),
    .X(_01832_));
 sky130_fd_sc_hd__mux2_1 _08975_ (.A0(net70),
    .A1(_04527_),
    .S(_04571_),
    .X(_04580_));
 sky130_fd_sc_hd__clkbuf_1 _08976_ (.A(_04580_),
    .X(_01833_));
 sky130_fd_sc_hd__mux2_1 _08977_ (.A0(net465),
    .A1(_04530_),
    .S(_04571_),
    .X(_04581_));
 sky130_fd_sc_hd__clkbuf_1 _08978_ (.A(_04581_),
    .X(_01834_));
 sky130_fd_sc_hd__mux2_1 _08979_ (.A0(net112),
    .A1(_04533_),
    .S(_04570_),
    .X(_04582_));
 sky130_fd_sc_hd__clkbuf_1 _08980_ (.A(_04582_),
    .X(_01835_));
 sky130_fd_sc_hd__mux2_1 _08981_ (.A0(net129),
    .A1(_04536_),
    .S(_04570_),
    .X(_04583_));
 sky130_fd_sc_hd__clkbuf_1 _08982_ (.A(_04583_),
    .X(_01836_));
 sky130_fd_sc_hd__mux2_1 _08983_ (.A0(net161),
    .A1(_04539_),
    .S(_04570_),
    .X(_04584_));
 sky130_fd_sc_hd__clkbuf_1 _08984_ (.A(_04584_),
    .X(_01837_));
 sky130_fd_sc_hd__mux2_1 _08985_ (.A0(net395),
    .A1(_04542_),
    .S(_04570_),
    .X(_04585_));
 sky130_fd_sc_hd__clkbuf_1 _08986_ (.A(_04585_),
    .X(_01838_));
 sky130_fd_sc_hd__mux2_1 _08987_ (.A0(net205),
    .A1(_04545_),
    .S(_04570_),
    .X(_04586_));
 sky130_fd_sc_hd__clkbuf_1 _08988_ (.A(_04586_),
    .X(_01839_));
 sky130_fd_sc_hd__mux2_1 _08989_ (.A0(net191),
    .A1(_04548_),
    .S(_04570_),
    .X(_04587_));
 sky130_fd_sc_hd__clkbuf_1 _08990_ (.A(_04587_),
    .X(_01840_));
 sky130_fd_sc_hd__nor2_4 _08991_ (.A(_04184_),
    .B(_04227_),
    .Y(_04588_));
 sky130_fd_sc_hd__buf_4 _08992_ (.A(_04588_),
    .X(_04589_));
 sky130_fd_sc_hd__mux2_1 _08993_ (.A0(net1615),
    .A1(_04499_),
    .S(_04589_),
    .X(_04590_));
 sky130_fd_sc_hd__clkbuf_1 _08994_ (.A(_04590_),
    .X(_01841_));
 sky130_fd_sc_hd__mux2_1 _08995_ (.A0(net202),
    .A1(_04506_),
    .S(_04589_),
    .X(_04591_));
 sky130_fd_sc_hd__clkbuf_1 _08996_ (.A(_04591_),
    .X(_01842_));
 sky130_fd_sc_hd__mux2_1 _08997_ (.A0(net397),
    .A1(_04509_),
    .S(_04589_),
    .X(_04592_));
 sky130_fd_sc_hd__clkbuf_1 _08998_ (.A(_04592_),
    .X(_01843_));
 sky130_fd_sc_hd__mux2_1 _08999_ (.A0(net583),
    .A1(_04512_),
    .S(_04589_),
    .X(_04593_));
 sky130_fd_sc_hd__clkbuf_1 _09000_ (.A(_04593_),
    .X(_01844_));
 sky130_fd_sc_hd__mux2_1 _09001_ (.A0(net644),
    .A1(_04515_),
    .S(_04589_),
    .X(_04594_));
 sky130_fd_sc_hd__clkbuf_1 _09002_ (.A(_04594_),
    .X(_01845_));
 sky130_fd_sc_hd__mux2_1 _09003_ (.A0(net981),
    .A1(_04518_),
    .S(_04589_),
    .X(_04595_));
 sky130_fd_sc_hd__clkbuf_1 _09004_ (.A(_04595_),
    .X(_01846_));
 sky130_fd_sc_hd__mux2_1 _09005_ (.A0(net1667),
    .A1(_04521_),
    .S(_04589_),
    .X(_04596_));
 sky130_fd_sc_hd__clkbuf_1 _09006_ (.A(_04596_),
    .X(_01847_));
 sky130_fd_sc_hd__mux2_1 _09007_ (.A0(net1850),
    .A1(_04524_),
    .S(_04589_),
    .X(_04597_));
 sky130_fd_sc_hd__clkbuf_1 _09008_ (.A(_04597_),
    .X(_01848_));
 sky130_fd_sc_hd__mux2_1 _09009_ (.A0(net980),
    .A1(_04527_),
    .S(_04589_),
    .X(_04598_));
 sky130_fd_sc_hd__clkbuf_1 _09010_ (.A(_04598_),
    .X(_01849_));
 sky130_fd_sc_hd__mux2_1 _09011_ (.A0(net1225),
    .A1(_04530_),
    .S(_04589_),
    .X(_04599_));
 sky130_fd_sc_hd__clkbuf_1 _09012_ (.A(_04599_),
    .X(_01850_));
 sky130_fd_sc_hd__mux2_1 _09013_ (.A0(net1077),
    .A1(_04533_),
    .S(_04588_),
    .X(_04600_));
 sky130_fd_sc_hd__clkbuf_1 _09014_ (.A(_04600_),
    .X(_01851_));
 sky130_fd_sc_hd__mux2_1 _09015_ (.A0(net755),
    .A1(_04536_),
    .S(_04588_),
    .X(_04601_));
 sky130_fd_sc_hd__clkbuf_1 _09016_ (.A(_04601_),
    .X(_01852_));
 sky130_fd_sc_hd__mux2_1 _09017_ (.A0(net658),
    .A1(_04539_),
    .S(_04588_),
    .X(_04602_));
 sky130_fd_sc_hd__clkbuf_1 _09018_ (.A(_04602_),
    .X(_01853_));
 sky130_fd_sc_hd__mux2_1 _09019_ (.A0(net463),
    .A1(_04542_),
    .S(_04588_),
    .X(_04603_));
 sky130_fd_sc_hd__clkbuf_1 _09020_ (.A(_04603_),
    .X(_01854_));
 sky130_fd_sc_hd__mux2_1 _09021_ (.A0(net263),
    .A1(_04545_),
    .S(_04588_),
    .X(_04604_));
 sky130_fd_sc_hd__clkbuf_1 _09022_ (.A(_04604_),
    .X(_01855_));
 sky130_fd_sc_hd__mux2_1 _09023_ (.A0(net894),
    .A1(_04548_),
    .S(_04588_),
    .X(_04605_));
 sky130_fd_sc_hd__clkbuf_1 _09024_ (.A(_04605_),
    .X(_01856_));
 sky130_fd_sc_hd__or3b_1 _09025_ (.A(_02497_),
    .B(_02645_),
    .C_N(_02617_),
    .X(_04606_));
 sky130_fd_sc_hd__buf_12 _09026_ (.A(_04606_),
    .X(_04607_));
 sky130_fd_sc_hd__nor2_8 _09027_ (.A(_04227_),
    .B(_04607_),
    .Y(_04608_));
 sky130_fd_sc_hd__buf_4 _09028_ (.A(_04608_),
    .X(_04609_));
 sky130_fd_sc_hd__mux2_1 _09029_ (.A0(net1012),
    .A1(_04499_),
    .S(_04609_),
    .X(_04610_));
 sky130_fd_sc_hd__clkbuf_1 _09030_ (.A(_04610_),
    .X(_01857_));
 sky130_fd_sc_hd__mux2_1 _09031_ (.A0(net875),
    .A1(_04506_),
    .S(_04609_),
    .X(_04611_));
 sky130_fd_sc_hd__clkbuf_1 _09032_ (.A(_04611_),
    .X(_01858_));
 sky130_fd_sc_hd__mux2_1 _09033_ (.A0(net1470),
    .A1(_04509_),
    .S(_04609_),
    .X(_04612_));
 sky130_fd_sc_hd__clkbuf_1 _09034_ (.A(_04612_),
    .X(_01859_));
 sky130_fd_sc_hd__mux2_1 _09035_ (.A0(net1356),
    .A1(_04512_),
    .S(_04609_),
    .X(_04613_));
 sky130_fd_sc_hd__clkbuf_1 _09036_ (.A(_04613_),
    .X(_01860_));
 sky130_fd_sc_hd__mux2_1 _09037_ (.A0(net1292),
    .A1(_04515_),
    .S(_04609_),
    .X(_04614_));
 sky130_fd_sc_hd__clkbuf_1 _09038_ (.A(_04614_),
    .X(_01861_));
 sky130_fd_sc_hd__mux2_1 _09039_ (.A0(net1710),
    .A1(_04518_),
    .S(_04609_),
    .X(_04615_));
 sky130_fd_sc_hd__clkbuf_1 _09040_ (.A(_04615_),
    .X(_01862_));
 sky130_fd_sc_hd__mux2_1 _09041_ (.A0(net870),
    .A1(_04521_),
    .S(_04609_),
    .X(_04616_));
 sky130_fd_sc_hd__clkbuf_1 _09042_ (.A(_04616_),
    .X(_01863_));
 sky130_fd_sc_hd__mux2_1 _09043_ (.A0(net926),
    .A1(_04524_),
    .S(_04609_),
    .X(_04617_));
 sky130_fd_sc_hd__clkbuf_1 _09044_ (.A(_04617_),
    .X(_01864_));
 sky130_fd_sc_hd__mux2_1 _09045_ (.A0(net1387),
    .A1(_04527_),
    .S(_04609_),
    .X(_04618_));
 sky130_fd_sc_hd__clkbuf_1 _09046_ (.A(_04618_),
    .X(_01865_));
 sky130_fd_sc_hd__mux2_1 _09047_ (.A0(net1747),
    .A1(_04530_),
    .S(_04609_),
    .X(_04619_));
 sky130_fd_sc_hd__clkbuf_1 _09048_ (.A(_04619_),
    .X(_01866_));
 sky130_fd_sc_hd__mux2_1 _09049_ (.A0(net1283),
    .A1(_04533_),
    .S(_04608_),
    .X(_04620_));
 sky130_fd_sc_hd__clkbuf_1 _09050_ (.A(_04620_),
    .X(_01867_));
 sky130_fd_sc_hd__mux2_1 _09051_ (.A0(net1392),
    .A1(_04536_),
    .S(_04608_),
    .X(_04621_));
 sky130_fd_sc_hd__clkbuf_1 _09052_ (.A(_04621_),
    .X(_01868_));
 sky130_fd_sc_hd__mux2_1 _09053_ (.A0(net1127),
    .A1(_04539_),
    .S(_04608_),
    .X(_04622_));
 sky130_fd_sc_hd__clkbuf_1 _09054_ (.A(_04622_),
    .X(_01869_));
 sky130_fd_sc_hd__mux2_1 _09055_ (.A0(net1324),
    .A1(_04542_),
    .S(_04608_),
    .X(_04623_));
 sky130_fd_sc_hd__clkbuf_1 _09056_ (.A(_04623_),
    .X(_01870_));
 sky130_fd_sc_hd__mux2_1 _09057_ (.A0(net1558),
    .A1(_04545_),
    .S(_04608_),
    .X(_04624_));
 sky130_fd_sc_hd__clkbuf_1 _09058_ (.A(_04624_),
    .X(_01871_));
 sky130_fd_sc_hd__mux2_1 _09059_ (.A0(net1152),
    .A1(_04548_),
    .S(_04608_),
    .X(_04625_));
 sky130_fd_sc_hd__clkbuf_1 _09060_ (.A(_04625_),
    .X(_01872_));
 sky130_fd_sc_hd__or3_1 _09061_ (.A(_02702_),
    .B(_03092_),
    .C(_04226_),
    .X(_04626_));
 sky130_fd_sc_hd__buf_4 _09062_ (.A(_04626_),
    .X(_04627_));
 sky130_fd_sc_hd__buf_4 _09063_ (.A(_04627_),
    .X(_04628_));
 sky130_fd_sc_hd__mux2_1 _09064_ (.A0(_04406_),
    .A1(net1958),
    .S(_04628_),
    .X(_04629_));
 sky130_fd_sc_hd__clkbuf_1 _09065_ (.A(_04629_),
    .X(_01873_));
 sky130_fd_sc_hd__mux2_1 _09066_ (.A0(_04412_),
    .A1(net1273),
    .S(_04628_),
    .X(_04630_));
 sky130_fd_sc_hd__clkbuf_1 _09067_ (.A(_04630_),
    .X(_01874_));
 sky130_fd_sc_hd__mux2_1 _09068_ (.A0(_04414_),
    .A1(net1697),
    .S(_04628_),
    .X(_04631_));
 sky130_fd_sc_hd__clkbuf_1 _09069_ (.A(_04631_),
    .X(_01875_));
 sky130_fd_sc_hd__mux2_1 _09070_ (.A0(_04416_),
    .A1(net1946),
    .S(_04628_),
    .X(_04632_));
 sky130_fd_sc_hd__clkbuf_1 _09071_ (.A(_04632_),
    .X(_01876_));
 sky130_fd_sc_hd__mux2_1 _09072_ (.A0(_04418_),
    .A1(net1483),
    .S(_04628_),
    .X(_04633_));
 sky130_fd_sc_hd__clkbuf_1 _09073_ (.A(_04633_),
    .X(_01877_));
 sky130_fd_sc_hd__mux2_1 _09074_ (.A0(_04420_),
    .A1(net1647),
    .S(_04628_),
    .X(_04634_));
 sky130_fd_sc_hd__clkbuf_1 _09075_ (.A(_04634_),
    .X(_01878_));
 sky130_fd_sc_hd__mux2_1 _09076_ (.A0(_04422_),
    .A1(net1693),
    .S(_04628_),
    .X(_04635_));
 sky130_fd_sc_hd__clkbuf_1 _09077_ (.A(_04635_),
    .X(_01879_));
 sky130_fd_sc_hd__mux2_1 _09078_ (.A0(_04424_),
    .A1(net1096),
    .S(_04628_),
    .X(_04636_));
 sky130_fd_sc_hd__clkbuf_1 _09079_ (.A(_04636_),
    .X(_01880_));
 sky130_fd_sc_hd__mux2_1 _09080_ (.A0(_04426_),
    .A1(net2005),
    .S(_04628_),
    .X(_04637_));
 sky130_fd_sc_hd__clkbuf_1 _09081_ (.A(_04637_),
    .X(_01881_));
 sky130_fd_sc_hd__mux2_1 _09082_ (.A0(_04428_),
    .A1(net1926),
    .S(_04628_),
    .X(_04638_));
 sky130_fd_sc_hd__clkbuf_1 _09083_ (.A(_04638_),
    .X(_01882_));
 sky130_fd_sc_hd__mux2_1 _09084_ (.A0(_04430_),
    .A1(net1576),
    .S(_04627_),
    .X(_04639_));
 sky130_fd_sc_hd__clkbuf_1 _09085_ (.A(_04639_),
    .X(_01883_));
 sky130_fd_sc_hd__mux2_1 _09086_ (.A0(_04432_),
    .A1(net1578),
    .S(_04627_),
    .X(_04640_));
 sky130_fd_sc_hd__clkbuf_1 _09087_ (.A(_04640_),
    .X(_01884_));
 sky130_fd_sc_hd__mux2_1 _09088_ (.A0(_04434_),
    .A1(net1731),
    .S(_04627_),
    .X(_04641_));
 sky130_fd_sc_hd__clkbuf_1 _09089_ (.A(_04641_),
    .X(_01885_));
 sky130_fd_sc_hd__mux2_1 _09090_ (.A0(_04436_),
    .A1(net1833),
    .S(_04627_),
    .X(_04642_));
 sky130_fd_sc_hd__clkbuf_1 _09091_ (.A(_04642_),
    .X(_01886_));
 sky130_fd_sc_hd__mux2_1 _09092_ (.A0(_04438_),
    .A1(net1685),
    .S(_04627_),
    .X(_04643_));
 sky130_fd_sc_hd__clkbuf_1 _09093_ (.A(_04643_),
    .X(_01887_));
 sky130_fd_sc_hd__mux2_1 _09094_ (.A0(_04440_),
    .A1(net1582),
    .S(_04627_),
    .X(_04644_));
 sky130_fd_sc_hd__clkbuf_1 _09095_ (.A(_04644_),
    .X(_01888_));
 sky130_fd_sc_hd__or3_1 _09096_ (.A(_02656_),
    .B(_02492_),
    .C(_02505_),
    .X(_04645_));
 sky130_fd_sc_hd__buf_12 _09097_ (.A(_04645_),
    .X(_04646_));
 sky130_fd_sc_hd__nor2_8 _09098_ (.A(_04227_),
    .B(_04646_),
    .Y(_04647_));
 sky130_fd_sc_hd__buf_6 _09099_ (.A(_04647_),
    .X(_04648_));
 sky130_fd_sc_hd__mux2_1 _09100_ (.A0(net1481),
    .A1(_04499_),
    .S(_04648_),
    .X(_04649_));
 sky130_fd_sc_hd__clkbuf_1 _09101_ (.A(_04649_),
    .X(_01889_));
 sky130_fd_sc_hd__mux2_1 _09102_ (.A0(net492),
    .A1(_04506_),
    .S(_04648_),
    .X(_04650_));
 sky130_fd_sc_hd__clkbuf_1 _09103_ (.A(_04650_),
    .X(_01890_));
 sky130_fd_sc_hd__mux2_1 _09104_ (.A0(net1525),
    .A1(_04509_),
    .S(_04648_),
    .X(_04651_));
 sky130_fd_sc_hd__clkbuf_1 _09105_ (.A(_04651_),
    .X(_01891_));
 sky130_fd_sc_hd__mux2_1 _09106_ (.A0(net785),
    .A1(_04512_),
    .S(_04648_),
    .X(_04652_));
 sky130_fd_sc_hd__clkbuf_1 _09107_ (.A(_04652_),
    .X(_01892_));
 sky130_fd_sc_hd__mux2_1 _09108_ (.A0(net1055),
    .A1(_04515_),
    .S(_04648_),
    .X(_04653_));
 sky130_fd_sc_hd__clkbuf_1 _09109_ (.A(_04653_),
    .X(_01893_));
 sky130_fd_sc_hd__mux2_1 _09110_ (.A0(net676),
    .A1(_04518_),
    .S(_04648_),
    .X(_04654_));
 sky130_fd_sc_hd__clkbuf_1 _09111_ (.A(_04654_),
    .X(_01894_));
 sky130_fd_sc_hd__mux2_1 _09112_ (.A0(net1596),
    .A1(_04521_),
    .S(_04648_),
    .X(_04655_));
 sky130_fd_sc_hd__clkbuf_1 _09113_ (.A(_04655_),
    .X(_01895_));
 sky130_fd_sc_hd__mux2_1 _09114_ (.A0(net1109),
    .A1(_04524_),
    .S(_04648_),
    .X(_04656_));
 sky130_fd_sc_hd__clkbuf_1 _09115_ (.A(_04656_),
    .X(_01896_));
 sky130_fd_sc_hd__mux2_1 _09116_ (.A0(net1113),
    .A1(_04527_),
    .S(_04648_),
    .X(_04657_));
 sky130_fd_sc_hd__clkbuf_1 _09117_ (.A(_04657_),
    .X(_01897_));
 sky130_fd_sc_hd__mux2_1 _09118_ (.A0(net1272),
    .A1(_04530_),
    .S(_04648_),
    .X(_04658_));
 sky130_fd_sc_hd__clkbuf_1 _09119_ (.A(_04658_),
    .X(_01898_));
 sky130_fd_sc_hd__mux2_1 _09120_ (.A0(net1655),
    .A1(_04533_),
    .S(_04647_),
    .X(_04659_));
 sky130_fd_sc_hd__clkbuf_1 _09121_ (.A(_04659_),
    .X(_01899_));
 sky130_fd_sc_hd__mux2_1 _09122_ (.A0(net1782),
    .A1(_04536_),
    .S(_04647_),
    .X(_04660_));
 sky130_fd_sc_hd__clkbuf_1 _09123_ (.A(_04660_),
    .X(_01900_));
 sky130_fd_sc_hd__mux2_1 _09124_ (.A0(net1957),
    .A1(_04539_),
    .S(_04647_),
    .X(_04661_));
 sky130_fd_sc_hd__clkbuf_1 _09125_ (.A(_04661_),
    .X(_01901_));
 sky130_fd_sc_hd__mux2_1 _09126_ (.A0(net219),
    .A1(_04542_),
    .S(_04647_),
    .X(_04662_));
 sky130_fd_sc_hd__clkbuf_1 _09127_ (.A(_04662_),
    .X(_01902_));
 sky130_fd_sc_hd__mux2_1 _09128_ (.A0(net1805),
    .A1(_04545_),
    .S(_04647_),
    .X(_04663_));
 sky130_fd_sc_hd__clkbuf_1 _09129_ (.A(_04663_),
    .X(_01903_));
 sky130_fd_sc_hd__mux2_1 _09130_ (.A0(net1130),
    .A1(_04548_),
    .S(_04647_),
    .X(_04664_));
 sky130_fd_sc_hd__clkbuf_1 _09131_ (.A(_04664_),
    .X(_01904_));
 sky130_fd_sc_hd__nor2_8 _09132_ (.A(_04127_),
    .B(_04227_),
    .Y(_04665_));
 sky130_fd_sc_hd__buf_6 _09133_ (.A(_04665_),
    .X(_04666_));
 sky130_fd_sc_hd__mux2_1 _09134_ (.A0(net1100),
    .A1(_04499_),
    .S(_04666_),
    .X(_04667_));
 sky130_fd_sc_hd__clkbuf_1 _09135_ (.A(_04667_),
    .X(_01905_));
 sky130_fd_sc_hd__mux2_1 _09136_ (.A0(net879),
    .A1(_04506_),
    .S(_04666_),
    .X(_04668_));
 sky130_fd_sc_hd__clkbuf_1 _09137_ (.A(_04668_),
    .X(_01906_));
 sky130_fd_sc_hd__mux2_1 _09138_ (.A0(net933),
    .A1(_04509_),
    .S(_04666_),
    .X(_04669_));
 sky130_fd_sc_hd__clkbuf_1 _09139_ (.A(_04669_),
    .X(_01907_));
 sky130_fd_sc_hd__mux2_1 _09140_ (.A0(net794),
    .A1(_04512_),
    .S(_04666_),
    .X(_04670_));
 sky130_fd_sc_hd__clkbuf_1 _09141_ (.A(_04670_),
    .X(_01908_));
 sky130_fd_sc_hd__mux2_1 _09142_ (.A0(net273),
    .A1(_04515_),
    .S(_04666_),
    .X(_04671_));
 sky130_fd_sc_hd__clkbuf_1 _09143_ (.A(_04671_),
    .X(_01909_));
 sky130_fd_sc_hd__mux2_1 _09144_ (.A0(net1347),
    .A1(_04518_),
    .S(_04666_),
    .X(_04672_));
 sky130_fd_sc_hd__clkbuf_1 _09145_ (.A(_04672_),
    .X(_01910_));
 sky130_fd_sc_hd__mux2_1 _09146_ (.A0(net1497),
    .A1(_04521_),
    .S(_04666_),
    .X(_04673_));
 sky130_fd_sc_hd__clkbuf_1 _09147_ (.A(_04673_),
    .X(_01911_));
 sky130_fd_sc_hd__mux2_1 _09148_ (.A0(net753),
    .A1(_04524_),
    .S(_04666_),
    .X(_04674_));
 sky130_fd_sc_hd__clkbuf_1 _09149_ (.A(_04674_),
    .X(_01912_));
 sky130_fd_sc_hd__mux2_1 _09150_ (.A0(net1422),
    .A1(_04527_),
    .S(_04666_),
    .X(_04675_));
 sky130_fd_sc_hd__clkbuf_1 _09151_ (.A(_04675_),
    .X(_01913_));
 sky130_fd_sc_hd__mux2_1 _09152_ (.A0(net1043),
    .A1(_04530_),
    .S(_04666_),
    .X(_04676_));
 sky130_fd_sc_hd__clkbuf_1 _09153_ (.A(_04676_),
    .X(_01914_));
 sky130_fd_sc_hd__mux2_1 _09154_ (.A0(net1847),
    .A1(_04533_),
    .S(_04665_),
    .X(_04677_));
 sky130_fd_sc_hd__clkbuf_1 _09155_ (.A(_04677_),
    .X(_01915_));
 sky130_fd_sc_hd__mux2_1 _09156_ (.A0(net1336),
    .A1(_04536_),
    .S(_04665_),
    .X(_04678_));
 sky130_fd_sc_hd__clkbuf_1 _09157_ (.A(_04678_),
    .X(_01916_));
 sky130_fd_sc_hd__mux2_1 _09158_ (.A0(net1744),
    .A1(_04539_),
    .S(_04665_),
    .X(_04679_));
 sky130_fd_sc_hd__clkbuf_1 _09159_ (.A(_04679_),
    .X(_01917_));
 sky130_fd_sc_hd__mux2_1 _09160_ (.A0(net1472),
    .A1(_04542_),
    .S(_04665_),
    .X(_04680_));
 sky130_fd_sc_hd__clkbuf_1 _09161_ (.A(_04680_),
    .X(_01918_));
 sky130_fd_sc_hd__mux2_1 _09162_ (.A0(net1762),
    .A1(_04545_),
    .S(_04665_),
    .X(_04681_));
 sky130_fd_sc_hd__clkbuf_1 _09163_ (.A(_04681_),
    .X(_01919_));
 sky130_fd_sc_hd__mux2_1 _09164_ (.A0(net1777),
    .A1(_04548_),
    .S(_04665_),
    .X(_04682_));
 sky130_fd_sc_hd__clkbuf_1 _09165_ (.A(_04682_),
    .X(_01920_));
 sky130_fd_sc_hd__or3b_1 _09166_ (.A(_02505_),
    .B(_02645_),
    .C_N(_02617_),
    .X(_04683_));
 sky130_fd_sc_hd__buf_12 _09167_ (.A(_04683_),
    .X(_04684_));
 sky130_fd_sc_hd__nor2_8 _09168_ (.A(_04227_),
    .B(_04684_),
    .Y(_04685_));
 sky130_fd_sc_hd__buf_6 _09169_ (.A(_04685_),
    .X(_04686_));
 sky130_fd_sc_hd__mux2_1 _09170_ (.A0(net802),
    .A1(_04499_),
    .S(_04686_),
    .X(_04687_));
 sky130_fd_sc_hd__clkbuf_1 _09171_ (.A(_04687_),
    .X(_01921_));
 sky130_fd_sc_hd__mux2_1 _09172_ (.A0(net213),
    .A1(_04506_),
    .S(_04686_),
    .X(_04688_));
 sky130_fd_sc_hd__clkbuf_1 _09173_ (.A(_04688_),
    .X(_01922_));
 sky130_fd_sc_hd__mux2_1 _09174_ (.A0(net1625),
    .A1(_04509_),
    .S(_04686_),
    .X(_04689_));
 sky130_fd_sc_hd__clkbuf_1 _09175_ (.A(_04689_),
    .X(_01923_));
 sky130_fd_sc_hd__mux2_1 _09176_ (.A0(net663),
    .A1(_04512_),
    .S(_04686_),
    .X(_04690_));
 sky130_fd_sc_hd__clkbuf_1 _09177_ (.A(_04690_),
    .X(_01924_));
 sky130_fd_sc_hd__mux2_1 _09178_ (.A0(net1177),
    .A1(_04515_),
    .S(_04686_),
    .X(_04691_));
 sky130_fd_sc_hd__clkbuf_1 _09179_ (.A(_04691_),
    .X(_01925_));
 sky130_fd_sc_hd__mux2_1 _09180_ (.A0(net370),
    .A1(_04518_),
    .S(_04686_),
    .X(_04692_));
 sky130_fd_sc_hd__clkbuf_1 _09181_ (.A(_04692_),
    .X(_01926_));
 sky130_fd_sc_hd__mux2_1 _09182_ (.A0(net943),
    .A1(_04521_),
    .S(_04686_),
    .X(_04693_));
 sky130_fd_sc_hd__clkbuf_1 _09183_ (.A(_04693_),
    .X(_01927_));
 sky130_fd_sc_hd__mux2_1 _09184_ (.A0(net846),
    .A1(_04524_),
    .S(_04686_),
    .X(_04694_));
 sky130_fd_sc_hd__clkbuf_1 _09185_ (.A(_04694_),
    .X(_01928_));
 sky130_fd_sc_hd__mux2_1 _09186_ (.A0(net1773),
    .A1(_04527_),
    .S(_04686_),
    .X(_04695_));
 sky130_fd_sc_hd__clkbuf_1 _09187_ (.A(_04695_),
    .X(_01929_));
 sky130_fd_sc_hd__mux2_1 _09188_ (.A0(net647),
    .A1(_04530_),
    .S(_04686_),
    .X(_04696_));
 sky130_fd_sc_hd__clkbuf_1 _09189_ (.A(_04696_),
    .X(_01930_));
 sky130_fd_sc_hd__mux2_1 _09190_ (.A0(net916),
    .A1(_04533_),
    .S(_04685_),
    .X(_04697_));
 sky130_fd_sc_hd__clkbuf_1 _09191_ (.A(_04697_),
    .X(_01931_));
 sky130_fd_sc_hd__mux2_1 _09192_ (.A0(net1598),
    .A1(_04536_),
    .S(_04685_),
    .X(_04698_));
 sky130_fd_sc_hd__clkbuf_1 _09193_ (.A(_04698_),
    .X(_01932_));
 sky130_fd_sc_hd__mux2_1 _09194_ (.A0(net1778),
    .A1(_04539_),
    .S(_04685_),
    .X(_04699_));
 sky130_fd_sc_hd__clkbuf_1 _09195_ (.A(_04699_),
    .X(_01933_));
 sky130_fd_sc_hd__mux2_1 _09196_ (.A0(net388),
    .A1(_04542_),
    .S(_04685_),
    .X(_04700_));
 sky130_fd_sc_hd__clkbuf_1 _09197_ (.A(_04700_),
    .X(_01934_));
 sky130_fd_sc_hd__mux2_1 _09198_ (.A0(net1252),
    .A1(_04545_),
    .S(_04685_),
    .X(_04701_));
 sky130_fd_sc_hd__clkbuf_1 _09199_ (.A(_04701_),
    .X(_01935_));
 sky130_fd_sc_hd__mux2_1 _09200_ (.A0(net1315),
    .A1(_04548_),
    .S(_04685_),
    .X(_04702_));
 sky130_fd_sc_hd__clkbuf_1 _09201_ (.A(_04702_),
    .X(_01936_));
 sky130_fd_sc_hd__or3_1 _09202_ (.A(_02707_),
    .B(_03092_),
    .C(_04226_),
    .X(_04703_));
 sky130_fd_sc_hd__buf_4 _09203_ (.A(_04703_),
    .X(_04704_));
 sky130_fd_sc_hd__buf_6 _09204_ (.A(_04704_),
    .X(_04705_));
 sky130_fd_sc_hd__mux2_1 _09205_ (.A0(_04406_),
    .A1(net1861),
    .S(_04705_),
    .X(_04706_));
 sky130_fd_sc_hd__clkbuf_1 _09206_ (.A(_04706_),
    .X(_01937_));
 sky130_fd_sc_hd__mux2_1 _09207_ (.A0(_04412_),
    .A1(net1852),
    .S(_04705_),
    .X(_04707_));
 sky130_fd_sc_hd__clkbuf_1 _09208_ (.A(_04707_),
    .X(_01938_));
 sky130_fd_sc_hd__mux2_1 _09209_ (.A0(_04414_),
    .A1(net1126),
    .S(_04705_),
    .X(_04708_));
 sky130_fd_sc_hd__clkbuf_1 _09210_ (.A(_04708_),
    .X(_01939_));
 sky130_fd_sc_hd__mux2_1 _09211_ (.A0(_04416_),
    .A1(net1793),
    .S(_04705_),
    .X(_04709_));
 sky130_fd_sc_hd__clkbuf_1 _09212_ (.A(_04709_),
    .X(_01940_));
 sky130_fd_sc_hd__mux2_1 _09213_ (.A0(_04418_),
    .A1(net1572),
    .S(_04705_),
    .X(_04710_));
 sky130_fd_sc_hd__clkbuf_1 _09214_ (.A(_04710_),
    .X(_01941_));
 sky130_fd_sc_hd__mux2_1 _09215_ (.A0(_04420_),
    .A1(net1823),
    .S(_04705_),
    .X(_04711_));
 sky130_fd_sc_hd__clkbuf_1 _09216_ (.A(_04711_),
    .X(_01942_));
 sky130_fd_sc_hd__mux2_1 _09217_ (.A0(_04422_),
    .A1(net1493),
    .S(_04705_),
    .X(_04712_));
 sky130_fd_sc_hd__clkbuf_1 _09218_ (.A(_04712_),
    .X(_01943_));
 sky130_fd_sc_hd__mux2_1 _09219_ (.A0(_04424_),
    .A1(net1864),
    .S(_04705_),
    .X(_04713_));
 sky130_fd_sc_hd__clkbuf_1 _09220_ (.A(_04713_),
    .X(_01944_));
 sky130_fd_sc_hd__mux2_1 _09221_ (.A0(_04426_),
    .A1(net1769),
    .S(_04705_),
    .X(_04714_));
 sky130_fd_sc_hd__clkbuf_1 _09222_ (.A(_04714_),
    .X(_01945_));
 sky130_fd_sc_hd__mux2_1 _09223_ (.A0(_04428_),
    .A1(net1459),
    .S(_04705_),
    .X(_04715_));
 sky130_fd_sc_hd__clkbuf_1 _09224_ (.A(_04715_),
    .X(_01946_));
 sky130_fd_sc_hd__mux2_1 _09225_ (.A0(_04430_),
    .A1(net1634),
    .S(_04704_),
    .X(_04716_));
 sky130_fd_sc_hd__clkbuf_1 _09226_ (.A(_04716_),
    .X(_01947_));
 sky130_fd_sc_hd__mux2_1 _09227_ (.A0(_04432_),
    .A1(net1689),
    .S(_04704_),
    .X(_04717_));
 sky130_fd_sc_hd__clkbuf_1 _09228_ (.A(_04717_),
    .X(_01948_));
 sky130_fd_sc_hd__mux2_1 _09229_ (.A0(_04434_),
    .A1(net1688),
    .S(_04704_),
    .X(_04718_));
 sky130_fd_sc_hd__clkbuf_1 _09230_ (.A(_04718_),
    .X(_01949_));
 sky130_fd_sc_hd__mux2_1 _09231_ (.A0(_04436_),
    .A1(net822),
    .S(_04704_),
    .X(_04719_));
 sky130_fd_sc_hd__clkbuf_1 _09232_ (.A(_04719_),
    .X(_01950_));
 sky130_fd_sc_hd__mux2_1 _09233_ (.A0(_04438_),
    .A1(net1661),
    .S(_04704_),
    .X(_04720_));
 sky130_fd_sc_hd__clkbuf_1 _09234_ (.A(_04720_),
    .X(_01951_));
 sky130_fd_sc_hd__mux2_1 _09235_ (.A0(_04440_),
    .A1(net1712),
    .S(_04704_),
    .X(_04721_));
 sky130_fd_sc_hd__clkbuf_1 _09236_ (.A(_04721_),
    .X(_01952_));
 sky130_fd_sc_hd__nor2_8 _09237_ (.A(_04226_),
    .B(_04365_),
    .Y(_04722_));
 sky130_fd_sc_hd__buf_4 _09238_ (.A(_04722_),
    .X(_04723_));
 sky130_fd_sc_hd__mux2_1 _09239_ (.A0(net137),
    .A1(_04499_),
    .S(_04723_),
    .X(_04724_));
 sky130_fd_sc_hd__clkbuf_1 _09240_ (.A(_04724_),
    .X(_01953_));
 sky130_fd_sc_hd__mux2_1 _09241_ (.A0(net595),
    .A1(_04506_),
    .S(_04723_),
    .X(_04725_));
 sky130_fd_sc_hd__clkbuf_1 _09242_ (.A(_04725_),
    .X(_01954_));
 sky130_fd_sc_hd__mux2_1 _09243_ (.A0(net206),
    .A1(_04509_),
    .S(_04723_),
    .X(_04726_));
 sky130_fd_sc_hd__clkbuf_1 _09244_ (.A(_04726_),
    .X(_01955_));
 sky130_fd_sc_hd__mux2_1 _09245_ (.A0(net864),
    .A1(_04512_),
    .S(_04723_),
    .X(_04727_));
 sky130_fd_sc_hd__clkbuf_1 _09246_ (.A(_04727_),
    .X(_01956_));
 sky130_fd_sc_hd__mux2_1 _09247_ (.A0(net960),
    .A1(_04515_),
    .S(_04723_),
    .X(_04728_));
 sky130_fd_sc_hd__clkbuf_1 _09248_ (.A(_04728_),
    .X(_01957_));
 sky130_fd_sc_hd__mux2_1 _09249_ (.A0(net1306),
    .A1(_04518_),
    .S(_04723_),
    .X(_04729_));
 sky130_fd_sc_hd__clkbuf_1 _09250_ (.A(_04729_),
    .X(_01958_));
 sky130_fd_sc_hd__mux2_1 _09251_ (.A0(net1916),
    .A1(_04521_),
    .S(_04723_),
    .X(_04730_));
 sky130_fd_sc_hd__clkbuf_1 _09252_ (.A(_04730_),
    .X(_01959_));
 sky130_fd_sc_hd__mux2_1 _09253_ (.A0(net277),
    .A1(_04524_),
    .S(_04723_),
    .X(_04731_));
 sky130_fd_sc_hd__clkbuf_1 _09254_ (.A(_04731_),
    .X(_01960_));
 sky130_fd_sc_hd__mux2_1 _09255_ (.A0(net1436),
    .A1(_04527_),
    .S(_04723_),
    .X(_04732_));
 sky130_fd_sc_hd__clkbuf_1 _09256_ (.A(_04732_),
    .X(_01961_));
 sky130_fd_sc_hd__mux2_1 _09257_ (.A0(net300),
    .A1(_04530_),
    .S(_04723_),
    .X(_04733_));
 sky130_fd_sc_hd__clkbuf_1 _09258_ (.A(_04733_),
    .X(_01962_));
 sky130_fd_sc_hd__mux2_1 _09259_ (.A0(net117),
    .A1(_04533_),
    .S(_04722_),
    .X(_04734_));
 sky130_fd_sc_hd__clkbuf_1 _09260_ (.A(_04734_),
    .X(_01963_));
 sky130_fd_sc_hd__mux2_1 _09261_ (.A0(net58),
    .A1(_04536_),
    .S(_04722_),
    .X(_04735_));
 sky130_fd_sc_hd__clkbuf_1 _09262_ (.A(_04735_),
    .X(_01964_));
 sky130_fd_sc_hd__mux2_1 _09263_ (.A0(net146),
    .A1(_04539_),
    .S(_04722_),
    .X(_04736_));
 sky130_fd_sc_hd__clkbuf_1 _09264_ (.A(_04736_),
    .X(_01965_));
 sky130_fd_sc_hd__mux2_1 _09265_ (.A0(net276),
    .A1(_04542_),
    .S(_04722_),
    .X(_04737_));
 sky130_fd_sc_hd__clkbuf_1 _09266_ (.A(_04737_),
    .X(_01966_));
 sky130_fd_sc_hd__mux2_1 _09267_ (.A0(net335),
    .A1(_04545_),
    .S(_04722_),
    .X(_04738_));
 sky130_fd_sc_hd__clkbuf_1 _09268_ (.A(_04738_),
    .X(_01967_));
 sky130_fd_sc_hd__mux2_1 _09269_ (.A0(net88),
    .A1(_04548_),
    .S(_04722_),
    .X(_04739_));
 sky130_fd_sc_hd__clkbuf_1 _09270_ (.A(_04739_),
    .X(_01968_));
 sky130_fd_sc_hd__nor2_4 _09271_ (.A(_04368_),
    .B(_04501_),
    .Y(_04740_));
 sky130_fd_sc_hd__buf_4 _09272_ (.A(_04740_),
    .X(_04741_));
 sky130_fd_sc_hd__mux2_1 _09273_ (.A0(net444),
    .A1(_04499_),
    .S(_04741_),
    .X(_04742_));
 sky130_fd_sc_hd__clkbuf_1 _09274_ (.A(_04742_),
    .X(_01969_));
 sky130_fd_sc_hd__mux2_1 _09275_ (.A0(net387),
    .A1(_04506_),
    .S(_04741_),
    .X(_04743_));
 sky130_fd_sc_hd__clkbuf_1 _09276_ (.A(_04743_),
    .X(_01970_));
 sky130_fd_sc_hd__mux2_1 _09277_ (.A0(net695),
    .A1(_04509_),
    .S(_04741_),
    .X(_04744_));
 sky130_fd_sc_hd__clkbuf_1 _09278_ (.A(_04744_),
    .X(_01971_));
 sky130_fd_sc_hd__mux2_1 _09279_ (.A0(net1844),
    .A1(_04512_),
    .S(_04741_),
    .X(_04745_));
 sky130_fd_sc_hd__clkbuf_1 _09280_ (.A(_04745_),
    .X(_01972_));
 sky130_fd_sc_hd__mux2_1 _09281_ (.A0(net220),
    .A1(_04515_),
    .S(_04741_),
    .X(_04746_));
 sky130_fd_sc_hd__clkbuf_1 _09282_ (.A(_04746_),
    .X(_01973_));
 sky130_fd_sc_hd__mux2_1 _09283_ (.A0(net507),
    .A1(_04518_),
    .S(_04741_),
    .X(_04747_));
 sky130_fd_sc_hd__clkbuf_1 _09284_ (.A(_04747_),
    .X(_01974_));
 sky130_fd_sc_hd__mux2_1 _09285_ (.A0(net443),
    .A1(_04521_),
    .S(_04741_),
    .X(_04748_));
 sky130_fd_sc_hd__clkbuf_1 _09286_ (.A(_04748_),
    .X(_01975_));
 sky130_fd_sc_hd__mux2_1 _09287_ (.A0(net826),
    .A1(_04524_),
    .S(_04741_),
    .X(_04749_));
 sky130_fd_sc_hd__clkbuf_1 _09288_ (.A(_04749_),
    .X(_01976_));
 sky130_fd_sc_hd__mux2_1 _09289_ (.A0(net552),
    .A1(_04527_),
    .S(_04741_),
    .X(_04750_));
 sky130_fd_sc_hd__clkbuf_1 _09290_ (.A(_04750_),
    .X(_01977_));
 sky130_fd_sc_hd__mux2_1 _09291_ (.A0(net491),
    .A1(_04530_),
    .S(_04741_),
    .X(_04751_));
 sky130_fd_sc_hd__clkbuf_1 _09292_ (.A(_04751_),
    .X(_01978_));
 sky130_fd_sc_hd__mux2_1 _09293_ (.A0(net1466),
    .A1(_04533_),
    .S(_04740_),
    .X(_04752_));
 sky130_fd_sc_hd__clkbuf_1 _09294_ (.A(_04752_),
    .X(_01979_));
 sky130_fd_sc_hd__mux2_1 _09295_ (.A0(net612),
    .A1(_04536_),
    .S(_04740_),
    .X(_04753_));
 sky130_fd_sc_hd__clkbuf_1 _09296_ (.A(_04753_),
    .X(_01980_));
 sky130_fd_sc_hd__mux2_1 _09297_ (.A0(net1162),
    .A1(_04539_),
    .S(_04740_),
    .X(_04754_));
 sky130_fd_sc_hd__clkbuf_1 _09298_ (.A(_04754_),
    .X(_01981_));
 sky130_fd_sc_hd__mux2_1 _09299_ (.A0(net256),
    .A1(_04542_),
    .S(_04740_),
    .X(_04755_));
 sky130_fd_sc_hd__clkbuf_1 _09300_ (.A(_04755_),
    .X(_01982_));
 sky130_fd_sc_hd__mux2_1 _09301_ (.A0(net1567),
    .A1(_04545_),
    .S(_04740_),
    .X(_04756_));
 sky130_fd_sc_hd__clkbuf_1 _09302_ (.A(_04756_),
    .X(_01983_));
 sky130_fd_sc_hd__mux2_1 _09303_ (.A0(net889),
    .A1(_04548_),
    .S(_04740_),
    .X(_04757_));
 sky130_fd_sc_hd__clkbuf_1 _09304_ (.A(_04757_),
    .X(_01984_));
 sky130_fd_sc_hd__nand2b_4 _09305_ (.A_N(_04226_),
    .B(_04408_),
    .Y(_04758_));
 sky130_fd_sc_hd__buf_4 _09306_ (.A(_04758_),
    .X(_04759_));
 sky130_fd_sc_hd__mux2_1 _09307_ (.A0(_04406_),
    .A1(net1509),
    .S(_04759_),
    .X(_04760_));
 sky130_fd_sc_hd__clkbuf_1 _09308_ (.A(_04760_),
    .X(_01985_));
 sky130_fd_sc_hd__mux2_1 _09309_ (.A0(_04412_),
    .A1(net1873),
    .S(_04759_),
    .X(_04761_));
 sky130_fd_sc_hd__clkbuf_1 _09310_ (.A(_04761_),
    .X(_01986_));
 sky130_fd_sc_hd__mux2_1 _09311_ (.A0(_04414_),
    .A1(net1763),
    .S(_04759_),
    .X(_04762_));
 sky130_fd_sc_hd__clkbuf_1 _09312_ (.A(_04762_),
    .X(_01987_));
 sky130_fd_sc_hd__mux2_1 _09313_ (.A0(_04416_),
    .A1(net1545),
    .S(_04759_),
    .X(_04763_));
 sky130_fd_sc_hd__clkbuf_1 _09314_ (.A(_04763_),
    .X(_01988_));
 sky130_fd_sc_hd__mux2_1 _09315_ (.A0(_04418_),
    .A1(net1530),
    .S(_04759_),
    .X(_04764_));
 sky130_fd_sc_hd__clkbuf_1 _09316_ (.A(_04764_),
    .X(_01989_));
 sky130_fd_sc_hd__mux2_1 _09317_ (.A0(_04420_),
    .A1(net1994),
    .S(_04759_),
    .X(_04765_));
 sky130_fd_sc_hd__clkbuf_1 _09318_ (.A(_04765_),
    .X(_01990_));
 sky130_fd_sc_hd__mux2_1 _09319_ (.A0(_04422_),
    .A1(net1832),
    .S(_04759_),
    .X(_04766_));
 sky130_fd_sc_hd__clkbuf_1 _09320_ (.A(_04766_),
    .X(_01991_));
 sky130_fd_sc_hd__mux2_1 _09321_ (.A0(_04424_),
    .A1(net1927),
    .S(_04759_),
    .X(_04767_));
 sky130_fd_sc_hd__clkbuf_1 _09322_ (.A(_04767_),
    .X(_01992_));
 sky130_fd_sc_hd__mux2_1 _09323_ (.A0(_04426_),
    .A1(net1934),
    .S(_04759_),
    .X(_04768_));
 sky130_fd_sc_hd__clkbuf_1 _09324_ (.A(_04768_),
    .X(_01993_));
 sky130_fd_sc_hd__mux2_1 _09325_ (.A0(_04428_),
    .A1(net1417),
    .S(_04759_),
    .X(_04769_));
 sky130_fd_sc_hd__clkbuf_1 _09326_ (.A(_04769_),
    .X(_01994_));
 sky130_fd_sc_hd__mux2_1 _09327_ (.A0(_04430_),
    .A1(net1666),
    .S(_04758_),
    .X(_04770_));
 sky130_fd_sc_hd__clkbuf_1 _09328_ (.A(_04770_),
    .X(_01995_));
 sky130_fd_sc_hd__mux2_1 _09329_ (.A0(_04432_),
    .A1(net1675),
    .S(_04758_),
    .X(_04771_));
 sky130_fd_sc_hd__clkbuf_1 _09330_ (.A(_04771_),
    .X(_01996_));
 sky130_fd_sc_hd__mux2_1 _09331_ (.A0(_04434_),
    .A1(net1888),
    .S(_04758_),
    .X(_04772_));
 sky130_fd_sc_hd__clkbuf_1 _09332_ (.A(_04772_),
    .X(_01997_));
 sky130_fd_sc_hd__mux2_1 _09333_ (.A0(_04436_),
    .A1(net1905),
    .S(_04758_),
    .X(_04773_));
 sky130_fd_sc_hd__clkbuf_1 _09334_ (.A(_04773_),
    .X(_01998_));
 sky130_fd_sc_hd__mux2_1 _09335_ (.A0(_04438_),
    .A1(net1229),
    .S(_04758_),
    .X(_04774_));
 sky130_fd_sc_hd__clkbuf_1 _09336_ (.A(_04774_),
    .X(_01999_));
 sky130_fd_sc_hd__mux2_1 _09337_ (.A0(_04440_),
    .A1(net1658),
    .S(_04758_),
    .X(_04775_));
 sky130_fd_sc_hd__clkbuf_1 _09338_ (.A(_04775_),
    .X(_02000_));
 sky130_fd_sc_hd__or3_1 _09339_ (.A(_04059_),
    .B(_03092_),
    .C(_04226_),
    .X(_04776_));
 sky130_fd_sc_hd__buf_4 _09340_ (.A(_04776_),
    .X(_04777_));
 sky130_fd_sc_hd__buf_4 _09341_ (.A(_04777_),
    .X(_04778_));
 sky130_fd_sc_hd__mux2_1 _09342_ (.A0(_04406_),
    .A1(net1668),
    .S(_04778_),
    .X(_04779_));
 sky130_fd_sc_hd__clkbuf_1 _09343_ (.A(_04779_),
    .X(_02001_));
 sky130_fd_sc_hd__mux2_1 _09344_ (.A0(_04412_),
    .A1(net1449),
    .S(_04778_),
    .X(_04780_));
 sky130_fd_sc_hd__clkbuf_1 _09345_ (.A(_04780_),
    .X(_02002_));
 sky130_fd_sc_hd__mux2_1 _09346_ (.A0(_04414_),
    .A1(net1329),
    .S(_04778_),
    .X(_04781_));
 sky130_fd_sc_hd__clkbuf_1 _09347_ (.A(_04781_),
    .X(_02003_));
 sky130_fd_sc_hd__mux2_1 _09348_ (.A0(_04416_),
    .A1(net1711),
    .S(_04778_),
    .X(_04782_));
 sky130_fd_sc_hd__clkbuf_1 _09349_ (.A(_04782_),
    .X(_02004_));
 sky130_fd_sc_hd__mux2_1 _09350_ (.A0(_04418_),
    .A1(net1851),
    .S(_04778_),
    .X(_04783_));
 sky130_fd_sc_hd__clkbuf_1 _09351_ (.A(_04783_),
    .X(_02005_));
 sky130_fd_sc_hd__mux2_1 _09352_ (.A0(_04420_),
    .A1(net1860),
    .S(_04778_),
    .X(_04784_));
 sky130_fd_sc_hd__clkbuf_1 _09353_ (.A(_04784_),
    .X(_02006_));
 sky130_fd_sc_hd__mux2_1 _09354_ (.A0(_04422_),
    .A1(net1240),
    .S(_04778_),
    .X(_04785_));
 sky130_fd_sc_hd__clkbuf_1 _09355_ (.A(_04785_),
    .X(_02007_));
 sky130_fd_sc_hd__mux2_1 _09356_ (.A0(_04424_),
    .A1(net1384),
    .S(_04778_),
    .X(_04786_));
 sky130_fd_sc_hd__clkbuf_1 _09357_ (.A(_04786_),
    .X(_02008_));
 sky130_fd_sc_hd__mux2_1 _09358_ (.A0(_04426_),
    .A1(net1700),
    .S(_04778_),
    .X(_04787_));
 sky130_fd_sc_hd__clkbuf_1 _09359_ (.A(_04787_),
    .X(_02009_));
 sky130_fd_sc_hd__mux2_1 _09360_ (.A0(_04428_),
    .A1(net1775),
    .S(_04778_),
    .X(_04788_));
 sky130_fd_sc_hd__clkbuf_1 _09361_ (.A(_04788_),
    .X(_02010_));
 sky130_fd_sc_hd__mux2_1 _09362_ (.A0(_04430_),
    .A1(net1742),
    .S(_04777_),
    .X(_04789_));
 sky130_fd_sc_hd__clkbuf_1 _09363_ (.A(_04789_),
    .X(_02011_));
 sky130_fd_sc_hd__mux2_1 _09364_ (.A0(_04432_),
    .A1(net1388),
    .S(_04777_),
    .X(_04790_));
 sky130_fd_sc_hd__clkbuf_1 _09365_ (.A(_04790_),
    .X(_02012_));
 sky130_fd_sc_hd__mux2_1 _09366_ (.A0(_04434_),
    .A1(net814),
    .S(_04777_),
    .X(_04791_));
 sky130_fd_sc_hd__clkbuf_1 _09367_ (.A(_04791_),
    .X(_02013_));
 sky130_fd_sc_hd__mux2_1 _09368_ (.A0(_04436_),
    .A1(net1890),
    .S(_04777_),
    .X(_04792_));
 sky130_fd_sc_hd__clkbuf_1 _09369_ (.A(_04792_),
    .X(_02014_));
 sky130_fd_sc_hd__mux2_1 _09370_ (.A0(_04438_),
    .A1(net1727),
    .S(_04777_),
    .X(_04793_));
 sky130_fd_sc_hd__clkbuf_1 _09371_ (.A(_04793_),
    .X(_02015_));
 sky130_fd_sc_hd__mux2_1 _09372_ (.A0(_04440_),
    .A1(net1893),
    .S(_04777_),
    .X(_04794_));
 sky130_fd_sc_hd__clkbuf_1 _09373_ (.A(_04794_),
    .X(_02016_));
 sky130_fd_sc_hd__clkbuf_4 _09374_ (.A(_04498_),
    .X(_04795_));
 sky130_fd_sc_hd__buf_8 _09375_ (.A(_04246_),
    .X(_04796_));
 sky130_fd_sc_hd__nor2_4 _09376_ (.A(_04796_),
    .B(_04461_),
    .Y(_04797_));
 sky130_fd_sc_hd__buf_6 _09377_ (.A(_04797_),
    .X(_04798_));
 sky130_fd_sc_hd__mux2_1 _09378_ (.A0(net827),
    .A1(_04795_),
    .S(_04798_),
    .X(_04799_));
 sky130_fd_sc_hd__clkbuf_1 _09379_ (.A(_04799_),
    .X(_02017_));
 sky130_fd_sc_hd__clkbuf_4 _09380_ (.A(_04505_),
    .X(_04800_));
 sky130_fd_sc_hd__mux2_1 _09381_ (.A0(net250),
    .A1(_04800_),
    .S(_04798_),
    .X(_04801_));
 sky130_fd_sc_hd__clkbuf_1 _09382_ (.A(_04801_),
    .X(_02018_));
 sky130_fd_sc_hd__clkbuf_4 _09383_ (.A(_04508_),
    .X(_04802_));
 sky130_fd_sc_hd__mux2_1 _09384_ (.A0(net233),
    .A1(_04802_),
    .S(_04798_),
    .X(_04803_));
 sky130_fd_sc_hd__clkbuf_1 _09385_ (.A(_04803_),
    .X(_02019_));
 sky130_fd_sc_hd__buf_4 _09386_ (.A(_04511_),
    .X(_04804_));
 sky130_fd_sc_hd__mux2_1 _09387_ (.A0(net376),
    .A1(_04804_),
    .S(_04798_),
    .X(_04805_));
 sky130_fd_sc_hd__clkbuf_1 _09388_ (.A(_04805_),
    .X(_02020_));
 sky130_fd_sc_hd__buf_4 _09389_ (.A(_04514_),
    .X(_04806_));
 sky130_fd_sc_hd__mux2_1 _09390_ (.A0(net1040),
    .A1(_04806_),
    .S(_04798_),
    .X(_04807_));
 sky130_fd_sc_hd__clkbuf_1 _09391_ (.A(_04807_),
    .X(_02021_));
 sky130_fd_sc_hd__clkbuf_4 _09392_ (.A(_04517_),
    .X(_04808_));
 sky130_fd_sc_hd__mux2_1 _09393_ (.A0(net208),
    .A1(_04808_),
    .S(_04798_),
    .X(_04809_));
 sky130_fd_sc_hd__clkbuf_1 _09394_ (.A(_04809_),
    .X(_02022_));
 sky130_fd_sc_hd__buf_4 _09395_ (.A(_04520_),
    .X(_04810_));
 sky130_fd_sc_hd__mux2_1 _09396_ (.A0(net1081),
    .A1(_04810_),
    .S(_04798_),
    .X(_04811_));
 sky130_fd_sc_hd__clkbuf_1 _09397_ (.A(_04811_),
    .X(_02023_));
 sky130_fd_sc_hd__buf_4 _09398_ (.A(_04523_),
    .X(_04812_));
 sky130_fd_sc_hd__mux2_1 _09399_ (.A0(net1054),
    .A1(_04812_),
    .S(_04798_),
    .X(_04813_));
 sky130_fd_sc_hd__clkbuf_1 _09400_ (.A(_04813_),
    .X(_02024_));
 sky130_fd_sc_hd__buf_4 _09401_ (.A(_04526_),
    .X(_04814_));
 sky130_fd_sc_hd__mux2_1 _09402_ (.A0(net1382),
    .A1(_04814_),
    .S(_04798_),
    .X(_04815_));
 sky130_fd_sc_hd__clkbuf_1 _09403_ (.A(_04815_),
    .X(_02025_));
 sky130_fd_sc_hd__buf_4 _09404_ (.A(_04529_),
    .X(_04816_));
 sky130_fd_sc_hd__mux2_1 _09405_ (.A0(net531),
    .A1(_04816_),
    .S(_04798_),
    .X(_04817_));
 sky130_fd_sc_hd__clkbuf_1 _09406_ (.A(_04817_),
    .X(_02026_));
 sky130_fd_sc_hd__clkbuf_4 _09407_ (.A(_04532_),
    .X(_04818_));
 sky130_fd_sc_hd__mux2_1 _09408_ (.A0(net498),
    .A1(_04818_),
    .S(_04797_),
    .X(_04819_));
 sky130_fd_sc_hd__clkbuf_1 _09409_ (.A(_04819_),
    .X(_02027_));
 sky130_fd_sc_hd__buf_4 _09410_ (.A(_04535_),
    .X(_04820_));
 sky130_fd_sc_hd__mux2_1 _09411_ (.A0(net1257),
    .A1(_04820_),
    .S(_04797_),
    .X(_04821_));
 sky130_fd_sc_hd__clkbuf_1 _09412_ (.A(_04821_),
    .X(_02028_));
 sky130_fd_sc_hd__buf_4 _09413_ (.A(_04538_),
    .X(_04822_));
 sky130_fd_sc_hd__mux2_1 _09414_ (.A0(net432),
    .A1(_04822_),
    .S(_04797_),
    .X(_04823_));
 sky130_fd_sc_hd__clkbuf_1 _09415_ (.A(_04823_),
    .X(_02029_));
 sky130_fd_sc_hd__clkbuf_4 _09416_ (.A(_04541_),
    .X(_04824_));
 sky130_fd_sc_hd__mux2_1 _09417_ (.A0(net599),
    .A1(_04824_),
    .S(_04797_),
    .X(_04825_));
 sky130_fd_sc_hd__clkbuf_1 _09418_ (.A(_04825_),
    .X(_02030_));
 sky130_fd_sc_hd__clkbuf_4 _09419_ (.A(_04544_),
    .X(_04826_));
 sky130_fd_sc_hd__mux2_1 _09420_ (.A0(net749),
    .A1(_04826_),
    .S(_04797_),
    .X(_04827_));
 sky130_fd_sc_hd__clkbuf_1 _09421_ (.A(_04827_),
    .X(_02031_));
 sky130_fd_sc_hd__clkbuf_4 _09422_ (.A(_04547_),
    .X(_04828_));
 sky130_fd_sc_hd__mux2_1 _09423_ (.A0(net435),
    .A1(_04828_),
    .S(_04797_),
    .X(_04829_));
 sky130_fd_sc_hd__clkbuf_1 _09424_ (.A(_04829_),
    .X(_02032_));
 sky130_fd_sc_hd__nor2_4 _09425_ (.A(_04072_),
    .B(_04796_),
    .Y(_04830_));
 sky130_fd_sc_hd__buf_6 _09426_ (.A(_04830_),
    .X(_04831_));
 sky130_fd_sc_hd__mux2_1 _09427_ (.A0(net302),
    .A1(_04795_),
    .S(_04831_),
    .X(_04832_));
 sky130_fd_sc_hd__clkbuf_1 _09428_ (.A(_04832_),
    .X(_02033_));
 sky130_fd_sc_hd__mux2_1 _09429_ (.A0(net207),
    .A1(_04800_),
    .S(_04831_),
    .X(_04833_));
 sky130_fd_sc_hd__clkbuf_1 _09430_ (.A(_04833_),
    .X(_02034_));
 sky130_fd_sc_hd__mux2_1 _09431_ (.A0(net579),
    .A1(_04802_),
    .S(_04831_),
    .X(_04834_));
 sky130_fd_sc_hd__clkbuf_1 _09432_ (.A(_04834_),
    .X(_02035_));
 sky130_fd_sc_hd__mux2_1 _09433_ (.A0(net801),
    .A1(_04804_),
    .S(_04831_),
    .X(_04835_));
 sky130_fd_sc_hd__clkbuf_1 _09434_ (.A(_04835_),
    .X(_02036_));
 sky130_fd_sc_hd__mux2_1 _09435_ (.A0(net681),
    .A1(_04806_),
    .S(_04831_),
    .X(_04836_));
 sky130_fd_sc_hd__clkbuf_1 _09436_ (.A(_04836_),
    .X(_02037_));
 sky130_fd_sc_hd__mux2_1 _09437_ (.A0(net416),
    .A1(_04808_),
    .S(_04831_),
    .X(_04837_));
 sky130_fd_sc_hd__clkbuf_1 _09438_ (.A(_04837_),
    .X(_02038_));
 sky130_fd_sc_hd__mux2_1 _09439_ (.A0(net453),
    .A1(_04810_),
    .S(_04831_),
    .X(_04838_));
 sky130_fd_sc_hd__clkbuf_1 _09440_ (.A(_04838_),
    .X(_02039_));
 sky130_fd_sc_hd__mux2_1 _09441_ (.A0(net1717),
    .A1(_04812_),
    .S(_04831_),
    .X(_04839_));
 sky130_fd_sc_hd__clkbuf_1 _09442_ (.A(_04839_),
    .X(_02040_));
 sky130_fd_sc_hd__mux2_1 _09443_ (.A0(net484),
    .A1(_04814_),
    .S(_04831_),
    .X(_04840_));
 sky130_fd_sc_hd__clkbuf_1 _09444_ (.A(_04840_),
    .X(_02041_));
 sky130_fd_sc_hd__mux2_1 _09445_ (.A0(net193),
    .A1(_04816_),
    .S(_04831_),
    .X(_04841_));
 sky130_fd_sc_hd__clkbuf_1 _09446_ (.A(_04841_),
    .X(_02042_));
 sky130_fd_sc_hd__mux2_1 _09447_ (.A0(net390),
    .A1(_04818_),
    .S(_04830_),
    .X(_04842_));
 sky130_fd_sc_hd__clkbuf_1 _09448_ (.A(_04842_),
    .X(_02043_));
 sky130_fd_sc_hd__mux2_1 _09449_ (.A0(net223),
    .A1(_04820_),
    .S(_04830_),
    .X(_04843_));
 sky130_fd_sc_hd__clkbuf_1 _09450_ (.A(_04843_),
    .X(_02044_));
 sky130_fd_sc_hd__mux2_1 _09451_ (.A0(net113),
    .A1(_04822_),
    .S(_04830_),
    .X(_04844_));
 sky130_fd_sc_hd__clkbuf_1 _09452_ (.A(_04844_),
    .X(_02045_));
 sky130_fd_sc_hd__mux2_1 _09453_ (.A0(net721),
    .A1(_04824_),
    .S(_04830_),
    .X(_04845_));
 sky130_fd_sc_hd__clkbuf_1 _09454_ (.A(_04845_),
    .X(_02046_));
 sky130_fd_sc_hd__mux2_1 _09455_ (.A0(net53),
    .A1(_04826_),
    .S(_04830_),
    .X(_04846_));
 sky130_fd_sc_hd__clkbuf_1 _09456_ (.A(_04846_),
    .X(_02047_));
 sky130_fd_sc_hd__mux2_1 _09457_ (.A0(net1199),
    .A1(_04828_),
    .S(_04830_),
    .X(_04847_));
 sky130_fd_sc_hd__clkbuf_1 _09458_ (.A(_04847_),
    .X(_02048_));
 sky130_fd_sc_hd__nor2_4 _09459_ (.A(_04796_),
    .B(_04501_),
    .Y(_04848_));
 sky130_fd_sc_hd__buf_6 _09460_ (.A(_04848_),
    .X(_04849_));
 sky130_fd_sc_hd__mux2_1 _09461_ (.A0(net1300),
    .A1(_04795_),
    .S(_04849_),
    .X(_04850_));
 sky130_fd_sc_hd__clkbuf_1 _09462_ (.A(_04850_),
    .X(_02049_));
 sky130_fd_sc_hd__mux2_1 _09463_ (.A0(net562),
    .A1(_04800_),
    .S(_04849_),
    .X(_04851_));
 sky130_fd_sc_hd__clkbuf_1 _09464_ (.A(_04851_),
    .X(_02050_));
 sky130_fd_sc_hd__mux2_1 _09465_ (.A0(net1457),
    .A1(_04802_),
    .S(_04849_),
    .X(_04852_));
 sky130_fd_sc_hd__clkbuf_1 _09466_ (.A(_04852_),
    .X(_02051_));
 sky130_fd_sc_hd__mux2_1 _09467_ (.A0(net354),
    .A1(_04804_),
    .S(_04849_),
    .X(_04853_));
 sky130_fd_sc_hd__clkbuf_1 _09468_ (.A(_04853_),
    .X(_02052_));
 sky130_fd_sc_hd__mux2_1 _09469_ (.A0(net1085),
    .A1(_04806_),
    .S(_04849_),
    .X(_04854_));
 sky130_fd_sc_hd__clkbuf_1 _09470_ (.A(_04854_),
    .X(_02053_));
 sky130_fd_sc_hd__mux2_1 _09471_ (.A0(net685),
    .A1(_04808_),
    .S(_04849_),
    .X(_04855_));
 sky130_fd_sc_hd__clkbuf_1 _09472_ (.A(_04855_),
    .X(_02054_));
 sky130_fd_sc_hd__mux2_1 _09473_ (.A0(net1088),
    .A1(_04810_),
    .S(_04849_),
    .X(_04856_));
 sky130_fd_sc_hd__clkbuf_1 _09474_ (.A(_04856_),
    .X(_02055_));
 sky130_fd_sc_hd__mux2_1 _09475_ (.A0(net626),
    .A1(_04812_),
    .S(_04849_),
    .X(_04857_));
 sky130_fd_sc_hd__clkbuf_1 _09476_ (.A(_04857_),
    .X(_02056_));
 sky130_fd_sc_hd__mux2_1 _09477_ (.A0(net1279),
    .A1(_04814_),
    .S(_04849_),
    .X(_04858_));
 sky130_fd_sc_hd__clkbuf_1 _09478_ (.A(_04858_),
    .X(_02057_));
 sky130_fd_sc_hd__mux2_1 _09479_ (.A0(net493),
    .A1(_04816_),
    .S(_04849_),
    .X(_04859_));
 sky130_fd_sc_hd__clkbuf_1 _09480_ (.A(_04859_),
    .X(_02058_));
 sky130_fd_sc_hd__mux2_1 _09481_ (.A0(net805),
    .A1(_04818_),
    .S(_04848_),
    .X(_04860_));
 sky130_fd_sc_hd__clkbuf_1 _09482_ (.A(_04860_),
    .X(_02059_));
 sky130_fd_sc_hd__mux2_1 _09483_ (.A0(net971),
    .A1(_04820_),
    .S(_04848_),
    .X(_04861_));
 sky130_fd_sc_hd__clkbuf_1 _09484_ (.A(_04861_),
    .X(_02060_));
 sky130_fd_sc_hd__mux2_1 _09485_ (.A0(net1758),
    .A1(_04822_),
    .S(_04848_),
    .X(_04862_));
 sky130_fd_sc_hd__clkbuf_1 _09486_ (.A(_04862_),
    .X(_02061_));
 sky130_fd_sc_hd__mux2_1 _09487_ (.A0(net296),
    .A1(_04824_),
    .S(_04848_),
    .X(_04863_));
 sky130_fd_sc_hd__clkbuf_1 _09488_ (.A(_04863_),
    .X(_02062_));
 sky130_fd_sc_hd__mux2_1 _09489_ (.A0(net1093),
    .A1(_04826_),
    .S(_04848_),
    .X(_04864_));
 sky130_fd_sc_hd__clkbuf_1 _09490_ (.A(_04864_),
    .X(_02063_));
 sky130_fd_sc_hd__mux2_1 _09491_ (.A0(net1437),
    .A1(_04828_),
    .S(_04848_),
    .X(_04865_));
 sky130_fd_sc_hd__clkbuf_1 _09492_ (.A(_04865_),
    .X(_00016_));
 sky130_fd_sc_hd__nor2_4 _09493_ (.A(_04225_),
    .B(_04796_),
    .Y(_04866_));
 sky130_fd_sc_hd__buf_6 _09494_ (.A(_04866_),
    .X(_04867_));
 sky130_fd_sc_hd__mux2_1 _09495_ (.A0(net68),
    .A1(_04795_),
    .S(_04867_),
    .X(_04868_));
 sky130_fd_sc_hd__clkbuf_1 _09496_ (.A(_04868_),
    .X(_00017_));
 sky130_fd_sc_hd__mux2_1 _09497_ (.A0(net196),
    .A1(_04800_),
    .S(_04867_),
    .X(_04869_));
 sky130_fd_sc_hd__clkbuf_1 _09498_ (.A(_04869_),
    .X(_00018_));
 sky130_fd_sc_hd__mux2_1 _09499_ (.A0(net576),
    .A1(_04802_),
    .S(_04867_),
    .X(_04870_));
 sky130_fd_sc_hd__clkbuf_1 _09500_ (.A(_04870_),
    .X(_00019_));
 sky130_fd_sc_hd__mux2_1 _09501_ (.A0(net437),
    .A1(_04804_),
    .S(_04867_),
    .X(_04871_));
 sky130_fd_sc_hd__clkbuf_1 _09502_ (.A(_04871_),
    .X(_00020_));
 sky130_fd_sc_hd__mux2_1 _09503_ (.A0(net886),
    .A1(_04806_),
    .S(_04867_),
    .X(_04872_));
 sky130_fd_sc_hd__clkbuf_1 _09504_ (.A(_04872_),
    .X(_00021_));
 sky130_fd_sc_hd__mux2_1 _09505_ (.A0(net235),
    .A1(_04808_),
    .S(_04867_),
    .X(_04873_));
 sky130_fd_sc_hd__clkbuf_1 _09506_ (.A(_04873_),
    .X(_00022_));
 sky130_fd_sc_hd__mux2_1 _09507_ (.A0(net292),
    .A1(_04810_),
    .S(_04867_),
    .X(_04874_));
 sky130_fd_sc_hd__clkbuf_1 _09508_ (.A(_04874_),
    .X(_00023_));
 sky130_fd_sc_hd__mux2_1 _09509_ (.A0(net769),
    .A1(_04812_),
    .S(_04867_),
    .X(_04875_));
 sky130_fd_sc_hd__clkbuf_1 _09510_ (.A(_04875_),
    .X(_00024_));
 sky130_fd_sc_hd__mux2_1 _09511_ (.A0(net895),
    .A1(_04814_),
    .S(_04867_),
    .X(_04876_));
 sky130_fd_sc_hd__clkbuf_1 _09512_ (.A(_04876_),
    .X(_00025_));
 sky130_fd_sc_hd__mux2_1 _09513_ (.A0(net311),
    .A1(_04816_),
    .S(_04867_),
    .X(_04877_));
 sky130_fd_sc_hd__clkbuf_1 _09514_ (.A(_04877_),
    .X(_00026_));
 sky130_fd_sc_hd__mux2_1 _09515_ (.A0(net481),
    .A1(_04818_),
    .S(_04866_),
    .X(_04878_));
 sky130_fd_sc_hd__clkbuf_1 _09516_ (.A(_04878_),
    .X(_00027_));
 sky130_fd_sc_hd__mux2_1 _09517_ (.A0(net722),
    .A1(_04820_),
    .S(_04866_),
    .X(_04879_));
 sky130_fd_sc_hd__clkbuf_1 _09518_ (.A(_04879_),
    .X(_00028_));
 sky130_fd_sc_hd__mux2_1 _09519_ (.A0(net1756),
    .A1(_04822_),
    .S(_04866_),
    .X(_04880_));
 sky130_fd_sc_hd__clkbuf_1 _09520_ (.A(_04880_),
    .X(_00029_));
 sky130_fd_sc_hd__mux2_1 _09521_ (.A0(net63),
    .A1(_04824_),
    .S(_04866_),
    .X(_04881_));
 sky130_fd_sc_hd__clkbuf_1 _09522_ (.A(_04881_),
    .X(_00030_));
 sky130_fd_sc_hd__mux2_1 _09523_ (.A0(net123),
    .A1(_04826_),
    .S(_04866_),
    .X(_04882_));
 sky130_fd_sc_hd__clkbuf_1 _09524_ (.A(_04882_),
    .X(_00031_));
 sky130_fd_sc_hd__mux2_1 _09525_ (.A0(net167),
    .A1(_04828_),
    .S(_04866_),
    .X(_04883_));
 sky130_fd_sc_hd__clkbuf_1 _09526_ (.A(_04883_),
    .X(_00032_));
 sky130_fd_sc_hd__nor2_4 _09527_ (.A(_04796_),
    .B(_04569_),
    .Y(_04884_));
 sky130_fd_sc_hd__buf_6 _09528_ (.A(_04884_),
    .X(_04885_));
 sky130_fd_sc_hd__mux2_1 _09529_ (.A0(net657),
    .A1(_04795_),
    .S(_04885_),
    .X(_04886_));
 sky130_fd_sc_hd__clkbuf_1 _09530_ (.A(_04886_),
    .X(_00033_));
 sky130_fd_sc_hd__mux2_1 _09531_ (.A0(net999),
    .A1(_04800_),
    .S(_04885_),
    .X(_04887_));
 sky130_fd_sc_hd__clkbuf_1 _09532_ (.A(_04887_),
    .X(_00034_));
 sky130_fd_sc_hd__mux2_1 _09533_ (.A0(net361),
    .A1(_04802_),
    .S(_04885_),
    .X(_04888_));
 sky130_fd_sc_hd__clkbuf_1 _09534_ (.A(_04888_),
    .X(_00035_));
 sky130_fd_sc_hd__mux2_1 _09535_ (.A0(net472),
    .A1(_04804_),
    .S(_04885_),
    .X(_04889_));
 sky130_fd_sc_hd__clkbuf_1 _09536_ (.A(_04889_),
    .X(_00036_));
 sky130_fd_sc_hd__mux2_1 _09537_ (.A0(net1223),
    .A1(_04806_),
    .S(_04885_),
    .X(_04890_));
 sky130_fd_sc_hd__clkbuf_1 _09538_ (.A(_04890_),
    .X(_00037_));
 sky130_fd_sc_hd__mux2_1 _09539_ (.A0(net775),
    .A1(_04808_),
    .S(_04885_),
    .X(_04891_));
 sky130_fd_sc_hd__clkbuf_1 _09540_ (.A(_04891_),
    .X(_00038_));
 sky130_fd_sc_hd__mux2_1 _09541_ (.A0(net299),
    .A1(_04810_),
    .S(_04885_),
    .X(_04892_));
 sky130_fd_sc_hd__clkbuf_1 _09542_ (.A(_04892_),
    .X(_00039_));
 sky130_fd_sc_hd__mux2_1 _09543_ (.A0(net372),
    .A1(_04812_),
    .S(_04885_),
    .X(_04893_));
 sky130_fd_sc_hd__clkbuf_1 _09544_ (.A(_04893_),
    .X(_00040_));
 sky130_fd_sc_hd__mux2_1 _09545_ (.A0(net953),
    .A1(_04814_),
    .S(_04885_),
    .X(_04894_));
 sky130_fd_sc_hd__clkbuf_1 _09546_ (.A(_04894_),
    .X(_00041_));
 sky130_fd_sc_hd__mux2_1 _09547_ (.A0(net262),
    .A1(_04816_),
    .S(_04885_),
    .X(_04895_));
 sky130_fd_sc_hd__clkbuf_1 _09548_ (.A(_04895_),
    .X(_00042_));
 sky130_fd_sc_hd__mux2_1 _09549_ (.A0(net976),
    .A1(_04818_),
    .S(_04884_),
    .X(_04896_));
 sky130_fd_sc_hd__clkbuf_1 _09550_ (.A(_04896_),
    .X(_00043_));
 sky130_fd_sc_hd__mux2_1 _09551_ (.A0(net290),
    .A1(_04820_),
    .S(_04884_),
    .X(_04897_));
 sky130_fd_sc_hd__clkbuf_1 _09552_ (.A(_04897_),
    .X(_00044_));
 sky130_fd_sc_hd__mux2_1 _09553_ (.A0(net254),
    .A1(_04822_),
    .S(_04884_),
    .X(_04898_));
 sky130_fd_sc_hd__clkbuf_1 _09554_ (.A(_04898_),
    .X(_00045_));
 sky130_fd_sc_hd__mux2_1 _09555_ (.A0(net1107),
    .A1(_04824_),
    .S(_04884_),
    .X(_04899_));
 sky130_fd_sc_hd__clkbuf_1 _09556_ (.A(_04899_),
    .X(_00046_));
 sky130_fd_sc_hd__mux2_1 _09557_ (.A0(net1027),
    .A1(_04826_),
    .S(_04884_),
    .X(_04900_));
 sky130_fd_sc_hd__clkbuf_1 _09558_ (.A(_04900_),
    .X(_00047_));
 sky130_fd_sc_hd__mux2_1 _09559_ (.A0(net142),
    .A1(_04828_),
    .S(_04884_),
    .X(_04901_));
 sky130_fd_sc_hd__clkbuf_1 _09560_ (.A(_04901_),
    .X(_00048_));
 sky130_fd_sc_hd__nor2_4 _09561_ (.A(_04184_),
    .B(_04796_),
    .Y(_04902_));
 sky130_fd_sc_hd__buf_6 _09562_ (.A(_04902_),
    .X(_04903_));
 sky130_fd_sc_hd__mux2_1 _09563_ (.A0(net188),
    .A1(_04795_),
    .S(_04903_),
    .X(_04904_));
 sky130_fd_sc_hd__clkbuf_1 _09564_ (.A(_04904_),
    .X(_00049_));
 sky130_fd_sc_hd__mux2_1 _09565_ (.A0(net103),
    .A1(_04800_),
    .S(_04903_),
    .X(_04905_));
 sky130_fd_sc_hd__clkbuf_1 _09566_ (.A(_04905_),
    .X(_00050_));
 sky130_fd_sc_hd__mux2_1 _09567_ (.A0(net99),
    .A1(_04802_),
    .S(_04903_),
    .X(_04906_));
 sky130_fd_sc_hd__clkbuf_1 _09568_ (.A(_04906_),
    .X(_00051_));
 sky130_fd_sc_hd__mux2_1 _09569_ (.A0(net118),
    .A1(_04804_),
    .S(_04903_),
    .X(_04907_));
 sky130_fd_sc_hd__clkbuf_1 _09570_ (.A(_04907_),
    .X(_00052_));
 sky130_fd_sc_hd__mux2_1 _09571_ (.A0(net419),
    .A1(_04806_),
    .S(_04903_),
    .X(_04908_));
 sky130_fd_sc_hd__clkbuf_1 _09572_ (.A(_04908_),
    .X(_00053_));
 sky130_fd_sc_hd__mux2_1 _09573_ (.A0(net48),
    .A1(_04808_),
    .S(_04903_),
    .X(_04909_));
 sky130_fd_sc_hd__clkbuf_1 _09574_ (.A(_04909_),
    .X(_00054_));
 sky130_fd_sc_hd__mux2_1 _09575_ (.A0(net51),
    .A1(_04810_),
    .S(_04903_),
    .X(_04910_));
 sky130_fd_sc_hd__clkbuf_1 _09576_ (.A(_04910_),
    .X(_00055_));
 sky130_fd_sc_hd__mux2_1 _09577_ (.A0(net211),
    .A1(_04812_),
    .S(_04903_),
    .X(_04911_));
 sky130_fd_sc_hd__clkbuf_1 _09578_ (.A(_04911_),
    .X(_00056_));
 sky130_fd_sc_hd__mux2_1 _09579_ (.A0(net64),
    .A1(_04814_),
    .S(_04903_),
    .X(_04912_));
 sky130_fd_sc_hd__clkbuf_1 _09580_ (.A(_04912_),
    .X(_00057_));
 sky130_fd_sc_hd__mux2_1 _09581_ (.A0(net267),
    .A1(_04816_),
    .S(_04903_),
    .X(_04913_));
 sky130_fd_sc_hd__clkbuf_1 _09582_ (.A(_04913_),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _09583_ (.A0(net417),
    .A1(_04818_),
    .S(_04902_),
    .X(_04914_));
 sky130_fd_sc_hd__clkbuf_1 _09584_ (.A(_04914_),
    .X(_00059_));
 sky130_fd_sc_hd__mux2_1 _09585_ (.A0(net374),
    .A1(_04820_),
    .S(_04902_),
    .X(_04915_));
 sky130_fd_sc_hd__clkbuf_1 _09586_ (.A(_04915_),
    .X(_00060_));
 sky130_fd_sc_hd__mux2_1 _09587_ (.A0(net629),
    .A1(_04822_),
    .S(_04902_),
    .X(_04916_));
 sky130_fd_sc_hd__clkbuf_1 _09588_ (.A(_04916_),
    .X(_00061_));
 sky130_fd_sc_hd__mux2_1 _09589_ (.A0(net434),
    .A1(_04824_),
    .S(_04902_),
    .X(_04917_));
 sky130_fd_sc_hd__clkbuf_1 _09590_ (.A(_04917_),
    .X(_00062_));
 sky130_fd_sc_hd__mux2_1 _09591_ (.A0(net181),
    .A1(_04826_),
    .S(_04902_),
    .X(_04918_));
 sky130_fd_sc_hd__clkbuf_1 _09592_ (.A(_04918_),
    .X(_00063_));
 sky130_fd_sc_hd__mux2_1 _09593_ (.A0(net572),
    .A1(_04828_),
    .S(_04902_),
    .X(_04919_));
 sky130_fd_sc_hd__clkbuf_1 _09594_ (.A(_04919_),
    .X(_00064_));
 sky130_fd_sc_hd__nor2_4 _09595_ (.A(_04796_),
    .B(_04607_),
    .Y(_04920_));
 sky130_fd_sc_hd__buf_6 _09596_ (.A(_04920_),
    .X(_04921_));
 sky130_fd_sc_hd__mux2_1 _09597_ (.A0(net378),
    .A1(_04795_),
    .S(_04921_),
    .X(_04922_));
 sky130_fd_sc_hd__clkbuf_1 _09598_ (.A(_04922_),
    .X(_00065_));
 sky130_fd_sc_hd__mux2_1 _09599_ (.A0(net412),
    .A1(_04800_),
    .S(_04921_),
    .X(_04923_));
 sky130_fd_sc_hd__clkbuf_1 _09600_ (.A(_04923_),
    .X(_00066_));
 sky130_fd_sc_hd__mux2_1 _09601_ (.A0(net132),
    .A1(_04802_),
    .S(_04921_),
    .X(_04924_));
 sky130_fd_sc_hd__clkbuf_1 _09602_ (.A(_04924_),
    .X(_00067_));
 sky130_fd_sc_hd__mux2_1 _09603_ (.A0(net344),
    .A1(_04804_),
    .S(_04921_),
    .X(_04925_));
 sky130_fd_sc_hd__clkbuf_1 _09604_ (.A(_04925_),
    .X(_00068_));
 sky130_fd_sc_hd__mux2_1 _09605_ (.A0(net350),
    .A1(_04806_),
    .S(_04921_),
    .X(_04926_));
 sky130_fd_sc_hd__clkbuf_1 _09606_ (.A(_04926_),
    .X(_00069_));
 sky130_fd_sc_hd__mux2_1 _09607_ (.A0(net1045),
    .A1(_04808_),
    .S(_04921_),
    .X(_04927_));
 sky130_fd_sc_hd__clkbuf_1 _09608_ (.A(_04927_),
    .X(_00070_));
 sky130_fd_sc_hd__mux2_1 _09609_ (.A0(net428),
    .A1(_04810_),
    .S(_04921_),
    .X(_04928_));
 sky130_fd_sc_hd__clkbuf_1 _09610_ (.A(_04928_),
    .X(_00071_));
 sky130_fd_sc_hd__mux2_1 _09611_ (.A0(net639),
    .A1(_04812_),
    .S(_04921_),
    .X(_04929_));
 sky130_fd_sc_hd__clkbuf_1 _09612_ (.A(_04929_),
    .X(_00072_));
 sky130_fd_sc_hd__mux2_1 _09613_ (.A0(net985),
    .A1(_04814_),
    .S(_04921_),
    .X(_04930_));
 sky130_fd_sc_hd__clkbuf_1 _09614_ (.A(_04930_),
    .X(_00073_));
 sky130_fd_sc_hd__mux2_1 _09615_ (.A0(net283),
    .A1(_04816_),
    .S(_04921_),
    .X(_04931_));
 sky130_fd_sc_hd__clkbuf_1 _09616_ (.A(_04931_),
    .X(_00074_));
 sky130_fd_sc_hd__mux2_1 _09617_ (.A0(net1099),
    .A1(_04818_),
    .S(_04920_),
    .X(_04932_));
 sky130_fd_sc_hd__clkbuf_1 _09618_ (.A(_04932_),
    .X(_00075_));
 sky130_fd_sc_hd__mux2_1 _09619_ (.A0(net334),
    .A1(_04820_),
    .S(_04920_),
    .X(_04933_));
 sky130_fd_sc_hd__clkbuf_1 _09620_ (.A(_04933_),
    .X(_00076_));
 sky130_fd_sc_hd__mux2_1 _09621_ (.A0(net471),
    .A1(_04822_),
    .S(_04920_),
    .X(_04934_));
 sky130_fd_sc_hd__clkbuf_1 _09622_ (.A(_04934_),
    .X(_00077_));
 sky130_fd_sc_hd__mux2_1 _09623_ (.A0(net265),
    .A1(_04824_),
    .S(_04920_),
    .X(_04935_));
 sky130_fd_sc_hd__clkbuf_1 _09624_ (.A(_04935_),
    .X(_00078_));
 sky130_fd_sc_hd__mux2_1 _09625_ (.A0(net1089),
    .A1(_04826_),
    .S(_04920_),
    .X(_04936_));
 sky130_fd_sc_hd__clkbuf_1 _09626_ (.A(_04936_),
    .X(_00079_));
 sky130_fd_sc_hd__mux2_1 _09627_ (.A0(net1868),
    .A1(_04828_),
    .S(_04920_),
    .X(_04937_));
 sky130_fd_sc_hd__clkbuf_1 _09628_ (.A(_04937_),
    .X(_00080_));
 sky130_fd_sc_hd__nor2_4 _09629_ (.A(_04225_),
    .B(_04368_),
    .Y(_04938_));
 sky130_fd_sc_hd__clkbuf_4 _09630_ (.A(_04938_),
    .X(_04939_));
 sky130_fd_sc_hd__mux2_1 _09631_ (.A0(net2069),
    .A1(_04795_),
    .S(_04939_),
    .X(_04940_));
 sky130_fd_sc_hd__clkbuf_1 _09632_ (.A(_04940_),
    .X(_00081_));
 sky130_fd_sc_hd__mux2_1 _09633_ (.A0(net1991),
    .A1(_04800_),
    .S(_04939_),
    .X(_04941_));
 sky130_fd_sc_hd__clkbuf_1 _09634_ (.A(_04941_),
    .X(_00082_));
 sky130_fd_sc_hd__mux2_1 _09635_ (.A0(net2066),
    .A1(_04802_),
    .S(_04939_),
    .X(_04942_));
 sky130_fd_sc_hd__clkbuf_1 _09636_ (.A(_04942_),
    .X(_00083_));
 sky130_fd_sc_hd__mux2_1 _09637_ (.A0(net2028),
    .A1(_04804_),
    .S(_04939_),
    .X(_04943_));
 sky130_fd_sc_hd__clkbuf_1 _09638_ (.A(_04943_),
    .X(_00084_));
 sky130_fd_sc_hd__mux2_1 _09639_ (.A0(net1594),
    .A1(_04806_),
    .S(_04939_),
    .X(_04944_));
 sky130_fd_sc_hd__clkbuf_1 _09640_ (.A(_04944_),
    .X(_00085_));
 sky130_fd_sc_hd__mux2_1 _09641_ (.A0(net1894),
    .A1(_04808_),
    .S(_04939_),
    .X(_04945_));
 sky130_fd_sc_hd__clkbuf_1 _09642_ (.A(_04945_),
    .X(_00086_));
 sky130_fd_sc_hd__mux2_1 _09643_ (.A0(net1917),
    .A1(_04810_),
    .S(_04939_),
    .X(_04946_));
 sky130_fd_sc_hd__clkbuf_1 _09644_ (.A(_04946_),
    .X(_00087_));
 sky130_fd_sc_hd__mux2_1 _09645_ (.A0(net1867),
    .A1(_04812_),
    .S(_04939_),
    .X(_04947_));
 sky130_fd_sc_hd__clkbuf_1 _09646_ (.A(_04947_),
    .X(_00088_));
 sky130_fd_sc_hd__mux2_1 _09647_ (.A0(net1840),
    .A1(_04814_),
    .S(_04939_),
    .X(_04948_));
 sky130_fd_sc_hd__clkbuf_1 _09648_ (.A(_04948_),
    .X(_00089_));
 sky130_fd_sc_hd__mux2_1 _09649_ (.A0(net2020),
    .A1(_04816_),
    .S(_04939_),
    .X(_04949_));
 sky130_fd_sc_hd__clkbuf_1 _09650_ (.A(_04949_),
    .X(_00090_));
 sky130_fd_sc_hd__mux2_1 _09651_ (.A0(net2074),
    .A1(_04818_),
    .S(_04938_),
    .X(_04950_));
 sky130_fd_sc_hd__clkbuf_1 _09652_ (.A(_04950_),
    .X(_00091_));
 sky130_fd_sc_hd__mux2_1 _09653_ (.A0(net2062),
    .A1(_04820_),
    .S(_04938_),
    .X(_04951_));
 sky130_fd_sc_hd__clkbuf_1 _09654_ (.A(_04951_),
    .X(_00092_));
 sky130_fd_sc_hd__mux2_1 _09655_ (.A0(net2080),
    .A1(_04822_),
    .S(_04938_),
    .X(_04952_));
 sky130_fd_sc_hd__clkbuf_1 _09656_ (.A(_04952_),
    .X(_00093_));
 sky130_fd_sc_hd__mux2_1 _09657_ (.A0(net2015),
    .A1(_04824_),
    .S(_04938_),
    .X(_04953_));
 sky130_fd_sc_hd__clkbuf_1 _09658_ (.A(_04953_),
    .X(_00094_));
 sky130_fd_sc_hd__mux2_1 _09659_ (.A0(net2087),
    .A1(_04826_),
    .S(_04938_),
    .X(_04954_));
 sky130_fd_sc_hd__clkbuf_1 _09660_ (.A(_04954_),
    .X(_00095_));
 sky130_fd_sc_hd__mux2_1 _09661_ (.A0(net2079),
    .A1(_04828_),
    .S(_04938_),
    .X(_04955_));
 sky130_fd_sc_hd__clkbuf_1 _09662_ (.A(_04955_),
    .X(_00096_));
 sky130_fd_sc_hd__nor2_4 _09663_ (.A(_04796_),
    .B(_04646_),
    .Y(_04956_));
 sky130_fd_sc_hd__buf_6 _09664_ (.A(_04956_),
    .X(_04957_));
 sky130_fd_sc_hd__mux2_1 _09665_ (.A0(net389),
    .A1(_04795_),
    .S(_04957_),
    .X(_04958_));
 sky130_fd_sc_hd__clkbuf_1 _09666_ (.A(_04958_),
    .X(_00097_));
 sky130_fd_sc_hd__mux2_1 _09667_ (.A0(net732),
    .A1(_04800_),
    .S(_04957_),
    .X(_04959_));
 sky130_fd_sc_hd__clkbuf_1 _09668_ (.A(_04959_),
    .X(_00098_));
 sky130_fd_sc_hd__mux2_1 _09669_ (.A0(net198),
    .A1(_04802_),
    .S(_04957_),
    .X(_04960_));
 sky130_fd_sc_hd__clkbuf_1 _09670_ (.A(_04960_),
    .X(_00099_));
 sky130_fd_sc_hd__mux2_1 _09671_ (.A0(net232),
    .A1(_04804_),
    .S(_04957_),
    .X(_04961_));
 sky130_fd_sc_hd__clkbuf_1 _09672_ (.A(_04961_),
    .X(_00100_));
 sky130_fd_sc_hd__mux2_1 _09673_ (.A0(net1076),
    .A1(_04806_),
    .S(_04957_),
    .X(_04962_));
 sky130_fd_sc_hd__clkbuf_1 _09674_ (.A(_04962_),
    .X(_00101_));
 sky130_fd_sc_hd__mux2_1 _09675_ (.A0(net850),
    .A1(_04808_),
    .S(_04957_),
    .X(_04963_));
 sky130_fd_sc_hd__clkbuf_1 _09676_ (.A(_04963_),
    .X(_00102_));
 sky130_fd_sc_hd__mux2_1 _09677_ (.A0(net174),
    .A1(_04810_),
    .S(_04957_),
    .X(_04964_));
 sky130_fd_sc_hd__clkbuf_1 _09678_ (.A(_04964_),
    .X(_00103_));
 sky130_fd_sc_hd__mux2_1 _09679_ (.A0(net176),
    .A1(_04812_),
    .S(_04957_),
    .X(_04965_));
 sky130_fd_sc_hd__clkbuf_1 _09680_ (.A(_04965_),
    .X(_00104_));
 sky130_fd_sc_hd__mux2_1 _09681_ (.A0(net659),
    .A1(_04814_),
    .S(_04957_),
    .X(_04966_));
 sky130_fd_sc_hd__clkbuf_1 _09682_ (.A(_04966_),
    .X(_00105_));
 sky130_fd_sc_hd__mux2_1 _09683_ (.A0(net272),
    .A1(_04816_),
    .S(_04957_),
    .X(_04967_));
 sky130_fd_sc_hd__clkbuf_1 _09684_ (.A(_04967_),
    .X(_00106_));
 sky130_fd_sc_hd__mux2_1 _09685_ (.A0(net1331),
    .A1(_04818_),
    .S(_04956_),
    .X(_04968_));
 sky130_fd_sc_hd__clkbuf_1 _09686_ (.A(_04968_),
    .X(_00107_));
 sky130_fd_sc_hd__mux2_1 _09687_ (.A0(net513),
    .A1(_04820_),
    .S(_04956_),
    .X(_04969_));
 sky130_fd_sc_hd__clkbuf_1 _09688_ (.A(_04969_),
    .X(_00108_));
 sky130_fd_sc_hd__mux2_1 _09689_ (.A0(net469),
    .A1(_04822_),
    .S(_04956_),
    .X(_04970_));
 sky130_fd_sc_hd__clkbuf_1 _09690_ (.A(_04970_),
    .X(_00109_));
 sky130_fd_sc_hd__mux2_1 _09691_ (.A0(net366),
    .A1(_04824_),
    .S(_04956_),
    .X(_04971_));
 sky130_fd_sc_hd__clkbuf_1 _09692_ (.A(_04971_),
    .X(_00110_));
 sky130_fd_sc_hd__mux2_1 _09693_ (.A0(net477),
    .A1(_04826_),
    .S(_04956_),
    .X(_04972_));
 sky130_fd_sc_hd__clkbuf_1 _09694_ (.A(_04972_),
    .X(_00111_));
 sky130_fd_sc_hd__mux2_1 _09695_ (.A0(net1962),
    .A1(_04828_),
    .S(_04956_),
    .X(_04973_));
 sky130_fd_sc_hd__clkbuf_1 _09696_ (.A(_04973_),
    .X(_00112_));
 sky130_fd_sc_hd__nor2_4 _09697_ (.A(_04127_),
    .B(_04796_),
    .Y(_04974_));
 sky130_fd_sc_hd__buf_6 _09698_ (.A(_04974_),
    .X(_04975_));
 sky130_fd_sc_hd__mux2_1 _09699_ (.A0(net539),
    .A1(_04795_),
    .S(_04975_),
    .X(_04976_));
 sky130_fd_sc_hd__clkbuf_1 _09700_ (.A(_04976_),
    .X(_00113_));
 sky130_fd_sc_hd__mux2_1 _09701_ (.A0(net281),
    .A1(_04800_),
    .S(_04975_),
    .X(_04977_));
 sky130_fd_sc_hd__clkbuf_1 _09702_ (.A(_04977_),
    .X(_00114_));
 sky130_fd_sc_hd__mux2_1 _09703_ (.A0(net758),
    .A1(_04802_),
    .S(_04975_),
    .X(_04978_));
 sky130_fd_sc_hd__clkbuf_1 _09704_ (.A(_04978_),
    .X(_00115_));
 sky130_fd_sc_hd__mux2_1 _09705_ (.A0(net225),
    .A1(_04804_),
    .S(_04975_),
    .X(_04979_));
 sky130_fd_sc_hd__clkbuf_1 _09706_ (.A(_04979_),
    .X(_00116_));
 sky130_fd_sc_hd__mux2_1 _09707_ (.A0(net104),
    .A1(_04806_),
    .S(_04975_),
    .X(_04980_));
 sky130_fd_sc_hd__clkbuf_1 _09708_ (.A(_04980_),
    .X(_00117_));
 sky130_fd_sc_hd__mux2_1 _09709_ (.A0(net1532),
    .A1(_04808_),
    .S(_04975_),
    .X(_04981_));
 sky130_fd_sc_hd__clkbuf_1 _09710_ (.A(_04981_),
    .X(_00118_));
 sky130_fd_sc_hd__mux2_1 _09711_ (.A0(net734),
    .A1(_04810_),
    .S(_04975_),
    .X(_04982_));
 sky130_fd_sc_hd__clkbuf_1 _09712_ (.A(_04982_),
    .X(_00119_));
 sky130_fd_sc_hd__mux2_1 _09713_ (.A0(net483),
    .A1(_04812_),
    .S(_04975_),
    .X(_04983_));
 sky130_fd_sc_hd__clkbuf_1 _09714_ (.A(_04983_),
    .X(_00120_));
 sky130_fd_sc_hd__mux2_1 _09715_ (.A0(net234),
    .A1(_04814_),
    .S(_04975_),
    .X(_04984_));
 sky130_fd_sc_hd__clkbuf_1 _09716_ (.A(_04984_),
    .X(_00121_));
 sky130_fd_sc_hd__mux2_1 _09717_ (.A0(net236),
    .A1(_04816_),
    .S(_04975_),
    .X(_04985_));
 sky130_fd_sc_hd__clkbuf_1 _09718_ (.A(_04985_),
    .X(_00122_));
 sky130_fd_sc_hd__mux2_1 _09719_ (.A0(net400),
    .A1(_04818_),
    .S(_04974_),
    .X(_04986_));
 sky130_fd_sc_hd__clkbuf_1 _09720_ (.A(_04986_),
    .X(_00123_));
 sky130_fd_sc_hd__mux2_1 _09721_ (.A0(net464),
    .A1(_04820_),
    .S(_04974_),
    .X(_04987_));
 sky130_fd_sc_hd__clkbuf_1 _09722_ (.A(_04987_),
    .X(_00124_));
 sky130_fd_sc_hd__mux2_1 _09723_ (.A0(net84),
    .A1(_04822_),
    .S(_04974_),
    .X(_04988_));
 sky130_fd_sc_hd__clkbuf_1 _09724_ (.A(_04988_),
    .X(_00125_));
 sky130_fd_sc_hd__mux2_1 _09725_ (.A0(net269),
    .A1(_04824_),
    .S(_04974_),
    .X(_04989_));
 sky130_fd_sc_hd__clkbuf_1 _09726_ (.A(_04989_),
    .X(_00126_));
 sky130_fd_sc_hd__mux2_1 _09727_ (.A0(net323),
    .A1(_04826_),
    .S(_04974_),
    .X(_04990_));
 sky130_fd_sc_hd__clkbuf_1 _09728_ (.A(_04990_),
    .X(_00127_));
 sky130_fd_sc_hd__mux2_1 _09729_ (.A0(net245),
    .A1(_04828_),
    .S(_04974_),
    .X(_04991_));
 sky130_fd_sc_hd__clkbuf_1 _09730_ (.A(_04991_),
    .X(_00128_));
 sky130_fd_sc_hd__buf_8 _09731_ (.A(_04069_),
    .X(_04992_));
 sky130_fd_sc_hd__nor2_4 _09732_ (.A(_04796_),
    .B(_04684_),
    .Y(_04993_));
 sky130_fd_sc_hd__buf_6 _09733_ (.A(_04993_),
    .X(_04994_));
 sky130_fd_sc_hd__mux2_1 _09734_ (.A0(net179),
    .A1(_04992_),
    .S(_04994_),
    .X(_04995_));
 sky130_fd_sc_hd__clkbuf_1 _09735_ (.A(_04995_),
    .X(_00129_));
 sky130_fd_sc_hd__buf_6 _09736_ (.A(_04080_),
    .X(_04996_));
 sky130_fd_sc_hd__mux2_1 _09737_ (.A0(net1260),
    .A1(_04996_),
    .S(_04994_),
    .X(_04997_));
 sky130_fd_sc_hd__clkbuf_1 _09738_ (.A(_04997_),
    .X(_00130_));
 sky130_fd_sc_hd__clkbuf_16 _09739_ (.A(_04083_),
    .X(_04998_));
 sky130_fd_sc_hd__mux2_1 _09740_ (.A0(net907),
    .A1(_04998_),
    .S(_04994_),
    .X(_04999_));
 sky130_fd_sc_hd__clkbuf_1 _09741_ (.A(_04999_),
    .X(_00131_));
 sky130_fd_sc_hd__buf_8 _09742_ (.A(_04086_),
    .X(_05000_));
 sky130_fd_sc_hd__mux2_1 _09743_ (.A0(net247),
    .A1(_05000_),
    .S(_04994_),
    .X(_05001_));
 sky130_fd_sc_hd__clkbuf_1 _09744_ (.A(_05001_),
    .X(_00132_));
 sky130_fd_sc_hd__buf_8 _09745_ (.A(_04089_),
    .X(_05002_));
 sky130_fd_sc_hd__mux2_1 _09746_ (.A0(net795),
    .A1(_05002_),
    .S(_04994_),
    .X(_05003_));
 sky130_fd_sc_hd__clkbuf_1 _09747_ (.A(_05003_),
    .X(_00133_));
 sky130_fd_sc_hd__buf_6 _09748_ (.A(_04092_),
    .X(_05004_));
 sky130_fd_sc_hd__mux2_1 _09749_ (.A0(net338),
    .A1(_05004_),
    .S(_04994_),
    .X(_05005_));
 sky130_fd_sc_hd__clkbuf_1 _09750_ (.A(_05005_),
    .X(_00134_));
 sky130_fd_sc_hd__buf_8 _09751_ (.A(_04095_),
    .X(_05006_));
 sky130_fd_sc_hd__mux2_1 _09752_ (.A0(net164),
    .A1(_05006_),
    .S(_04994_),
    .X(_05007_));
 sky130_fd_sc_hd__clkbuf_1 _09753_ (.A(_05007_),
    .X(_00135_));
 sky130_fd_sc_hd__buf_8 _09754_ (.A(_04098_),
    .X(_05008_));
 sky130_fd_sc_hd__mux2_1 _09755_ (.A0(net41),
    .A1(_05008_),
    .S(_04994_),
    .X(_05009_));
 sky130_fd_sc_hd__clkbuf_1 _09756_ (.A(_05009_),
    .X(_00136_));
 sky130_fd_sc_hd__buf_8 _09757_ (.A(_04101_),
    .X(_05010_));
 sky130_fd_sc_hd__mux2_1 _09758_ (.A0(net301),
    .A1(_05010_),
    .S(_04994_),
    .X(_05011_));
 sky130_fd_sc_hd__clkbuf_1 _09759_ (.A(_05011_),
    .X(_00137_));
 sky130_fd_sc_hd__buf_8 _09760_ (.A(_04104_),
    .X(_05012_));
 sky130_fd_sc_hd__mux2_1 _09761_ (.A0(net398),
    .A1(_05012_),
    .S(_04994_),
    .X(_05013_));
 sky130_fd_sc_hd__clkbuf_1 _09762_ (.A(_05013_),
    .X(_00138_));
 sky130_fd_sc_hd__buf_8 _09763_ (.A(_04107_),
    .X(_05014_));
 sky130_fd_sc_hd__mux2_1 _09764_ (.A0(net287),
    .A1(_05014_),
    .S(_04993_),
    .X(_05015_));
 sky130_fd_sc_hd__clkbuf_1 _09765_ (.A(_05015_),
    .X(_00139_));
 sky130_fd_sc_hd__buf_8 _09766_ (.A(_04110_),
    .X(_05016_));
 sky130_fd_sc_hd__mux2_1 _09767_ (.A0(net497),
    .A1(_05016_),
    .S(_04993_),
    .X(_05017_));
 sky130_fd_sc_hd__clkbuf_1 _09768_ (.A(_05017_),
    .X(_00140_));
 sky130_fd_sc_hd__buf_8 _09769_ (.A(_04113_),
    .X(_05018_));
 sky130_fd_sc_hd__mux2_1 _09770_ (.A0(net1372),
    .A1(_05018_),
    .S(_04993_),
    .X(_05019_));
 sky130_fd_sc_hd__clkbuf_1 _09771_ (.A(_05019_),
    .X(_00141_));
 sky130_fd_sc_hd__buf_6 _09772_ (.A(_04116_),
    .X(_05020_));
 sky130_fd_sc_hd__mux2_1 _09773_ (.A0(net1064),
    .A1(_05020_),
    .S(_04993_),
    .X(_05021_));
 sky130_fd_sc_hd__clkbuf_1 _09774_ (.A(_05021_),
    .X(_00142_));
 sky130_fd_sc_hd__buf_8 _09775_ (.A(_04119_),
    .X(_05022_));
 sky130_fd_sc_hd__mux2_1 _09776_ (.A0(net1613),
    .A1(_05022_),
    .S(_04993_),
    .X(_05023_));
 sky130_fd_sc_hd__clkbuf_1 _09777_ (.A(_05023_),
    .X(_00143_));
 sky130_fd_sc_hd__buf_6 _09778_ (.A(_04122_),
    .X(_05024_));
 sky130_fd_sc_hd__mux2_1 _09779_ (.A0(net743),
    .A1(_05024_),
    .S(_04993_),
    .X(_05025_));
 sky130_fd_sc_hd__clkbuf_1 _09780_ (.A(_05025_),
    .X(_00144_));
 sky130_fd_sc_hd__buf_6 _09781_ (.A(_02442_),
    .X(_05026_));
 sky130_fd_sc_hd__or3_1 _09782_ (.A(_02707_),
    .B(_05026_),
    .C(_04246_),
    .X(_05027_));
 sky130_fd_sc_hd__clkbuf_4 _09783_ (.A(_05027_),
    .X(_05028_));
 sky130_fd_sc_hd__buf_6 _09784_ (.A(_05028_),
    .X(_05029_));
 sky130_fd_sc_hd__mux2_1 _09785_ (.A0(_04406_),
    .A1(net646),
    .S(_05029_),
    .X(_05030_));
 sky130_fd_sc_hd__clkbuf_1 _09786_ (.A(_05030_),
    .X(_00145_));
 sky130_fd_sc_hd__mux2_1 _09787_ (.A0(_04412_),
    .A1(net1809),
    .S(_05029_),
    .X(_05031_));
 sky130_fd_sc_hd__clkbuf_1 _09788_ (.A(_05031_),
    .X(_00146_));
 sky130_fd_sc_hd__mux2_1 _09789_ (.A0(_04414_),
    .A1(net1350),
    .S(_05029_),
    .X(_05032_));
 sky130_fd_sc_hd__clkbuf_1 _09790_ (.A(_05032_),
    .X(_00147_));
 sky130_fd_sc_hd__mux2_1 _09791_ (.A0(_04416_),
    .A1(net1869),
    .S(_05029_),
    .X(_05033_));
 sky130_fd_sc_hd__clkbuf_1 _09792_ (.A(_05033_),
    .X(_00148_));
 sky130_fd_sc_hd__mux2_1 _09793_ (.A0(_04418_),
    .A1(net1404),
    .S(_05029_),
    .X(_05034_));
 sky130_fd_sc_hd__clkbuf_1 _09794_ (.A(_05034_),
    .X(_00149_));
 sky130_fd_sc_hd__mux2_1 _09795_ (.A0(_04420_),
    .A1(net1446),
    .S(_05029_),
    .X(_05035_));
 sky130_fd_sc_hd__clkbuf_1 _09796_ (.A(_05035_),
    .X(_00150_));
 sky130_fd_sc_hd__mux2_1 _09797_ (.A0(_04422_),
    .A1(net1147),
    .S(_05029_),
    .X(_05036_));
 sky130_fd_sc_hd__clkbuf_1 _09798_ (.A(_05036_),
    .X(_00151_));
 sky130_fd_sc_hd__mux2_1 _09799_ (.A0(_04424_),
    .A1(net1393),
    .S(_05029_),
    .X(_05037_));
 sky130_fd_sc_hd__clkbuf_1 _09800_ (.A(_05037_),
    .X(_00152_));
 sky130_fd_sc_hd__mux2_1 _09801_ (.A0(_04426_),
    .A1(net603),
    .S(_05029_),
    .X(_05038_));
 sky130_fd_sc_hd__clkbuf_1 _09802_ (.A(_05038_),
    .X(_00153_));
 sky130_fd_sc_hd__mux2_1 _09803_ (.A0(_04428_),
    .A1(net649),
    .S(_05029_),
    .X(_05039_));
 sky130_fd_sc_hd__clkbuf_1 _09804_ (.A(_05039_),
    .X(_00154_));
 sky130_fd_sc_hd__mux2_1 _09805_ (.A0(_04430_),
    .A1(net1910),
    .S(_05028_),
    .X(_05040_));
 sky130_fd_sc_hd__clkbuf_1 _09806_ (.A(_05040_),
    .X(_00155_));
 sky130_fd_sc_hd__mux2_1 _09807_ (.A0(_04432_),
    .A1(net1168),
    .S(_05028_),
    .X(_05041_));
 sky130_fd_sc_hd__clkbuf_1 _09808_ (.A(_05041_),
    .X(_00156_));
 sky130_fd_sc_hd__mux2_1 _09809_ (.A0(_04434_),
    .A1(net1086),
    .S(_05028_),
    .X(_05042_));
 sky130_fd_sc_hd__clkbuf_1 _09810_ (.A(_05042_),
    .X(_00157_));
 sky130_fd_sc_hd__mux2_1 _09811_ (.A0(_04436_),
    .A1(net906),
    .S(_05028_),
    .X(_05043_));
 sky130_fd_sc_hd__clkbuf_1 _09812_ (.A(_05043_),
    .X(_00158_));
 sky130_fd_sc_hd__mux2_1 _09813_ (.A0(_04438_),
    .A1(net786),
    .S(_05028_),
    .X(_05044_));
 sky130_fd_sc_hd__clkbuf_1 _09814_ (.A(_05044_),
    .X(_00159_));
 sky130_fd_sc_hd__mux2_1 _09815_ (.A0(_04440_),
    .A1(net598),
    .S(_05028_),
    .X(_05045_));
 sky130_fd_sc_hd__clkbuf_1 _09816_ (.A(_05045_),
    .X(_00160_));
 sky130_fd_sc_hd__nor2_4 _09817_ (.A(_04246_),
    .B(_04365_),
    .Y(_05046_));
 sky130_fd_sc_hd__buf_6 _09818_ (.A(_05046_),
    .X(_05047_));
 sky130_fd_sc_hd__mux2_1 _09819_ (.A0(net178),
    .A1(_04992_),
    .S(_05047_),
    .X(_05048_));
 sky130_fd_sc_hd__clkbuf_1 _09820_ (.A(_05048_),
    .X(_00161_));
 sky130_fd_sc_hd__mux2_1 _09821_ (.A0(net759),
    .A1(_04996_),
    .S(_05047_),
    .X(_05049_));
 sky130_fd_sc_hd__clkbuf_1 _09822_ (.A(_05049_),
    .X(_00162_));
 sky130_fd_sc_hd__mux2_1 _09823_ (.A0(net904),
    .A1(_04998_),
    .S(_05047_),
    .X(_05050_));
 sky130_fd_sc_hd__clkbuf_1 _09824_ (.A(_05050_),
    .X(_00163_));
 sky130_fd_sc_hd__mux2_1 _09825_ (.A0(net1439),
    .A1(_05000_),
    .S(_05047_),
    .X(_05051_));
 sky130_fd_sc_hd__clkbuf_1 _09826_ (.A(_05051_),
    .X(_00164_));
 sky130_fd_sc_hd__mux2_1 _09827_ (.A0(net840),
    .A1(_05002_),
    .S(_05047_),
    .X(_05052_));
 sky130_fd_sc_hd__clkbuf_1 _09828_ (.A(_05052_),
    .X(_00165_));
 sky130_fd_sc_hd__mux2_1 _09829_ (.A0(net87),
    .A1(_05004_),
    .S(_05047_),
    .X(_05053_));
 sky130_fd_sc_hd__clkbuf_1 _09830_ (.A(_05053_),
    .X(_00166_));
 sky130_fd_sc_hd__mux2_1 _09831_ (.A0(net1364),
    .A1(_05006_),
    .S(_05047_),
    .X(_05054_));
 sky130_fd_sc_hd__clkbuf_1 _09832_ (.A(_05054_),
    .X(_00167_));
 sky130_fd_sc_hd__mux2_1 _09833_ (.A0(net845),
    .A1(_05008_),
    .S(_05047_),
    .X(_05055_));
 sky130_fd_sc_hd__clkbuf_1 _09834_ (.A(_05055_),
    .X(_00168_));
 sky130_fd_sc_hd__mux2_1 _09835_ (.A0(net1899),
    .A1(_05010_),
    .S(_05047_),
    .X(_05056_));
 sky130_fd_sc_hd__clkbuf_1 _09836_ (.A(_05056_),
    .X(_00169_));
 sky130_fd_sc_hd__mux2_1 _09837_ (.A0(net589),
    .A1(_05012_),
    .S(_05047_),
    .X(_05057_));
 sky130_fd_sc_hd__clkbuf_1 _09838_ (.A(_05057_),
    .X(_00170_));
 sky130_fd_sc_hd__mux2_1 _09839_ (.A0(net536),
    .A1(_05014_),
    .S(_05046_),
    .X(_05058_));
 sky130_fd_sc_hd__clkbuf_1 _09840_ (.A(_05058_),
    .X(_00171_));
 sky130_fd_sc_hd__mux2_1 _09841_ (.A0(net524),
    .A1(_05016_),
    .S(_05046_),
    .X(_05059_));
 sky130_fd_sc_hd__clkbuf_1 _09842_ (.A(_05059_),
    .X(_00172_));
 sky130_fd_sc_hd__mux2_1 _09843_ (.A0(net402),
    .A1(_05018_),
    .S(_05046_),
    .X(_05060_));
 sky130_fd_sc_hd__clkbuf_1 _09844_ (.A(_05060_),
    .X(_00173_));
 sky130_fd_sc_hd__mux2_1 _09845_ (.A0(net653),
    .A1(_05020_),
    .S(_05046_),
    .X(_05061_));
 sky130_fd_sc_hd__clkbuf_1 _09846_ (.A(_05061_),
    .X(_00174_));
 sky130_fd_sc_hd__mux2_1 _09847_ (.A0(net487),
    .A1(_05022_),
    .S(_05046_),
    .X(_05062_));
 sky130_fd_sc_hd__clkbuf_1 _09848_ (.A(_05062_),
    .X(_00175_));
 sky130_fd_sc_hd__mux2_1 _09849_ (.A0(net337),
    .A1(_05024_),
    .S(_05046_),
    .X(_05063_));
 sky130_fd_sc_hd__clkbuf_1 _09850_ (.A(_05063_),
    .X(_00176_));
 sky130_fd_sc_hd__or3_1 _09851_ (.A(_04059_),
    .B(_02737_),
    .C(_04246_),
    .X(_05064_));
 sky130_fd_sc_hd__clkbuf_4 _09852_ (.A(_05064_),
    .X(_05065_));
 sky130_fd_sc_hd__buf_6 _09853_ (.A(_05065_),
    .X(_05066_));
 sky130_fd_sc_hd__mux2_1 _09854_ (.A0(_04406_),
    .A1(net616),
    .S(_05066_),
    .X(_05067_));
 sky130_fd_sc_hd__clkbuf_1 _09855_ (.A(_05067_),
    .X(_00177_));
 sky130_fd_sc_hd__mux2_1 _09856_ (.A0(_04412_),
    .A1(net741),
    .S(_05066_),
    .X(_05068_));
 sky130_fd_sc_hd__clkbuf_1 _09857_ (.A(_05068_),
    .X(_00178_));
 sky130_fd_sc_hd__mux2_1 _09858_ (.A0(_04414_),
    .A1(net565),
    .S(_05066_),
    .X(_05069_));
 sky130_fd_sc_hd__clkbuf_1 _09859_ (.A(_05069_),
    .X(_00179_));
 sky130_fd_sc_hd__mux2_1 _09860_ (.A0(_04416_),
    .A1(net133),
    .S(_05066_),
    .X(_05070_));
 sky130_fd_sc_hd__clkbuf_1 _09861_ (.A(_05070_),
    .X(_00180_));
 sky130_fd_sc_hd__mux2_1 _09862_ (.A0(_04418_),
    .A1(net950),
    .S(_05066_),
    .X(_05071_));
 sky130_fd_sc_hd__clkbuf_1 _09863_ (.A(_05071_),
    .X(_00181_));
 sky130_fd_sc_hd__mux2_1 _09864_ (.A0(_04420_),
    .A1(net496),
    .S(_05066_),
    .X(_05072_));
 sky130_fd_sc_hd__clkbuf_1 _09865_ (.A(_05072_),
    .X(_00182_));
 sky130_fd_sc_hd__mux2_1 _09866_ (.A0(_04422_),
    .A1(net282),
    .S(_05066_),
    .X(_05073_));
 sky130_fd_sc_hd__clkbuf_1 _09867_ (.A(_05073_),
    .X(_00183_));
 sky130_fd_sc_hd__mux2_1 _09868_ (.A0(_04424_),
    .A1(net730),
    .S(_05066_),
    .X(_05074_));
 sky130_fd_sc_hd__clkbuf_1 _09869_ (.A(_05074_),
    .X(_00184_));
 sky130_fd_sc_hd__mux2_1 _09870_ (.A0(_04426_),
    .A1(net849),
    .S(_05066_),
    .X(_05075_));
 sky130_fd_sc_hd__clkbuf_1 _09871_ (.A(_05075_),
    .X(_00185_));
 sky130_fd_sc_hd__mux2_1 _09872_ (.A0(_04428_),
    .A1(net382),
    .S(_05066_),
    .X(_05076_));
 sky130_fd_sc_hd__clkbuf_1 _09873_ (.A(_05076_),
    .X(_00186_));
 sky130_fd_sc_hd__mux2_1 _09874_ (.A0(_04430_),
    .A1(net1496),
    .S(_05065_),
    .X(_05077_));
 sky130_fd_sc_hd__clkbuf_1 _09875_ (.A(_05077_),
    .X(_00187_));
 sky130_fd_sc_hd__mux2_1 _09876_ (.A0(_04432_),
    .A1(net503),
    .S(_05065_),
    .X(_05078_));
 sky130_fd_sc_hd__clkbuf_1 _09877_ (.A(_05078_),
    .X(_00188_));
 sky130_fd_sc_hd__mux2_1 _09878_ (.A0(_04434_),
    .A1(net381),
    .S(_05065_),
    .X(_05079_));
 sky130_fd_sc_hd__clkbuf_1 _09879_ (.A(_05079_),
    .X(_00189_));
 sky130_fd_sc_hd__mux2_1 _09880_ (.A0(_04436_),
    .A1(net1557),
    .S(_05065_),
    .X(_05080_));
 sky130_fd_sc_hd__clkbuf_1 _09881_ (.A(_05080_),
    .X(_00190_));
 sky130_fd_sc_hd__mux2_1 _09882_ (.A0(_04438_),
    .A1(net1681),
    .S(_05065_),
    .X(_05081_));
 sky130_fd_sc_hd__clkbuf_1 _09883_ (.A(_05081_),
    .X(_00191_));
 sky130_fd_sc_hd__mux2_1 _09884_ (.A0(_04440_),
    .A1(net394),
    .S(_05065_),
    .X(_05082_));
 sky130_fd_sc_hd__clkbuf_1 _09885_ (.A(_05082_),
    .X(_00192_));
 sky130_fd_sc_hd__nand2b_4 _09886_ (.A_N(_04246_),
    .B(_04408_),
    .Y(_05083_));
 sky130_fd_sc_hd__buf_6 _09887_ (.A(_05083_),
    .X(_05084_));
 sky130_fd_sc_hd__mux2_1 _09888_ (.A0(_04406_),
    .A1(net908),
    .S(_05084_),
    .X(_05085_));
 sky130_fd_sc_hd__clkbuf_1 _09889_ (.A(_05085_),
    .X(_00193_));
 sky130_fd_sc_hd__mux2_1 _09890_ (.A0(_04412_),
    .A1(net1254),
    .S(_05084_),
    .X(_05086_));
 sky130_fd_sc_hd__clkbuf_1 _09891_ (.A(_05086_),
    .X(_00194_));
 sky130_fd_sc_hd__mux2_1 _09892_ (.A0(_04414_),
    .A1(net1813),
    .S(_05084_),
    .X(_05087_));
 sky130_fd_sc_hd__clkbuf_1 _09893_ (.A(_05087_),
    .X(_00195_));
 sky130_fd_sc_hd__mux2_1 _09894_ (.A0(_04416_),
    .A1(net855),
    .S(_05084_),
    .X(_05088_));
 sky130_fd_sc_hd__clkbuf_1 _09895_ (.A(_05088_),
    .X(_00196_));
 sky130_fd_sc_hd__mux2_1 _09896_ (.A0(_04418_),
    .A1(net1190),
    .S(_05084_),
    .X(_05089_));
 sky130_fd_sc_hd__clkbuf_1 _09897_ (.A(_05089_),
    .X(_00197_));
 sky130_fd_sc_hd__mux2_1 _09898_ (.A0(_04420_),
    .A1(net1352),
    .S(_05084_),
    .X(_05090_));
 sky130_fd_sc_hd__clkbuf_1 _09899_ (.A(_05090_),
    .X(_00198_));
 sky130_fd_sc_hd__mux2_1 _09900_ (.A0(_04422_),
    .A1(net678),
    .S(_05084_),
    .X(_05091_));
 sky130_fd_sc_hd__clkbuf_1 _09901_ (.A(_05091_),
    .X(_00199_));
 sky130_fd_sc_hd__mux2_1 _09902_ (.A0(_04424_),
    .A1(net1125),
    .S(_05084_),
    .X(_05092_));
 sky130_fd_sc_hd__clkbuf_1 _09903_ (.A(_05092_),
    .X(_00200_));
 sky130_fd_sc_hd__mux2_1 _09904_ (.A0(_04426_),
    .A1(net856),
    .S(_05084_),
    .X(_05093_));
 sky130_fd_sc_hd__clkbuf_1 _09905_ (.A(_05093_),
    .X(_00201_));
 sky130_fd_sc_hd__mux2_1 _09906_ (.A0(_04428_),
    .A1(net1471),
    .S(_05084_),
    .X(_05094_));
 sky130_fd_sc_hd__clkbuf_1 _09907_ (.A(_05094_),
    .X(_00202_));
 sky130_fd_sc_hd__mux2_1 _09908_ (.A0(_04430_),
    .A1(net533),
    .S(_05083_),
    .X(_05095_));
 sky130_fd_sc_hd__clkbuf_1 _09909_ (.A(_05095_),
    .X(_00203_));
 sky130_fd_sc_hd__mux2_1 _09910_ (.A0(_04432_),
    .A1(net1624),
    .S(_05083_),
    .X(_05096_));
 sky130_fd_sc_hd__clkbuf_1 _09911_ (.A(_05096_),
    .X(_00204_));
 sky130_fd_sc_hd__mux2_1 _09912_ (.A0(_04434_),
    .A1(net1195),
    .S(_05083_),
    .X(_05097_));
 sky130_fd_sc_hd__clkbuf_1 _09913_ (.A(_05097_),
    .X(_00205_));
 sky130_fd_sc_hd__mux2_1 _09914_ (.A0(_04436_),
    .A1(net986),
    .S(_05083_),
    .X(_05098_));
 sky130_fd_sc_hd__clkbuf_1 _09915_ (.A(_05098_),
    .X(_00206_));
 sky130_fd_sc_hd__mux2_1 _09916_ (.A0(_04438_),
    .A1(net1492),
    .S(_05083_),
    .X(_05099_));
 sky130_fd_sc_hd__clkbuf_1 _09917_ (.A(_05099_),
    .X(_00207_));
 sky130_fd_sc_hd__mux2_1 _09918_ (.A0(_04440_),
    .A1(net1327),
    .S(_05083_),
    .X(_05100_));
 sky130_fd_sc_hd__clkbuf_1 _09919_ (.A(_05100_),
    .X(_00208_));
 sky130_fd_sc_hd__or3_1 _09920_ (.A(_04059_),
    .B(_05026_),
    .C(_04246_),
    .X(_05101_));
 sky130_fd_sc_hd__clkbuf_4 _09921_ (.A(_05101_),
    .X(_05102_));
 sky130_fd_sc_hd__buf_6 _09922_ (.A(_05102_),
    .X(_05103_));
 sky130_fd_sc_hd__mux2_1 _09923_ (.A0(_04406_),
    .A1(net995),
    .S(_05103_),
    .X(_05104_));
 sky130_fd_sc_hd__clkbuf_1 _09924_ (.A(_05104_),
    .X(_00209_));
 sky130_fd_sc_hd__mux2_1 _09925_ (.A0(_04412_),
    .A1(net1617),
    .S(_05103_),
    .X(_05105_));
 sky130_fd_sc_hd__clkbuf_1 _09926_ (.A(_05105_),
    .X(_00210_));
 sky130_fd_sc_hd__mux2_1 _09927_ (.A0(_04414_),
    .A1(net1538),
    .S(_05103_),
    .X(_05106_));
 sky130_fd_sc_hd__clkbuf_1 _09928_ (.A(_05106_),
    .X(_00211_));
 sky130_fd_sc_hd__mux2_1 _09929_ (.A0(_04416_),
    .A1(net1034),
    .S(_05103_),
    .X(_05107_));
 sky130_fd_sc_hd__clkbuf_1 _09930_ (.A(_05107_),
    .X(_00212_));
 sky130_fd_sc_hd__mux2_1 _09931_ (.A0(_04418_),
    .A1(net546),
    .S(_05103_),
    .X(_05108_));
 sky130_fd_sc_hd__clkbuf_1 _09932_ (.A(_05108_),
    .X(_00213_));
 sky130_fd_sc_hd__mux2_1 _09933_ (.A0(_04420_),
    .A1(net1610),
    .S(_05103_),
    .X(_05109_));
 sky130_fd_sc_hd__clkbuf_1 _09934_ (.A(_05109_),
    .X(_00214_));
 sky130_fd_sc_hd__mux2_1 _09935_ (.A0(_04422_),
    .A1(net534),
    .S(_05103_),
    .X(_05110_));
 sky130_fd_sc_hd__clkbuf_1 _09936_ (.A(_05110_),
    .X(_00215_));
 sky130_fd_sc_hd__mux2_1 _09937_ (.A0(_04424_),
    .A1(net905),
    .S(_05103_),
    .X(_05111_));
 sky130_fd_sc_hd__clkbuf_1 _09938_ (.A(_05111_),
    .X(_00216_));
 sky130_fd_sc_hd__mux2_1 _09939_ (.A0(_04426_),
    .A1(net1001),
    .S(_05103_),
    .X(_05112_));
 sky130_fd_sc_hd__clkbuf_1 _09940_ (.A(_05112_),
    .X(_00217_));
 sky130_fd_sc_hd__mux2_1 _09941_ (.A0(_04428_),
    .A1(net1247),
    .S(_05103_),
    .X(_05113_));
 sky130_fd_sc_hd__clkbuf_1 _09942_ (.A(_05113_),
    .X(_00218_));
 sky130_fd_sc_hd__mux2_1 _09943_ (.A0(_04430_),
    .A1(net304),
    .S(_05102_),
    .X(_05114_));
 sky130_fd_sc_hd__clkbuf_1 _09944_ (.A(_05114_),
    .X(_00219_));
 sky130_fd_sc_hd__mux2_1 _09945_ (.A0(_04432_),
    .A1(net1560),
    .S(_05102_),
    .X(_05115_));
 sky130_fd_sc_hd__clkbuf_1 _09946_ (.A(_05115_),
    .X(_00220_));
 sky130_fd_sc_hd__mux2_1 _09947_ (.A0(_04434_),
    .A1(net1146),
    .S(_05102_),
    .X(_05116_));
 sky130_fd_sc_hd__clkbuf_1 _09948_ (.A(_05116_),
    .X(_00221_));
 sky130_fd_sc_hd__mux2_1 _09949_ (.A0(_04436_),
    .A1(net1931),
    .S(_05102_),
    .X(_05117_));
 sky130_fd_sc_hd__clkbuf_1 _09950_ (.A(_05117_),
    .X(_00222_));
 sky130_fd_sc_hd__mux2_1 _09951_ (.A0(_04438_),
    .A1(net1798),
    .S(_05102_),
    .X(_05118_));
 sky130_fd_sc_hd__clkbuf_1 _09952_ (.A(_05118_),
    .X(_00223_));
 sky130_fd_sc_hd__mux2_1 _09953_ (.A0(_04440_),
    .A1(net880),
    .S(_05102_),
    .X(_05119_));
 sky130_fd_sc_hd__clkbuf_1 _09954_ (.A(_05119_),
    .X(_00224_));
 sky130_fd_sc_hd__nor2_4 _09955_ (.A(_04076_),
    .B(_04461_),
    .Y(_05120_));
 sky130_fd_sc_hd__buf_4 _09956_ (.A(_05120_),
    .X(_05121_));
 sky130_fd_sc_hd__mux2_1 _09957_ (.A0(net86),
    .A1(_04992_),
    .S(_05121_),
    .X(_05122_));
 sky130_fd_sc_hd__clkbuf_1 _09958_ (.A(_05122_),
    .X(_00225_));
 sky130_fd_sc_hd__mux2_1 _09959_ (.A0(net156),
    .A1(_04996_),
    .S(_05121_),
    .X(_05123_));
 sky130_fd_sc_hd__clkbuf_1 _09960_ (.A(_05123_),
    .X(_00226_));
 sky130_fd_sc_hd__mux2_1 _09961_ (.A0(net351),
    .A1(_04998_),
    .S(_05121_),
    .X(_05124_));
 sky130_fd_sc_hd__clkbuf_1 _09962_ (.A(_05124_),
    .X(_00227_));
 sky130_fd_sc_hd__mux2_1 _09963_ (.A0(net451),
    .A1(_05000_),
    .S(_05121_),
    .X(_05125_));
 sky130_fd_sc_hd__clkbuf_1 _09964_ (.A(_05125_),
    .X(_00228_));
 sky130_fd_sc_hd__mux2_1 _09965_ (.A0(net369),
    .A1(_05002_),
    .S(_05121_),
    .X(_05126_));
 sky130_fd_sc_hd__clkbuf_1 _09966_ (.A(_05126_),
    .X(_00229_));
 sky130_fd_sc_hd__mux2_1 _09967_ (.A0(net82),
    .A1(_05004_),
    .S(_05121_),
    .X(_05127_));
 sky130_fd_sc_hd__clkbuf_1 _09968_ (.A(_05127_),
    .X(_00230_));
 sky130_fd_sc_hd__mux2_1 _09969_ (.A0(net243),
    .A1(_05006_),
    .S(_05121_),
    .X(_05128_));
 sky130_fd_sc_hd__clkbuf_1 _09970_ (.A(_05128_),
    .X(_00231_));
 sky130_fd_sc_hd__mux2_1 _09971_ (.A0(net384),
    .A1(_05008_),
    .S(_05121_),
    .X(_05129_));
 sky130_fd_sc_hd__clkbuf_1 _09972_ (.A(_05129_),
    .X(_00232_));
 sky130_fd_sc_hd__mux2_1 _09973_ (.A0(net183),
    .A1(_05010_),
    .S(_05121_),
    .X(_05130_));
 sky130_fd_sc_hd__clkbuf_1 _09974_ (.A(_05130_),
    .X(_00233_));
 sky130_fd_sc_hd__mux2_1 _09975_ (.A0(net239),
    .A1(_05012_),
    .S(_05121_),
    .X(_05131_));
 sky130_fd_sc_hd__clkbuf_1 _09976_ (.A(_05131_),
    .X(_00234_));
 sky130_fd_sc_hd__mux2_1 _09977_ (.A0(net557),
    .A1(_05014_),
    .S(_05120_),
    .X(_05132_));
 sky130_fd_sc_hd__clkbuf_1 _09978_ (.A(_05132_),
    .X(_00235_));
 sky130_fd_sc_hd__mux2_1 _09979_ (.A0(net119),
    .A1(_05016_),
    .S(_05120_),
    .X(_05133_));
 sky130_fd_sc_hd__clkbuf_1 _09980_ (.A(_05133_),
    .X(_00236_));
 sky130_fd_sc_hd__mux2_1 _09981_ (.A0(net139),
    .A1(_05018_),
    .S(_05120_),
    .X(_05134_));
 sky130_fd_sc_hd__clkbuf_1 _09982_ (.A(_05134_),
    .X(_00237_));
 sky130_fd_sc_hd__mux2_1 _09983_ (.A0(net266),
    .A1(_05020_),
    .S(_05120_),
    .X(_05135_));
 sky130_fd_sc_hd__clkbuf_1 _09984_ (.A(_05135_),
    .X(_00238_));
 sky130_fd_sc_hd__mux2_1 _09985_ (.A0(net72),
    .A1(_05022_),
    .S(_05120_),
    .X(_05136_));
 sky130_fd_sc_hd__clkbuf_1 _09986_ (.A(_05136_),
    .X(_00239_));
 sky130_fd_sc_hd__mux2_1 _09987_ (.A0(net954),
    .A1(_05024_),
    .S(_05120_),
    .X(_05137_));
 sky130_fd_sc_hd__clkbuf_1 _09988_ (.A(_05137_),
    .X(_00240_));
 sky130_fd_sc_hd__nor2_4 _09989_ (.A(_04368_),
    .B(_04569_),
    .Y(_05138_));
 sky130_fd_sc_hd__buf_4 _09990_ (.A(_05138_),
    .X(_05139_));
 sky130_fd_sc_hd__mux2_1 _09991_ (.A0(net128),
    .A1(_04992_),
    .S(_05139_),
    .X(_05140_));
 sky130_fd_sc_hd__clkbuf_1 _09992_ (.A(_05140_),
    .X(_00241_));
 sky130_fd_sc_hd__mux2_1 _09993_ (.A0(net767),
    .A1(_04996_),
    .S(_05139_),
    .X(_05141_));
 sky130_fd_sc_hd__clkbuf_1 _09994_ (.A(_05141_),
    .X(_00242_));
 sky130_fd_sc_hd__mux2_1 _09995_ (.A0(net415),
    .A1(_04998_),
    .S(_05139_),
    .X(_05142_));
 sky130_fd_sc_hd__clkbuf_1 _09996_ (.A(_05142_),
    .X(_00243_));
 sky130_fd_sc_hd__mux2_1 _09997_ (.A0(net226),
    .A1(_05000_),
    .S(_05139_),
    .X(_05143_));
 sky130_fd_sc_hd__clkbuf_1 _09998_ (.A(_05143_),
    .X(_00244_));
 sky130_fd_sc_hd__mux2_1 _09999_ (.A0(net212),
    .A1(_05002_),
    .S(_05139_),
    .X(_05144_));
 sky130_fd_sc_hd__clkbuf_1 _10000_ (.A(_05144_),
    .X(_00245_));
 sky130_fd_sc_hd__mux2_1 _10001_ (.A0(net241),
    .A1(_05004_),
    .S(_05139_),
    .X(_05145_));
 sky130_fd_sc_hd__clkbuf_1 _10002_ (.A(_05145_),
    .X(_00246_));
 sky130_fd_sc_hd__mux2_1 _10003_ (.A0(net709),
    .A1(_05006_),
    .S(_05139_),
    .X(_05146_));
 sky130_fd_sc_hd__clkbuf_1 _10004_ (.A(_05146_),
    .X(_00247_));
 sky130_fd_sc_hd__mux2_1 _10005_ (.A0(net270),
    .A1(_05008_),
    .S(_05139_),
    .X(_05147_));
 sky130_fd_sc_hd__clkbuf_1 _10006_ (.A(_05147_),
    .X(_00248_));
 sky130_fd_sc_hd__mux2_1 _10007_ (.A0(net581),
    .A1(_05010_),
    .S(_05139_),
    .X(_05148_));
 sky130_fd_sc_hd__clkbuf_1 _10008_ (.A(_05148_),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_1 _10009_ (.A0(net489),
    .A1(_05012_),
    .S(_05139_),
    .X(_05149_));
 sky130_fd_sc_hd__clkbuf_1 _10010_ (.A(_05149_),
    .X(_00250_));
 sky130_fd_sc_hd__mux2_1 _10011_ (.A0(net392),
    .A1(_05014_),
    .S(_05138_),
    .X(_05150_));
 sky130_fd_sc_hd__clkbuf_1 _10012_ (.A(_05150_),
    .X(_00251_));
 sky130_fd_sc_hd__mux2_1 _10013_ (.A0(net170),
    .A1(_05016_),
    .S(_05138_),
    .X(_05151_));
 sky130_fd_sc_hd__clkbuf_1 _10014_ (.A(_05151_),
    .X(_00252_));
 sky130_fd_sc_hd__mux2_1 _10015_ (.A0(net309),
    .A1(_05018_),
    .S(_05138_),
    .X(_05152_));
 sky130_fd_sc_hd__clkbuf_1 _10016_ (.A(_05152_),
    .X(_00253_));
 sky130_fd_sc_hd__mux2_1 _10017_ (.A0(net613),
    .A1(_05020_),
    .S(_05138_),
    .X(_05153_));
 sky130_fd_sc_hd__clkbuf_1 _10018_ (.A(_05153_),
    .X(_00254_));
 sky130_fd_sc_hd__mux2_1 _10019_ (.A0(net54),
    .A1(_05022_),
    .S(_05138_),
    .X(_05154_));
 sky130_fd_sc_hd__clkbuf_1 _10020_ (.A(_05154_),
    .X(_00255_));
 sky130_fd_sc_hd__mux2_1 _10021_ (.A0(net725),
    .A1(_05024_),
    .S(_05138_),
    .X(_05155_));
 sky130_fd_sc_hd__clkbuf_1 _10022_ (.A(_05155_),
    .X(_00256_));
 sky130_fd_sc_hd__nor2_4 _10023_ (.A(_04076_),
    .B(_04501_),
    .Y(_05156_));
 sky130_fd_sc_hd__buf_4 _10024_ (.A(_05156_),
    .X(_05157_));
 sky130_fd_sc_hd__mux2_1 _10025_ (.A0(net363),
    .A1(_04992_),
    .S(_05157_),
    .X(_05158_));
 sky130_fd_sc_hd__clkbuf_1 _10026_ (.A(_05158_),
    .X(_00257_));
 sky130_fd_sc_hd__mux2_1 _10027_ (.A0(net371),
    .A1(_04996_),
    .S(_05157_),
    .X(_05159_));
 sky130_fd_sc_hd__clkbuf_1 _10028_ (.A(_05159_),
    .X(_00258_));
 sky130_fd_sc_hd__mux2_1 _10029_ (.A0(net1516),
    .A1(_04998_),
    .S(_05157_),
    .X(_05160_));
 sky130_fd_sc_hd__clkbuf_1 _10030_ (.A(_05160_),
    .X(_00259_));
 sky130_fd_sc_hd__mux2_1 _10031_ (.A0(net820),
    .A1(_05000_),
    .S(_05157_),
    .X(_05161_));
 sky130_fd_sc_hd__clkbuf_1 _10032_ (.A(_05161_),
    .X(_00260_));
 sky130_fd_sc_hd__mux2_1 _10033_ (.A0(net1019),
    .A1(_05002_),
    .S(_05157_),
    .X(_05162_));
 sky130_fd_sc_hd__clkbuf_1 _10034_ (.A(_05162_),
    .X(_00261_));
 sky130_fd_sc_hd__mux2_1 _10035_ (.A0(net320),
    .A1(_05004_),
    .S(_05157_),
    .X(_05163_));
 sky130_fd_sc_hd__clkbuf_1 _10036_ (.A(_05163_),
    .X(_00262_));
 sky130_fd_sc_hd__mux2_1 _10037_ (.A0(net261),
    .A1(_05006_),
    .S(_05157_),
    .X(_05164_));
 sky130_fd_sc_hd__clkbuf_1 _10038_ (.A(_05164_),
    .X(_00263_));
 sky130_fd_sc_hd__mux2_1 _10039_ (.A0(net714),
    .A1(_05008_),
    .S(_05157_),
    .X(_05165_));
 sky130_fd_sc_hd__clkbuf_1 _10040_ (.A(_05165_),
    .X(_00264_));
 sky130_fd_sc_hd__mux2_1 _10041_ (.A0(net125),
    .A1(_05010_),
    .S(_05157_),
    .X(_05166_));
 sky130_fd_sc_hd__clkbuf_1 _10042_ (.A(_05166_),
    .X(_00265_));
 sky130_fd_sc_hd__mux2_1 _10043_ (.A0(net454),
    .A1(_05012_),
    .S(_05157_),
    .X(_05167_));
 sky130_fd_sc_hd__clkbuf_1 _10044_ (.A(_05167_),
    .X(_00266_));
 sky130_fd_sc_hd__mux2_1 _10045_ (.A0(net200),
    .A1(_05014_),
    .S(_05156_),
    .X(_05168_));
 sky130_fd_sc_hd__clkbuf_1 _10046_ (.A(_05168_),
    .X(_00267_));
 sky130_fd_sc_hd__mux2_1 _10047_ (.A0(net298),
    .A1(_05016_),
    .S(_05156_),
    .X(_05169_));
 sky130_fd_sc_hd__clkbuf_1 _10048_ (.A(_05169_),
    .X(_00268_));
 sky130_fd_sc_hd__mux2_1 _10049_ (.A0(net326),
    .A1(_05018_),
    .S(_05156_),
    .X(_05170_));
 sky130_fd_sc_hd__clkbuf_1 _10050_ (.A(_05170_),
    .X(_00269_));
 sky130_fd_sc_hd__mux2_1 _10051_ (.A0(net96),
    .A1(_05020_),
    .S(_05156_),
    .X(_05171_));
 sky130_fd_sc_hd__clkbuf_1 _10052_ (.A(_05171_),
    .X(_00270_));
 sky130_fd_sc_hd__mux2_1 _10053_ (.A0(net404),
    .A1(_05022_),
    .S(_05156_),
    .X(_05172_));
 sky130_fd_sc_hd__clkbuf_1 _10054_ (.A(_05172_),
    .X(_00271_));
 sky130_fd_sc_hd__mux2_1 _10055_ (.A0(net362),
    .A1(_05024_),
    .S(_05156_),
    .X(_05173_));
 sky130_fd_sc_hd__clkbuf_1 _10056_ (.A(_05173_),
    .X(_00272_));
 sky130_fd_sc_hd__or2_1 _10057_ (.A(_04076_),
    .B(_04225_),
    .X(_05174_));
 sky130_fd_sc_hd__clkbuf_4 _10058_ (.A(_05174_),
    .X(_05175_));
 sky130_fd_sc_hd__buf_4 _10059_ (.A(_05175_),
    .X(_05176_));
 sky130_fd_sc_hd__mux2_1 _10060_ (.A0(_04406_),
    .A1(net1764),
    .S(_05176_),
    .X(_05177_));
 sky130_fd_sc_hd__clkbuf_1 _10061_ (.A(_05177_),
    .X(_00273_));
 sky130_fd_sc_hd__mux2_1 _10062_ (.A0(_04412_),
    .A1(net1289),
    .S(_05176_),
    .X(_05178_));
 sky130_fd_sc_hd__clkbuf_1 _10063_ (.A(_05178_),
    .X(_00274_));
 sky130_fd_sc_hd__mux2_1 _10064_ (.A0(_04414_),
    .A1(net726),
    .S(_05176_),
    .X(_05179_));
 sky130_fd_sc_hd__clkbuf_1 _10065_ (.A(_05179_),
    .X(_00275_));
 sky130_fd_sc_hd__mux2_1 _10066_ (.A0(_04416_),
    .A1(net1296),
    .S(_05176_),
    .X(_05180_));
 sky130_fd_sc_hd__clkbuf_1 _10067_ (.A(_05180_),
    .X(_00276_));
 sky130_fd_sc_hd__mux2_1 _10068_ (.A0(_04418_),
    .A1(net738),
    .S(_05176_),
    .X(_05181_));
 sky130_fd_sc_hd__clkbuf_1 _10069_ (.A(_05181_),
    .X(_00277_));
 sky130_fd_sc_hd__mux2_1 _10070_ (.A0(_04420_),
    .A1(net2047),
    .S(_05176_),
    .X(_05182_));
 sky130_fd_sc_hd__clkbuf_1 _10071_ (.A(_05182_),
    .X(_00278_));
 sky130_fd_sc_hd__mux2_1 _10072_ (.A0(_04422_),
    .A1(net1514),
    .S(_05176_),
    .X(_05183_));
 sky130_fd_sc_hd__clkbuf_1 _10073_ (.A(_05183_),
    .X(_00279_));
 sky130_fd_sc_hd__mux2_1 _10074_ (.A0(_04424_),
    .A1(net1042),
    .S(_05176_),
    .X(_05184_));
 sky130_fd_sc_hd__clkbuf_1 _10075_ (.A(_05184_),
    .X(_00280_));
 sky130_fd_sc_hd__mux2_1 _10076_ (.A0(_04426_),
    .A1(net1923),
    .S(_05176_),
    .X(_05185_));
 sky130_fd_sc_hd__clkbuf_1 _10077_ (.A(_05185_),
    .X(_00281_));
 sky130_fd_sc_hd__mux2_1 _10078_ (.A0(_04428_),
    .A1(net927),
    .S(_05176_),
    .X(_05186_));
 sky130_fd_sc_hd__clkbuf_1 _10079_ (.A(_05186_),
    .X(_00282_));
 sky130_fd_sc_hd__mux2_1 _10080_ (.A0(_04430_),
    .A1(net982),
    .S(_05175_),
    .X(_05187_));
 sky130_fd_sc_hd__clkbuf_1 _10081_ (.A(_05187_),
    .X(_00283_));
 sky130_fd_sc_hd__mux2_1 _10082_ (.A0(_04432_),
    .A1(net1148),
    .S(_05175_),
    .X(_05188_));
 sky130_fd_sc_hd__clkbuf_1 _10083_ (.A(_05188_),
    .X(_00284_));
 sky130_fd_sc_hd__mux2_1 _10084_ (.A0(_04434_),
    .A1(net1547),
    .S(_05175_),
    .X(_05189_));
 sky130_fd_sc_hd__clkbuf_1 _10085_ (.A(_05189_),
    .X(_00285_));
 sky130_fd_sc_hd__mux2_1 _10086_ (.A0(_04436_),
    .A1(net772),
    .S(_05175_),
    .X(_05190_));
 sky130_fd_sc_hd__clkbuf_1 _10087_ (.A(_05190_),
    .X(_00286_));
 sky130_fd_sc_hd__mux2_1 _10088_ (.A0(_04438_),
    .A1(net1970),
    .S(_05175_),
    .X(_05191_));
 sky130_fd_sc_hd__clkbuf_1 _10089_ (.A(_05191_),
    .X(_00287_));
 sky130_fd_sc_hd__mux2_1 _10090_ (.A0(_04440_),
    .A1(net580),
    .S(_05175_),
    .X(_05192_));
 sky130_fd_sc_hd__clkbuf_1 _10091_ (.A(_05192_),
    .X(_00288_));
 sky130_fd_sc_hd__nor2_4 _10092_ (.A(_04076_),
    .B(_04569_),
    .Y(_05193_));
 sky130_fd_sc_hd__buf_4 _10093_ (.A(_05193_),
    .X(_05194_));
 sky130_fd_sc_hd__mux2_1 _10094_ (.A0(net1124),
    .A1(_04992_),
    .S(_05194_),
    .X(_05195_));
 sky130_fd_sc_hd__clkbuf_1 _10095_ (.A(_05195_),
    .X(_00289_));
 sky130_fd_sc_hd__mux2_1 _10096_ (.A0(net89),
    .A1(_04996_),
    .S(_05194_),
    .X(_05196_));
 sky130_fd_sc_hd__clkbuf_1 _10097_ (.A(_05196_),
    .X(_00290_));
 sky130_fd_sc_hd__mux2_1 _10098_ (.A0(net990),
    .A1(_04998_),
    .S(_05194_),
    .X(_05197_));
 sky130_fd_sc_hd__clkbuf_1 _10099_ (.A(_05197_),
    .X(_00291_));
 sky130_fd_sc_hd__mux2_1 _10100_ (.A0(net459),
    .A1(_05000_),
    .S(_05194_),
    .X(_05198_));
 sky130_fd_sc_hd__clkbuf_1 _10101_ (.A(_05198_),
    .X(_00292_));
 sky130_fd_sc_hd__mux2_1 _10102_ (.A0(net462),
    .A1(_05002_),
    .S(_05194_),
    .X(_05199_));
 sky130_fd_sc_hd__clkbuf_1 _10103_ (.A(_05199_),
    .X(_00293_));
 sky130_fd_sc_hd__mux2_1 _10104_ (.A0(net819),
    .A1(_05004_),
    .S(_05194_),
    .X(_05200_));
 sky130_fd_sc_hd__clkbuf_1 _10105_ (.A(_05200_),
    .X(_00294_));
 sky130_fd_sc_hd__mux2_1 _10106_ (.A0(net747),
    .A1(_05006_),
    .S(_05194_),
    .X(_05201_));
 sky130_fd_sc_hd__clkbuf_1 _10107_ (.A(_05201_),
    .X(_00295_));
 sky130_fd_sc_hd__mux2_1 _10108_ (.A0(net604),
    .A1(_05008_),
    .S(_05194_),
    .X(_05202_));
 sky130_fd_sc_hd__clkbuf_1 _10109_ (.A(_05202_),
    .X(_00296_));
 sky130_fd_sc_hd__mux2_1 _10110_ (.A0(net352),
    .A1(_05010_),
    .S(_05194_),
    .X(_05203_));
 sky130_fd_sc_hd__clkbuf_1 _10111_ (.A(_05203_),
    .X(_00297_));
 sky130_fd_sc_hd__mux2_1 _10112_ (.A0(net748),
    .A1(_05012_),
    .S(_05194_),
    .X(_05204_));
 sky130_fd_sc_hd__clkbuf_1 _10113_ (.A(_05204_),
    .X(_00298_));
 sky130_fd_sc_hd__mux2_1 _10114_ (.A0(net1765),
    .A1(_05014_),
    .S(_05193_),
    .X(_05205_));
 sky130_fd_sc_hd__clkbuf_1 _10115_ (.A(_05205_),
    .X(_00299_));
 sky130_fd_sc_hd__mux2_1 _10116_ (.A0(net172),
    .A1(_05016_),
    .S(_05193_),
    .X(_05206_));
 sky130_fd_sc_hd__clkbuf_1 _10117_ (.A(_05206_),
    .X(_00300_));
 sky130_fd_sc_hd__mux2_1 _10118_ (.A0(net756),
    .A1(_05018_),
    .S(_05193_),
    .X(_05207_));
 sky130_fd_sc_hd__clkbuf_1 _10119_ (.A(_05207_),
    .X(_00301_));
 sky130_fd_sc_hd__mux2_1 _10120_ (.A0(net411),
    .A1(_05020_),
    .S(_05193_),
    .X(_05208_));
 sky130_fd_sc_hd__clkbuf_1 _10121_ (.A(_05208_),
    .X(_00302_));
 sky130_fd_sc_hd__mux2_1 _10122_ (.A0(net339),
    .A1(_05022_),
    .S(_05193_),
    .X(_05209_));
 sky130_fd_sc_hd__clkbuf_1 _10123_ (.A(_05209_),
    .X(_00303_));
 sky130_fd_sc_hd__mux2_1 _10124_ (.A0(net347),
    .A1(_05024_),
    .S(_05193_),
    .X(_05210_));
 sky130_fd_sc_hd__clkbuf_1 _10125_ (.A(_05210_),
    .X(_00304_));
 sky130_fd_sc_hd__buf_6 _10126_ (.A(_04069_),
    .X(_05211_));
 sky130_fd_sc_hd__or2_1 _10127_ (.A(_04076_),
    .B(_04184_),
    .X(_05212_));
 sky130_fd_sc_hd__clkbuf_4 _10128_ (.A(_05212_),
    .X(_05213_));
 sky130_fd_sc_hd__buf_4 _10129_ (.A(_05213_),
    .X(_05214_));
 sky130_fd_sc_hd__mux2_1 _10130_ (.A0(_05211_),
    .A1(net843),
    .S(_05214_),
    .X(_05215_));
 sky130_fd_sc_hd__clkbuf_1 _10131_ (.A(_05215_),
    .X(_00305_));
 sky130_fd_sc_hd__buf_4 _10132_ (.A(_04080_),
    .X(_05216_));
 sky130_fd_sc_hd__mux2_1 _10133_ (.A0(_05216_),
    .A1(net957),
    .S(_05214_),
    .X(_05217_));
 sky130_fd_sc_hd__clkbuf_1 _10134_ (.A(_05217_),
    .X(_00306_));
 sky130_fd_sc_hd__buf_6 _10135_ (.A(_04083_),
    .X(_05218_));
 sky130_fd_sc_hd__mux2_1 _10136_ (.A0(_05218_),
    .A1(net941),
    .S(_05214_),
    .X(_05219_));
 sky130_fd_sc_hd__clkbuf_1 _10137_ (.A(_05219_),
    .X(_00307_));
 sky130_fd_sc_hd__buf_6 _10138_ (.A(_04086_),
    .X(_05220_));
 sky130_fd_sc_hd__mux2_1 _10139_ (.A0(_05220_),
    .A1(net765),
    .S(_05214_),
    .X(_05221_));
 sky130_fd_sc_hd__clkbuf_1 _10140_ (.A(_05221_),
    .X(_00308_));
 sky130_fd_sc_hd__buf_6 _10141_ (.A(_04089_),
    .X(_05222_));
 sky130_fd_sc_hd__mux2_1 _10142_ (.A0(_05222_),
    .A1(net1154),
    .S(_05214_),
    .X(_05223_));
 sky130_fd_sc_hd__clkbuf_1 _10143_ (.A(_05223_),
    .X(_00309_));
 sky130_fd_sc_hd__buf_4 _10144_ (.A(_04092_),
    .X(_05224_));
 sky130_fd_sc_hd__mux2_1 _10145_ (.A0(_05224_),
    .A1(net548),
    .S(_05214_),
    .X(_05225_));
 sky130_fd_sc_hd__clkbuf_1 _10146_ (.A(_05225_),
    .X(_00310_));
 sky130_fd_sc_hd__clkbuf_8 _10147_ (.A(_04095_),
    .X(_05226_));
 sky130_fd_sc_hd__mux2_1 _10148_ (.A0(_05226_),
    .A1(net745),
    .S(_05214_),
    .X(_05227_));
 sky130_fd_sc_hd__clkbuf_1 _10149_ (.A(_05227_),
    .X(_00311_));
 sky130_fd_sc_hd__buf_6 _10150_ (.A(_04098_),
    .X(_05228_));
 sky130_fd_sc_hd__mux2_1 _10151_ (.A0(_05228_),
    .A1(net403),
    .S(_05214_),
    .X(_05229_));
 sky130_fd_sc_hd__clkbuf_1 _10152_ (.A(_05229_),
    .X(_00312_));
 sky130_fd_sc_hd__buf_6 _10153_ (.A(_04101_),
    .X(_05230_));
 sky130_fd_sc_hd__mux2_1 _10154_ (.A0(_05230_),
    .A1(net691),
    .S(_05214_),
    .X(_05231_));
 sky130_fd_sc_hd__clkbuf_1 _10155_ (.A(_05231_),
    .X(_00313_));
 sky130_fd_sc_hd__buf_6 _10156_ (.A(_04104_),
    .X(_05232_));
 sky130_fd_sc_hd__mux2_1 _10157_ (.A0(_05232_),
    .A1(net610),
    .S(_05214_),
    .X(_05233_));
 sky130_fd_sc_hd__clkbuf_1 _10158_ (.A(_05233_),
    .X(_00314_));
 sky130_fd_sc_hd__buf_4 _10159_ (.A(_04107_),
    .X(_05234_));
 sky130_fd_sc_hd__mux2_1 _10160_ (.A0(_05234_),
    .A1(net1482),
    .S(_05213_),
    .X(_05235_));
 sky130_fd_sc_hd__clkbuf_1 _10161_ (.A(_05235_),
    .X(_00315_));
 sky130_fd_sc_hd__buf_4 _10162_ (.A(_04110_),
    .X(_05236_));
 sky130_fd_sc_hd__mux2_1 _10163_ (.A0(_05236_),
    .A1(net804),
    .S(_05213_),
    .X(_05237_));
 sky130_fd_sc_hd__clkbuf_1 _10164_ (.A(_05237_),
    .X(_00316_));
 sky130_fd_sc_hd__buf_4 _10165_ (.A(_04113_),
    .X(_05238_));
 sky130_fd_sc_hd__mux2_1 _10166_ (.A0(_05238_),
    .A1(net1041),
    .S(_05213_),
    .X(_05239_));
 sky130_fd_sc_hd__clkbuf_1 _10167_ (.A(_05239_),
    .X(_00317_));
 sky130_fd_sc_hd__buf_4 _10168_ (.A(_04116_),
    .X(_05240_));
 sky130_fd_sc_hd__mux2_1 _10169_ (.A0(_05240_),
    .A1(net1276),
    .S(_05213_),
    .X(_05241_));
 sky130_fd_sc_hd__clkbuf_1 _10170_ (.A(_05241_),
    .X(_00318_));
 sky130_fd_sc_hd__buf_4 _10171_ (.A(_04119_),
    .X(_05242_));
 sky130_fd_sc_hd__mux2_1 _10172_ (.A0(_05242_),
    .A1(net1465),
    .S(_05213_),
    .X(_05243_));
 sky130_fd_sc_hd__clkbuf_1 _10173_ (.A(_05243_),
    .X(_00319_));
 sky130_fd_sc_hd__buf_4 _10174_ (.A(_04122_),
    .X(_05244_));
 sky130_fd_sc_hd__mux2_1 _10175_ (.A0(_05244_),
    .A1(net1709),
    .S(_05213_),
    .X(_05245_));
 sky130_fd_sc_hd__clkbuf_1 _10176_ (.A(_05245_),
    .X(_00320_));
 sky130_fd_sc_hd__or2_1 _10177_ (.A(_04076_),
    .B(_04607_),
    .X(_05246_));
 sky130_fd_sc_hd__clkbuf_4 _10178_ (.A(_05246_),
    .X(_05247_));
 sky130_fd_sc_hd__buf_4 _10179_ (.A(_05247_),
    .X(_05248_));
 sky130_fd_sc_hd__mux2_1 _10180_ (.A0(_05211_),
    .A1(net974),
    .S(_05248_),
    .X(_05249_));
 sky130_fd_sc_hd__clkbuf_1 _10181_ (.A(_05249_),
    .X(_00321_));
 sky130_fd_sc_hd__mux2_1 _10182_ (.A0(_05216_),
    .A1(net1559),
    .S(_05248_),
    .X(_05250_));
 sky130_fd_sc_hd__clkbuf_1 _10183_ (.A(_05250_),
    .X(_00322_));
 sky130_fd_sc_hd__mux2_1 _10184_ (.A0(_05218_),
    .A1(net559),
    .S(_05248_),
    .X(_05251_));
 sky130_fd_sc_hd__clkbuf_1 _10185_ (.A(_05251_),
    .X(_00323_));
 sky130_fd_sc_hd__mux2_1 _10186_ (.A0(_05220_),
    .A1(net883),
    .S(_05248_),
    .X(_05252_));
 sky130_fd_sc_hd__clkbuf_1 _10187_ (.A(_05252_),
    .X(_00324_));
 sky130_fd_sc_hd__mux2_1 _10188_ (.A0(_05222_),
    .A1(net1770),
    .S(_05248_),
    .X(_05253_));
 sky130_fd_sc_hd__clkbuf_1 _10189_ (.A(_05253_),
    .X(_00325_));
 sky130_fd_sc_hd__mux2_1 _10190_ (.A0(_05224_),
    .A1(net1123),
    .S(_05248_),
    .X(_05254_));
 sky130_fd_sc_hd__clkbuf_1 _10191_ (.A(_05254_),
    .X(_00326_));
 sky130_fd_sc_hd__mux2_1 _10192_ (.A0(_05226_),
    .A1(net538),
    .S(_05248_),
    .X(_05255_));
 sky130_fd_sc_hd__clkbuf_1 _10193_ (.A(_05255_),
    .X(_00327_));
 sky130_fd_sc_hd__mux2_1 _10194_ (.A0(_05228_),
    .A1(net1810),
    .S(_05248_),
    .X(_05256_));
 sky130_fd_sc_hd__clkbuf_1 _10195_ (.A(_05256_),
    .X(_00328_));
 sky130_fd_sc_hd__mux2_1 _10196_ (.A0(_05230_),
    .A1(net1825),
    .S(_05248_),
    .X(_05257_));
 sky130_fd_sc_hd__clkbuf_1 _10197_ (.A(_05257_),
    .X(_00329_));
 sky130_fd_sc_hd__mux2_1 _10198_ (.A0(_05232_),
    .A1(net1789),
    .S(_05248_),
    .X(_05258_));
 sky130_fd_sc_hd__clkbuf_1 _10199_ (.A(_05258_),
    .X(_00330_));
 sky130_fd_sc_hd__mux2_1 _10200_ (.A0(_05234_),
    .A1(net1002),
    .S(_05247_),
    .X(_05259_));
 sky130_fd_sc_hd__clkbuf_1 _10201_ (.A(_05259_),
    .X(_00331_));
 sky130_fd_sc_hd__mux2_1 _10202_ (.A0(_05236_),
    .A1(net1139),
    .S(_05247_),
    .X(_05260_));
 sky130_fd_sc_hd__clkbuf_1 _10203_ (.A(_05260_),
    .X(_00332_));
 sky130_fd_sc_hd__mux2_1 _10204_ (.A0(_05238_),
    .A1(net876),
    .S(_05247_),
    .X(_05261_));
 sky130_fd_sc_hd__clkbuf_1 _10205_ (.A(_05261_),
    .X(_00333_));
 sky130_fd_sc_hd__mux2_1 _10206_ (.A0(_05240_),
    .A1(net1883),
    .S(_05247_),
    .X(_05262_));
 sky130_fd_sc_hd__clkbuf_1 _10207_ (.A(_05262_),
    .X(_00334_));
 sky130_fd_sc_hd__mux2_1 _10208_ (.A0(_05242_),
    .A1(net1171),
    .S(_05247_),
    .X(_05263_));
 sky130_fd_sc_hd__clkbuf_1 _10209_ (.A(_05263_),
    .X(_00335_));
 sky130_fd_sc_hd__mux2_1 _10210_ (.A0(_05244_),
    .A1(net1672),
    .S(_05247_),
    .X(_05264_));
 sky130_fd_sc_hd__clkbuf_1 _10211_ (.A(_05264_),
    .X(_00336_));
 sky130_fd_sc_hd__or3_1 _10212_ (.A(_02702_),
    .B(_05026_),
    .C(_04075_),
    .X(_05265_));
 sky130_fd_sc_hd__clkbuf_4 _10213_ (.A(_05265_),
    .X(_05266_));
 sky130_fd_sc_hd__buf_4 _10214_ (.A(_05266_),
    .X(_05267_));
 sky130_fd_sc_hd__mux2_1 _10215_ (.A0(_05211_),
    .A1(net1005),
    .S(_05267_),
    .X(_05268_));
 sky130_fd_sc_hd__clkbuf_1 _10216_ (.A(_05268_),
    .X(_00337_));
 sky130_fd_sc_hd__mux2_1 _10217_ (.A0(_05216_),
    .A1(net1627),
    .S(_05267_),
    .X(_05269_));
 sky130_fd_sc_hd__clkbuf_1 _10218_ (.A(_05269_),
    .X(_00338_));
 sky130_fd_sc_hd__mux2_1 _10219_ (.A0(_05218_),
    .A1(net1792),
    .S(_05267_),
    .X(_05270_));
 sky130_fd_sc_hd__clkbuf_1 _10220_ (.A(_05270_),
    .X(_00339_));
 sky130_fd_sc_hd__mux2_1 _10221_ (.A0(_05220_),
    .A1(net1739),
    .S(_05267_),
    .X(_05271_));
 sky130_fd_sc_hd__clkbuf_1 _10222_ (.A(_05271_),
    .X(_00340_));
 sky130_fd_sc_hd__mux2_1 _10223_ (.A0(_05222_),
    .A1(net1485),
    .S(_05267_),
    .X(_05272_));
 sky130_fd_sc_hd__clkbuf_1 _10224_ (.A(_05272_),
    .X(_00341_));
 sky130_fd_sc_hd__mux2_1 _10225_ (.A0(_05224_),
    .A1(net717),
    .S(_05267_),
    .X(_05273_));
 sky130_fd_sc_hd__clkbuf_1 _10226_ (.A(_05273_),
    .X(_00342_));
 sky130_fd_sc_hd__mux2_1 _10227_ (.A0(_05226_),
    .A1(net1748),
    .S(_05267_),
    .X(_05274_));
 sky130_fd_sc_hd__clkbuf_1 _10228_ (.A(_05274_),
    .X(_00343_));
 sky130_fd_sc_hd__mux2_1 _10229_ (.A0(_05228_),
    .A1(net1239),
    .S(_05267_),
    .X(_05275_));
 sky130_fd_sc_hd__clkbuf_1 _10230_ (.A(_05275_),
    .X(_00344_));
 sky130_fd_sc_hd__mux2_1 _10231_ (.A0(_05230_),
    .A1(net330),
    .S(_05267_),
    .X(_05276_));
 sky130_fd_sc_hd__clkbuf_1 _10232_ (.A(_05276_),
    .X(_00345_));
 sky130_fd_sc_hd__mux2_1 _10233_ (.A0(_05232_),
    .A1(net475),
    .S(_05267_),
    .X(_05277_));
 sky130_fd_sc_hd__clkbuf_1 _10234_ (.A(_05277_),
    .X(_00346_));
 sky130_fd_sc_hd__mux2_1 _10235_ (.A0(_05234_),
    .A1(net942),
    .S(_05266_),
    .X(_05278_));
 sky130_fd_sc_hd__clkbuf_1 _10236_ (.A(_05278_),
    .X(_00347_));
 sky130_fd_sc_hd__mux2_1 _10237_ (.A0(_05236_),
    .A1(net1907),
    .S(_05266_),
    .X(_05279_));
 sky130_fd_sc_hd__clkbuf_1 _10238_ (.A(_05279_),
    .X(_00348_));
 sky130_fd_sc_hd__mux2_1 _10239_ (.A0(_05238_),
    .A1(net1848),
    .S(_05266_),
    .X(_05280_));
 sky130_fd_sc_hd__clkbuf_1 _10240_ (.A(_05280_),
    .X(_00349_));
 sky130_fd_sc_hd__mux2_1 _10241_ (.A0(_05240_),
    .A1(net544),
    .S(_05266_),
    .X(_05281_));
 sky130_fd_sc_hd__clkbuf_1 _10242_ (.A(_05281_),
    .X(_00350_));
 sky130_fd_sc_hd__mux2_1 _10243_ (.A0(_05242_),
    .A1(net1651),
    .S(_05266_),
    .X(_05282_));
 sky130_fd_sc_hd__clkbuf_1 _10244_ (.A(_05282_),
    .X(_00351_));
 sky130_fd_sc_hd__mux2_1 _10245_ (.A0(_05244_),
    .A1(net1708),
    .S(_05266_),
    .X(_05283_));
 sky130_fd_sc_hd__clkbuf_1 _10246_ (.A(_05283_),
    .X(_00352_));
 sky130_fd_sc_hd__nor2_4 _10247_ (.A(_04076_),
    .B(_04646_),
    .Y(_05284_));
 sky130_fd_sc_hd__buf_4 _10248_ (.A(_05284_),
    .X(_05285_));
 sky130_fd_sc_hd__mux2_1 _10249_ (.A0(net1038),
    .A1(_04992_),
    .S(_05285_),
    .X(_05286_));
 sky130_fd_sc_hd__clkbuf_1 _10250_ (.A(_05286_),
    .X(_00353_));
 sky130_fd_sc_hd__mux2_1 _10251_ (.A0(net711),
    .A1(_04996_),
    .S(_05285_),
    .X(_05287_));
 sky130_fd_sc_hd__clkbuf_1 _10252_ (.A(_05287_),
    .X(_00354_));
 sky130_fd_sc_hd__mux2_1 _10253_ (.A0(net342),
    .A1(_04998_),
    .S(_05285_),
    .X(_05288_));
 sky130_fd_sc_hd__clkbuf_1 _10254_ (.A(_05288_),
    .X(_00355_));
 sky130_fd_sc_hd__mux2_1 _10255_ (.A0(net1699),
    .A1(_05000_),
    .S(_05285_),
    .X(_05289_));
 sky130_fd_sc_hd__clkbuf_1 _10256_ (.A(_05289_),
    .X(_00356_));
 sky130_fd_sc_hd__mux2_1 _10257_ (.A0(net835),
    .A1(_05002_),
    .S(_05285_),
    .X(_05290_));
 sky130_fd_sc_hd__clkbuf_1 _10258_ (.A(_05290_),
    .X(_00357_));
 sky130_fd_sc_hd__mux2_1 _10259_ (.A0(net1165),
    .A1(_05004_),
    .S(_05285_),
    .X(_05291_));
 sky130_fd_sc_hd__clkbuf_1 _10260_ (.A(_05291_),
    .X(_00358_));
 sky130_fd_sc_hd__mux2_1 _10261_ (.A0(net606),
    .A1(_05006_),
    .S(_05285_),
    .X(_05292_));
 sky130_fd_sc_hd__clkbuf_1 _10262_ (.A(_05292_),
    .X(_00359_));
 sky130_fd_sc_hd__mux2_1 _10263_ (.A0(net151),
    .A1(_05008_),
    .S(_05285_),
    .X(_05293_));
 sky130_fd_sc_hd__clkbuf_1 _10264_ (.A(_05293_),
    .X(_00360_));
 sky130_fd_sc_hd__mux2_1 _10265_ (.A0(net811),
    .A1(_05010_),
    .S(_05285_),
    .X(_05294_));
 sky130_fd_sc_hd__clkbuf_1 _10266_ (.A(_05294_),
    .X(_00361_));
 sky130_fd_sc_hd__mux2_1 _10267_ (.A0(net504),
    .A1(_05012_),
    .S(_05285_),
    .X(_05295_));
 sky130_fd_sc_hd__clkbuf_1 _10268_ (.A(_05295_),
    .X(_00362_));
 sky130_fd_sc_hd__mux2_1 _10269_ (.A0(net349),
    .A1(_05014_),
    .S(_05284_),
    .X(_05296_));
 sky130_fd_sc_hd__clkbuf_1 _10270_ (.A(_05296_),
    .X(_00363_));
 sky130_fd_sc_hd__mux2_1 _10271_ (.A0(net258),
    .A1(_05016_),
    .S(_05284_),
    .X(_05297_));
 sky130_fd_sc_hd__clkbuf_1 _10272_ (.A(_05297_),
    .X(_00364_));
 sky130_fd_sc_hd__mux2_1 _10273_ (.A0(net288),
    .A1(_05018_),
    .S(_05284_),
    .X(_05298_));
 sky130_fd_sc_hd__clkbuf_1 _10274_ (.A(_05298_),
    .X(_00365_));
 sky130_fd_sc_hd__mux2_1 _10275_ (.A0(net163),
    .A1(_05020_),
    .S(_05284_),
    .X(_05299_));
 sky130_fd_sc_hd__clkbuf_1 _10276_ (.A(_05299_),
    .X(_00366_));
 sky130_fd_sc_hd__mux2_1 _10277_ (.A0(net618),
    .A1(_05022_),
    .S(_05284_),
    .X(_05300_));
 sky130_fd_sc_hd__clkbuf_1 _10278_ (.A(_05300_),
    .X(_00367_));
 sky130_fd_sc_hd__mux2_1 _10279_ (.A0(net1646),
    .A1(_05024_),
    .S(_05284_),
    .X(_05301_));
 sky130_fd_sc_hd__clkbuf_1 _10280_ (.A(_05301_),
    .X(_00368_));
 sky130_fd_sc_hd__or2_1 _10281_ (.A(_04076_),
    .B(_04127_),
    .X(_05302_));
 sky130_fd_sc_hd__clkbuf_4 _10282_ (.A(_05302_),
    .X(_05303_));
 sky130_fd_sc_hd__clkbuf_8 _10283_ (.A(_05303_),
    .X(_05304_));
 sky130_fd_sc_hd__mux2_1 _10284_ (.A0(_05211_),
    .A1(net1314),
    .S(_05304_),
    .X(_05305_));
 sky130_fd_sc_hd__clkbuf_1 _10285_ (.A(_05305_),
    .X(_00369_));
 sky130_fd_sc_hd__mux2_1 _10286_ (.A0(_05216_),
    .A1(net1361),
    .S(_05304_),
    .X(_05306_));
 sky130_fd_sc_hd__clkbuf_1 _10287_ (.A(_05306_),
    .X(_00370_));
 sky130_fd_sc_hd__mux2_1 _10288_ (.A0(_05218_),
    .A1(net892),
    .S(_05304_),
    .X(_05307_));
 sky130_fd_sc_hd__clkbuf_1 _10289_ (.A(_05307_),
    .X(_00371_));
 sky130_fd_sc_hd__mux2_1 _10290_ (.A0(_05220_),
    .A1(net859),
    .S(_05304_),
    .X(_05308_));
 sky130_fd_sc_hd__clkbuf_1 _10291_ (.A(_05308_),
    .X(_00372_));
 sky130_fd_sc_hd__mux2_1 _10292_ (.A0(_05222_),
    .A1(net862),
    .S(_05304_),
    .X(_05309_));
 sky130_fd_sc_hd__clkbuf_1 _10293_ (.A(_05309_),
    .X(_00373_));
 sky130_fd_sc_hd__mux2_1 _10294_ (.A0(_05224_),
    .A1(net973),
    .S(_05304_),
    .X(_05310_));
 sky130_fd_sc_hd__clkbuf_1 _10295_ (.A(_05310_),
    .X(_00374_));
 sky130_fd_sc_hd__mux2_1 _10296_ (.A0(_05226_),
    .A1(net689),
    .S(_05304_),
    .X(_05311_));
 sky130_fd_sc_hd__clkbuf_1 _10297_ (.A(_05311_),
    .X(_00375_));
 sky130_fd_sc_hd__mux2_1 _10298_ (.A0(_05228_),
    .A1(net858),
    .S(_05304_),
    .X(_05312_));
 sky130_fd_sc_hd__clkbuf_1 _10299_ (.A(_05312_),
    .X(_00376_));
 sky130_fd_sc_hd__mux2_1 _10300_ (.A0(_05230_),
    .A1(net911),
    .S(_05304_),
    .X(_05313_));
 sky130_fd_sc_hd__clkbuf_1 _10301_ (.A(_05313_),
    .X(_00377_));
 sky130_fd_sc_hd__mux2_1 _10302_ (.A0(_05232_),
    .A1(net1084),
    .S(_05304_),
    .X(_05314_));
 sky130_fd_sc_hd__clkbuf_1 _10303_ (.A(_05314_),
    .X(_00378_));
 sky130_fd_sc_hd__mux2_1 _10304_ (.A0(_05234_),
    .A1(net588),
    .S(_05303_),
    .X(_05315_));
 sky130_fd_sc_hd__clkbuf_1 _10305_ (.A(_05315_),
    .X(_00379_));
 sky130_fd_sc_hd__mux2_1 _10306_ (.A0(_05236_),
    .A1(net570),
    .S(_05303_),
    .X(_05316_));
 sky130_fd_sc_hd__clkbuf_1 _10307_ (.A(_05316_),
    .X(_00380_));
 sky130_fd_sc_hd__mux2_1 _10308_ (.A0(_05238_),
    .A1(net1141),
    .S(_05303_),
    .X(_05317_));
 sky130_fd_sc_hd__clkbuf_1 _10309_ (.A(_05317_),
    .X(_00381_));
 sky130_fd_sc_hd__mux2_1 _10310_ (.A0(_05240_),
    .A1(net978),
    .S(_05303_),
    .X(_05318_));
 sky130_fd_sc_hd__clkbuf_1 _10311_ (.A(_05318_),
    .X(_00382_));
 sky130_fd_sc_hd__mux2_1 _10312_ (.A0(_05242_),
    .A1(net1032),
    .S(_05303_),
    .X(_05319_));
 sky130_fd_sc_hd__clkbuf_1 _10313_ (.A(_05319_),
    .X(_00383_));
 sky130_fd_sc_hd__mux2_1 _10314_ (.A0(_05244_),
    .A1(net571),
    .S(_05303_),
    .X(_05320_));
 sky130_fd_sc_hd__clkbuf_1 _10315_ (.A(_05320_),
    .X(_00384_));
 sky130_fd_sc_hd__or2_1 _10316_ (.A(_04075_),
    .B(_04684_),
    .X(_05321_));
 sky130_fd_sc_hd__clkbuf_4 _10317_ (.A(_05321_),
    .X(_05322_));
 sky130_fd_sc_hd__buf_4 _10318_ (.A(_05322_),
    .X(_05323_));
 sky130_fd_sc_hd__mux2_1 _10319_ (.A0(_05211_),
    .A1(net1430),
    .S(_05323_),
    .X(_05324_));
 sky130_fd_sc_hd__clkbuf_1 _10320_ (.A(_05324_),
    .X(_00385_));
 sky130_fd_sc_hd__mux2_1 _10321_ (.A0(_05216_),
    .A1(net1056),
    .S(_05323_),
    .X(_05325_));
 sky130_fd_sc_hd__clkbuf_1 _10322_ (.A(_05325_),
    .X(_00386_));
 sky130_fd_sc_hd__mux2_1 _10323_ (.A0(_05218_),
    .A1(net1900),
    .S(_05323_),
    .X(_05326_));
 sky130_fd_sc_hd__clkbuf_1 _10324_ (.A(_05326_),
    .X(_00387_));
 sky130_fd_sc_hd__mux2_1 _10325_ (.A0(_05220_),
    .A1(net1500),
    .S(_05323_),
    .X(_05327_));
 sky130_fd_sc_hd__clkbuf_1 _10326_ (.A(_05327_),
    .X(_00388_));
 sky130_fd_sc_hd__mux2_1 _10327_ (.A0(_05222_),
    .A1(net1932),
    .S(_05323_),
    .X(_05328_));
 sky130_fd_sc_hd__clkbuf_1 _10328_ (.A(_05328_),
    .X(_00389_));
 sky130_fd_sc_hd__mux2_1 _10329_ (.A0(_05224_),
    .A1(net1884),
    .S(_05323_),
    .X(_05329_));
 sky130_fd_sc_hd__clkbuf_1 _10330_ (.A(_05329_),
    .X(_00390_));
 sky130_fd_sc_hd__mux2_1 _10331_ (.A0(_05226_),
    .A1(net1421),
    .S(_05323_),
    .X(_05330_));
 sky130_fd_sc_hd__clkbuf_1 _10332_ (.A(_05330_),
    .X(_00391_));
 sky130_fd_sc_hd__mux2_1 _10333_ (.A0(_05228_),
    .A1(net575),
    .S(_05323_),
    .X(_05331_));
 sky130_fd_sc_hd__clkbuf_1 _10334_ (.A(_05331_),
    .X(_00392_));
 sky130_fd_sc_hd__mux2_1 _10335_ (.A0(_05230_),
    .A1(net1947),
    .S(_05323_),
    .X(_05332_));
 sky130_fd_sc_hd__clkbuf_1 _10336_ (.A(_05332_),
    .X(_00393_));
 sky130_fd_sc_hd__mux2_1 _10337_ (.A0(_05232_),
    .A1(net1476),
    .S(_05323_),
    .X(_05333_));
 sky130_fd_sc_hd__clkbuf_1 _10338_ (.A(_05333_),
    .X(_00394_));
 sky130_fd_sc_hd__mux2_1 _10339_ (.A0(_05234_),
    .A1(net1467),
    .S(_05322_),
    .X(_05334_));
 sky130_fd_sc_hd__clkbuf_1 _10340_ (.A(_05334_),
    .X(_00395_));
 sky130_fd_sc_hd__mux2_1 _10341_ (.A0(_05236_),
    .A1(net634),
    .S(_05322_),
    .X(_05335_));
 sky130_fd_sc_hd__clkbuf_1 _10342_ (.A(_05335_),
    .X(_00396_));
 sky130_fd_sc_hd__mux2_1 _10343_ (.A0(_05238_),
    .A1(net696),
    .S(_05322_),
    .X(_05336_));
 sky130_fd_sc_hd__clkbuf_1 _10344_ (.A(_05336_),
    .X(_00397_));
 sky130_fd_sc_hd__mux2_1 _10345_ (.A0(_05240_),
    .A1(net1515),
    .S(_05322_),
    .X(_05337_));
 sky130_fd_sc_hd__clkbuf_1 _10346_ (.A(_05337_),
    .X(_00398_));
 sky130_fd_sc_hd__mux2_1 _10347_ (.A0(_05242_),
    .A1(net1486),
    .S(_05322_),
    .X(_05338_));
 sky130_fd_sc_hd__clkbuf_1 _10348_ (.A(_05338_),
    .X(_00399_));
 sky130_fd_sc_hd__mux2_1 _10349_ (.A0(_05244_),
    .A1(net1377),
    .S(_05322_),
    .X(_05339_));
 sky130_fd_sc_hd__clkbuf_1 _10350_ (.A(_05339_),
    .X(_00400_));
 sky130_fd_sc_hd__nor2_4 _10351_ (.A(_04184_),
    .B(_04368_),
    .Y(_05340_));
 sky130_fd_sc_hd__buf_4 _10352_ (.A(_05340_),
    .X(_05341_));
 sky130_fd_sc_hd__mux2_1 _10353_ (.A0(net2073),
    .A1(_04992_),
    .S(_05341_),
    .X(_05342_));
 sky130_fd_sc_hd__clkbuf_1 _10354_ (.A(_05342_),
    .X(_00401_));
 sky130_fd_sc_hd__mux2_1 _10355_ (.A0(net1450),
    .A1(_04996_),
    .S(_05341_),
    .X(_05343_));
 sky130_fd_sc_hd__clkbuf_1 _10356_ (.A(_05343_),
    .X(_00402_));
 sky130_fd_sc_hd__mux2_1 _10357_ (.A0(net1405),
    .A1(_04998_),
    .S(_05341_),
    .X(_05344_));
 sky130_fd_sc_hd__clkbuf_1 _10358_ (.A(_05344_),
    .X(_00403_));
 sky130_fd_sc_hd__mux2_1 _10359_ (.A0(net547),
    .A1(_05000_),
    .S(_05341_),
    .X(_05345_));
 sky130_fd_sc_hd__clkbuf_1 _10360_ (.A(_05345_),
    .X(_00404_));
 sky130_fd_sc_hd__mux2_1 _10361_ (.A0(net457),
    .A1(_05002_),
    .S(_05341_),
    .X(_05346_));
 sky130_fd_sc_hd__clkbuf_1 _10362_ (.A(_05346_),
    .X(_00405_));
 sky130_fd_sc_hd__mux2_1 _10363_ (.A0(net143),
    .A1(_05004_),
    .S(_05341_),
    .X(_05347_));
 sky130_fd_sc_hd__clkbuf_1 _10364_ (.A(_05347_),
    .X(_00406_));
 sky130_fd_sc_hd__mux2_1 _10365_ (.A0(net1023),
    .A1(_05006_),
    .S(_05341_),
    .X(_05348_));
 sky130_fd_sc_hd__clkbuf_1 _10366_ (.A(_05348_),
    .X(_00407_));
 sky130_fd_sc_hd__mux2_1 _10367_ (.A0(net1233),
    .A1(_05008_),
    .S(_05341_),
    .X(_05349_));
 sky130_fd_sc_hd__clkbuf_1 _10368_ (.A(_05349_),
    .X(_00408_));
 sky130_fd_sc_hd__mux2_1 _10369_ (.A0(net1135),
    .A1(_05010_),
    .S(_05341_),
    .X(_05350_));
 sky130_fd_sc_hd__clkbuf_1 _10370_ (.A(_05350_),
    .X(_00409_));
 sky130_fd_sc_hd__mux2_1 _10371_ (.A0(net650),
    .A1(_05012_),
    .S(_05341_),
    .X(_05351_));
 sky130_fd_sc_hd__clkbuf_1 _10372_ (.A(_05351_),
    .X(_00410_));
 sky130_fd_sc_hd__mux2_1 _10373_ (.A0(net1297),
    .A1(_05014_),
    .S(_05340_),
    .X(_05352_));
 sky130_fd_sc_hd__clkbuf_1 _10374_ (.A(_05352_),
    .X(_00411_));
 sky130_fd_sc_hd__mux2_1 _10375_ (.A0(net648),
    .A1(_05016_),
    .S(_05340_),
    .X(_05353_));
 sky130_fd_sc_hd__clkbuf_1 _10376_ (.A(_05353_),
    .X(_00412_));
 sky130_fd_sc_hd__mux2_1 _10377_ (.A0(net866),
    .A1(_05018_),
    .S(_05340_),
    .X(_05354_));
 sky130_fd_sc_hd__clkbuf_1 _10378_ (.A(_05354_),
    .X(_00413_));
 sky130_fd_sc_hd__mux2_1 _10379_ (.A0(net1101),
    .A1(_05020_),
    .S(_05340_),
    .X(_05355_));
 sky130_fd_sc_hd__clkbuf_1 _10380_ (.A(_05355_),
    .X(_00414_));
 sky130_fd_sc_hd__mux2_1 _10381_ (.A0(net997),
    .A1(_05022_),
    .S(_05340_),
    .X(_05356_));
 sky130_fd_sc_hd__clkbuf_1 _10382_ (.A(_05356_),
    .X(_00415_));
 sky130_fd_sc_hd__mux2_1 _10383_ (.A0(net341),
    .A1(_05024_),
    .S(_05340_),
    .X(_05357_));
 sky130_fd_sc_hd__clkbuf_1 _10384_ (.A(_05357_),
    .X(_00416_));
 sky130_fd_sc_hd__or2_1 _10385_ (.A(_04075_),
    .B(_04365_),
    .X(_05358_));
 sky130_fd_sc_hd__clkbuf_4 _10386_ (.A(_05358_),
    .X(_05359_));
 sky130_fd_sc_hd__buf_4 _10387_ (.A(_05359_),
    .X(_05360_));
 sky130_fd_sc_hd__mux2_1 _10388_ (.A0(_05211_),
    .A1(net1366),
    .S(_05360_),
    .X(_05361_));
 sky130_fd_sc_hd__clkbuf_1 _10389_ (.A(_05361_),
    .X(_00417_));
 sky130_fd_sc_hd__mux2_1 _10390_ (.A0(_05216_),
    .A1(net1222),
    .S(_05360_),
    .X(_05362_));
 sky130_fd_sc_hd__clkbuf_1 _10391_ (.A(_05362_),
    .X(_00418_));
 sky130_fd_sc_hd__mux2_1 _10392_ (.A0(_05218_),
    .A1(net1301),
    .S(_05360_),
    .X(_05363_));
 sky130_fd_sc_hd__clkbuf_1 _10393_ (.A(_05363_),
    .X(_00419_));
 sky130_fd_sc_hd__mux2_1 _10394_ (.A0(_05220_),
    .A1(net967),
    .S(_05360_),
    .X(_05364_));
 sky130_fd_sc_hd__clkbuf_1 _10395_ (.A(_05364_),
    .X(_00420_));
 sky130_fd_sc_hd__mux2_1 _10396_ (.A0(_05222_),
    .A1(net1073),
    .S(_05360_),
    .X(_05365_));
 sky130_fd_sc_hd__clkbuf_1 _10397_ (.A(_05365_),
    .X(_00421_));
 sky130_fd_sc_hd__mux2_1 _10398_ (.A0(_05224_),
    .A1(net1303),
    .S(_05360_),
    .X(_05366_));
 sky130_fd_sc_hd__clkbuf_1 _10399_ (.A(_05366_),
    .X(_00422_));
 sky130_fd_sc_hd__mux2_1 _10400_ (.A0(_05226_),
    .A1(net1586),
    .S(_05360_),
    .X(_05367_));
 sky130_fd_sc_hd__clkbuf_1 _10401_ (.A(_05367_),
    .X(_00423_));
 sky130_fd_sc_hd__mux2_1 _10402_ (.A0(_05228_),
    .A1(net1236),
    .S(_05360_),
    .X(_05368_));
 sky130_fd_sc_hd__clkbuf_1 _10403_ (.A(_05368_),
    .X(_00424_));
 sky130_fd_sc_hd__mux2_1 _10404_ (.A0(_05230_),
    .A1(net712),
    .S(_05360_),
    .X(_05369_));
 sky130_fd_sc_hd__clkbuf_1 _10405_ (.A(_05369_),
    .X(_00425_));
 sky130_fd_sc_hd__mux2_1 _10406_ (.A0(_05232_),
    .A1(net1656),
    .S(_05360_),
    .X(_05370_));
 sky130_fd_sc_hd__clkbuf_1 _10407_ (.A(_05370_),
    .X(_00426_));
 sky130_fd_sc_hd__mux2_1 _10408_ (.A0(_05234_),
    .A1(net742),
    .S(_05359_),
    .X(_05371_));
 sky130_fd_sc_hd__clkbuf_1 _10409_ (.A(_05371_),
    .X(_00427_));
 sky130_fd_sc_hd__mux2_1 _10410_ (.A0(_05236_),
    .A1(net1394),
    .S(_05359_),
    .X(_05372_));
 sky130_fd_sc_hd__clkbuf_1 _10411_ (.A(_05372_),
    .X(_00428_));
 sky130_fd_sc_hd__mux2_1 _10412_ (.A0(_05238_),
    .A1(net609),
    .S(_05359_),
    .X(_05373_));
 sky130_fd_sc_hd__clkbuf_1 _10413_ (.A(_05373_),
    .X(_00429_));
 sky130_fd_sc_hd__mux2_1 _10414_ (.A0(_05240_),
    .A1(net1489),
    .S(_05359_),
    .X(_05374_));
 sky130_fd_sc_hd__clkbuf_1 _10415_ (.A(_05374_),
    .X(_00430_));
 sky130_fd_sc_hd__mux2_1 _10416_ (.A0(_05242_),
    .A1(net1402),
    .S(_05359_),
    .X(_05375_));
 sky130_fd_sc_hd__clkbuf_1 _10417_ (.A(_05375_),
    .X(_00431_));
 sky130_fd_sc_hd__mux2_1 _10418_ (.A0(_05244_),
    .A1(net1176),
    .S(_05359_),
    .X(_05376_));
 sky130_fd_sc_hd__clkbuf_1 _10419_ (.A(_05376_),
    .X(_00432_));
 sky130_fd_sc_hd__or3_1 _10420_ (.A(_04059_),
    .B(_02737_),
    .C(_04075_),
    .X(_05377_));
 sky130_fd_sc_hd__clkbuf_4 _10421_ (.A(_05377_),
    .X(_05378_));
 sky130_fd_sc_hd__buf_4 _10422_ (.A(_05378_),
    .X(_05379_));
 sky130_fd_sc_hd__mux2_1 _10423_ (.A0(_05211_),
    .A1(net515),
    .S(_05379_),
    .X(_05380_));
 sky130_fd_sc_hd__clkbuf_1 _10424_ (.A(_05380_),
    .X(_00433_));
 sky130_fd_sc_hd__mux2_1 _10425_ (.A0(_05216_),
    .A1(net638),
    .S(_05379_),
    .X(_05381_));
 sky130_fd_sc_hd__clkbuf_1 _10426_ (.A(_05381_),
    .X(_00434_));
 sky130_fd_sc_hd__mux2_1 _10427_ (.A0(_05218_),
    .A1(net1499),
    .S(_05379_),
    .X(_05382_));
 sky130_fd_sc_hd__clkbuf_1 _10428_ (.A(_05382_),
    .X(_00435_));
 sky130_fd_sc_hd__mux2_1 _10429_ (.A0(_05220_),
    .A1(net1192),
    .S(_05379_),
    .X(_05383_));
 sky130_fd_sc_hd__clkbuf_1 _10430_ (.A(_05383_),
    .X(_00436_));
 sky130_fd_sc_hd__mux2_1 _10431_ (.A0(_05222_),
    .A1(net280),
    .S(_05379_),
    .X(_05384_));
 sky130_fd_sc_hd__clkbuf_1 _10432_ (.A(_05384_),
    .X(_00437_));
 sky130_fd_sc_hd__mux2_1 _10433_ (.A0(_05224_),
    .A1(net764),
    .S(_05379_),
    .X(_05385_));
 sky130_fd_sc_hd__clkbuf_1 _10434_ (.A(_05385_),
    .X(_00438_));
 sky130_fd_sc_hd__mux2_1 _10435_ (.A0(_05226_),
    .A1(net799),
    .S(_05379_),
    .X(_05386_));
 sky130_fd_sc_hd__clkbuf_1 _10436_ (.A(_05386_),
    .X(_00439_));
 sky130_fd_sc_hd__mux2_1 _10437_ (.A0(_05228_),
    .A1(net393),
    .S(_05379_),
    .X(_05387_));
 sky130_fd_sc_hd__clkbuf_1 _10438_ (.A(_05387_),
    .X(_00440_));
 sky130_fd_sc_hd__mux2_1 _10439_ (.A0(_05230_),
    .A1(net937),
    .S(_05379_),
    .X(_05388_));
 sky130_fd_sc_hd__clkbuf_1 _10440_ (.A(_05388_),
    .X(_00441_));
 sky130_fd_sc_hd__mux2_1 _10441_ (.A0(_05232_),
    .A1(net615),
    .S(_05379_),
    .X(_05389_));
 sky130_fd_sc_hd__clkbuf_1 _10442_ (.A(_05389_),
    .X(_00442_));
 sky130_fd_sc_hd__mux2_1 _10443_ (.A0(_05234_),
    .A1(net1581),
    .S(_05378_),
    .X(_05390_));
 sky130_fd_sc_hd__clkbuf_1 _10444_ (.A(_05390_),
    .X(_00443_));
 sky130_fd_sc_hd__mux2_1 _10445_ (.A0(_05236_),
    .A1(net424),
    .S(_05378_),
    .X(_05391_));
 sky130_fd_sc_hd__clkbuf_1 _10446_ (.A(_05391_),
    .X(_00444_));
 sky130_fd_sc_hd__mux2_1 _10447_ (.A0(_05238_),
    .A1(net1660),
    .S(_05378_),
    .X(_05392_));
 sky130_fd_sc_hd__clkbuf_1 _10448_ (.A(_05392_),
    .X(_00445_));
 sky130_fd_sc_hd__mux2_1 _10449_ (.A0(_05240_),
    .A1(net1407),
    .S(_05378_),
    .X(_05393_));
 sky130_fd_sc_hd__clkbuf_1 _10450_ (.A(_05393_),
    .X(_00446_));
 sky130_fd_sc_hd__mux2_1 _10451_ (.A0(_05242_),
    .A1(net1197),
    .S(_05378_),
    .X(_05394_));
 sky130_fd_sc_hd__clkbuf_1 _10452_ (.A(_05394_),
    .X(_00447_));
 sky130_fd_sc_hd__mux2_1 _10453_ (.A0(_05244_),
    .A1(net887),
    .S(_05378_),
    .X(_05395_));
 sky130_fd_sc_hd__clkbuf_1 _10454_ (.A(_05395_),
    .X(_00448_));
 sky130_fd_sc_hd__nand2b_4 _10455_ (.A_N(_04076_),
    .B(_04408_),
    .Y(_05396_));
 sky130_fd_sc_hd__buf_4 _10456_ (.A(_05396_),
    .X(_05397_));
 sky130_fd_sc_hd__mux2_1 _10457_ (.A0(_05211_),
    .A1(net1741),
    .S(_05397_),
    .X(_05398_));
 sky130_fd_sc_hd__clkbuf_1 _10458_ (.A(_05398_),
    .X(_00449_));
 sky130_fd_sc_hd__mux2_1 _10459_ (.A0(_05216_),
    .A1(net1746),
    .S(_05397_),
    .X(_05399_));
 sky130_fd_sc_hd__clkbuf_1 _10460_ (.A(_05399_),
    .X(_00450_));
 sky130_fd_sc_hd__mux2_1 _10461_ (.A0(_05218_),
    .A1(net1542),
    .S(_05397_),
    .X(_05400_));
 sky130_fd_sc_hd__clkbuf_1 _10462_ (.A(_05400_),
    .X(_00451_));
 sky130_fd_sc_hd__mux2_1 _10463_ (.A0(_05220_),
    .A1(net1268),
    .S(_05397_),
    .X(_05401_));
 sky130_fd_sc_hd__clkbuf_1 _10464_ (.A(_05401_),
    .X(_00452_));
 sky130_fd_sc_hd__mux2_1 _10465_ (.A0(_05222_),
    .A1(net687),
    .S(_05397_),
    .X(_05402_));
 sky130_fd_sc_hd__clkbuf_1 _10466_ (.A(_05402_),
    .X(_00453_));
 sky130_fd_sc_hd__mux2_1 _10467_ (.A0(_05224_),
    .A1(net1215),
    .S(_05397_),
    .X(_05403_));
 sky130_fd_sc_hd__clkbuf_1 _10468_ (.A(_05403_),
    .X(_00454_));
 sky130_fd_sc_hd__mux2_1 _10469_ (.A0(_05226_),
    .A1(net1716),
    .S(_05397_),
    .X(_05404_));
 sky130_fd_sc_hd__clkbuf_1 _10470_ (.A(_05404_),
    .X(_00455_));
 sky130_fd_sc_hd__mux2_1 _10471_ (.A0(_05228_),
    .A1(net720),
    .S(_05397_),
    .X(_05405_));
 sky130_fd_sc_hd__clkbuf_1 _10472_ (.A(_05405_),
    .X(_00456_));
 sky130_fd_sc_hd__mux2_1 _10473_ (.A0(_05230_),
    .A1(net1420),
    .S(_05397_),
    .X(_05406_));
 sky130_fd_sc_hd__clkbuf_1 _10474_ (.A(_05406_),
    .X(_00457_));
 sky130_fd_sc_hd__mux2_1 _10475_ (.A0(_05232_),
    .A1(net1337),
    .S(_05397_),
    .X(_05407_));
 sky130_fd_sc_hd__clkbuf_1 _10476_ (.A(_05407_),
    .X(_00458_));
 sky130_fd_sc_hd__mux2_1 _10477_ (.A0(_05234_),
    .A1(net1258),
    .S(_05396_),
    .X(_05408_));
 sky130_fd_sc_hd__clkbuf_1 _10478_ (.A(_05408_),
    .X(_00459_));
 sky130_fd_sc_hd__mux2_1 _10479_ (.A0(_05236_),
    .A1(net812),
    .S(_05396_),
    .X(_05409_));
 sky130_fd_sc_hd__clkbuf_1 _10480_ (.A(_05409_),
    .X(_00460_));
 sky130_fd_sc_hd__mux2_1 _10481_ (.A0(_05238_),
    .A1(net1228),
    .S(_05396_),
    .X(_05410_));
 sky130_fd_sc_hd__clkbuf_1 _10482_ (.A(_05410_),
    .X(_00461_));
 sky130_fd_sc_hd__mux2_1 _10483_ (.A0(_05240_),
    .A1(net1945),
    .S(_05396_),
    .X(_05411_));
 sky130_fd_sc_hd__clkbuf_1 _10484_ (.A(_05411_),
    .X(_00462_));
 sky130_fd_sc_hd__mux2_1 _10485_ (.A0(_05242_),
    .A1(net1590),
    .S(_05396_),
    .X(_05412_));
 sky130_fd_sc_hd__clkbuf_1 _10486_ (.A(_05412_),
    .X(_00463_));
 sky130_fd_sc_hd__mux2_1 _10487_ (.A0(_05244_),
    .A1(net1663),
    .S(_05396_),
    .X(_05413_));
 sky130_fd_sc_hd__clkbuf_1 _10488_ (.A(_05413_),
    .X(_00464_));
 sky130_fd_sc_hd__or3_1 _10489_ (.A(_02484_),
    .B(_05026_),
    .C(_04075_),
    .X(_05414_));
 sky130_fd_sc_hd__clkbuf_4 _10490_ (.A(_05414_),
    .X(_05415_));
 sky130_fd_sc_hd__buf_4 _10491_ (.A(_05415_),
    .X(_05416_));
 sky130_fd_sc_hd__mux2_1 _10492_ (.A0(_05211_),
    .A1(net923),
    .S(_05416_),
    .X(_05417_));
 sky130_fd_sc_hd__clkbuf_1 _10493_ (.A(_05417_),
    .X(_00465_));
 sky130_fd_sc_hd__mux2_1 _10494_ (.A0(_05216_),
    .A1(net776),
    .S(_05416_),
    .X(_05418_));
 sky130_fd_sc_hd__clkbuf_1 _10495_ (.A(_05418_),
    .X(_00466_));
 sky130_fd_sc_hd__mux2_1 _10496_ (.A0(_05218_),
    .A1(net1453),
    .S(_05416_),
    .X(_05419_));
 sky130_fd_sc_hd__clkbuf_1 _10497_ (.A(_05419_),
    .X(_00467_));
 sky130_fd_sc_hd__mux2_1 _10498_ (.A0(_05220_),
    .A1(net1004),
    .S(_05416_),
    .X(_05420_));
 sky130_fd_sc_hd__clkbuf_1 _10499_ (.A(_05420_),
    .X(_00468_));
 sky130_fd_sc_hd__mux2_1 _10500_ (.A0(_05222_),
    .A1(net1807),
    .S(_05416_),
    .X(_05421_));
 sky130_fd_sc_hd__clkbuf_1 _10501_ (.A(_05421_),
    .X(_00469_));
 sky130_fd_sc_hd__mux2_1 _10502_ (.A0(_05224_),
    .A1(net1342),
    .S(_05416_),
    .X(_05422_));
 sky130_fd_sc_hd__clkbuf_1 _10503_ (.A(_05422_),
    .X(_00470_));
 sky130_fd_sc_hd__mux2_1 _10504_ (.A0(_05226_),
    .A1(net1753),
    .S(_05416_),
    .X(_05423_));
 sky130_fd_sc_hd__clkbuf_1 _10505_ (.A(_05423_),
    .X(_00471_));
 sky130_fd_sc_hd__mux2_1 _10506_ (.A0(_05228_),
    .A1(net731),
    .S(_05416_),
    .X(_05424_));
 sky130_fd_sc_hd__clkbuf_1 _10507_ (.A(_05424_),
    .X(_00472_));
 sky130_fd_sc_hd__mux2_1 _10508_ (.A0(_05230_),
    .A1(net1295),
    .S(_05416_),
    .X(_05425_));
 sky130_fd_sc_hd__clkbuf_1 _10509_ (.A(_05425_),
    .X(_00473_));
 sky130_fd_sc_hd__mux2_1 _10510_ (.A0(_05232_),
    .A1(net1302),
    .S(_05416_),
    .X(_05426_));
 sky130_fd_sc_hd__clkbuf_1 _10511_ (.A(_05426_),
    .X(_00474_));
 sky130_fd_sc_hd__mux2_1 _10512_ (.A0(_05234_),
    .A1(net1461),
    .S(_05415_),
    .X(_05427_));
 sky130_fd_sc_hd__clkbuf_1 _10513_ (.A(_05427_),
    .X(_00475_));
 sky130_fd_sc_hd__mux2_1 _10514_ (.A0(_05236_),
    .A1(net1761),
    .S(_05415_),
    .X(_05428_));
 sky130_fd_sc_hd__clkbuf_1 _10515_ (.A(_05428_),
    .X(_00476_));
 sky130_fd_sc_hd__mux2_1 _10516_ (.A0(_05238_),
    .A1(net934),
    .S(_05415_),
    .X(_05429_));
 sky130_fd_sc_hd__clkbuf_1 _10517_ (.A(_05429_),
    .X(_00477_));
 sky130_fd_sc_hd__mux2_1 _10518_ (.A0(_05240_),
    .A1(net1858),
    .S(_05415_),
    .X(_05430_));
 sky130_fd_sc_hd__clkbuf_1 _10519_ (.A(_05430_),
    .X(_00478_));
 sky130_fd_sc_hd__mux2_1 _10520_ (.A0(_05242_),
    .A1(net752),
    .S(_05415_),
    .X(_05431_));
 sky130_fd_sc_hd__clkbuf_1 _10521_ (.A(_05431_),
    .X(_00479_));
 sky130_fd_sc_hd__mux2_1 _10522_ (.A0(_05244_),
    .A1(net1652),
    .S(_05415_),
    .X(_05432_));
 sky130_fd_sc_hd__clkbuf_1 _10523_ (.A(_05432_),
    .X(_00480_));
 sky130_fd_sc_hd__nor2_4 _10524_ (.A(_04186_),
    .B(_04461_),
    .Y(_05433_));
 sky130_fd_sc_hd__buf_4 _10525_ (.A(_05433_),
    .X(_05434_));
 sky130_fd_sc_hd__mux2_1 _10526_ (.A0(net1183),
    .A1(_04992_),
    .S(_05434_),
    .X(_05435_));
 sky130_fd_sc_hd__clkbuf_1 _10527_ (.A(_05435_),
    .X(_00481_));
 sky130_fd_sc_hd__mux2_1 _10528_ (.A0(net1448),
    .A1(_04996_),
    .S(_05434_),
    .X(_05436_));
 sky130_fd_sc_hd__clkbuf_1 _10529_ (.A(_05436_),
    .X(_00482_));
 sky130_fd_sc_hd__mux2_1 _10530_ (.A0(net331),
    .A1(_04998_),
    .S(_05434_),
    .X(_05437_));
 sky130_fd_sc_hd__clkbuf_1 _10531_ (.A(_05437_),
    .X(_00483_));
 sky130_fd_sc_hd__mux2_1 _10532_ (.A0(net841),
    .A1(_05000_),
    .S(_05434_),
    .X(_05438_));
 sky130_fd_sc_hd__clkbuf_1 _10533_ (.A(_05438_),
    .X(_00484_));
 sky130_fd_sc_hd__mux2_1 _10534_ (.A0(net959),
    .A1(_05002_),
    .S(_05434_),
    .X(_05439_));
 sky130_fd_sc_hd__clkbuf_1 _10535_ (.A(_05439_),
    .X(_00485_));
 sky130_fd_sc_hd__mux2_1 _10536_ (.A0(net925),
    .A1(_05004_),
    .S(_05434_),
    .X(_05440_));
 sky130_fd_sc_hd__clkbuf_1 _10537_ (.A(_05440_),
    .X(_00486_));
 sky130_fd_sc_hd__mux2_1 _10538_ (.A0(net1294),
    .A1(_05006_),
    .S(_05434_),
    .X(_05441_));
 sky130_fd_sc_hd__clkbuf_1 _10539_ (.A(_05441_),
    .X(_00487_));
 sky130_fd_sc_hd__mux2_1 _10540_ (.A0(net723),
    .A1(_05008_),
    .S(_05434_),
    .X(_05442_));
 sky130_fd_sc_hd__clkbuf_1 _10541_ (.A(_05442_),
    .X(_00488_));
 sky130_fd_sc_hd__mux2_1 _10542_ (.A0(net829),
    .A1(_05010_),
    .S(_05434_),
    .X(_05443_));
 sky130_fd_sc_hd__clkbuf_1 _10543_ (.A(_05443_),
    .X(_00489_));
 sky130_fd_sc_hd__mux2_1 _10544_ (.A0(net1246),
    .A1(_05012_),
    .S(_05434_),
    .X(_05444_));
 sky130_fd_sc_hd__clkbuf_1 _10545_ (.A(_05444_),
    .X(_00490_));
 sky130_fd_sc_hd__mux2_1 _10546_ (.A0(net1212),
    .A1(_05014_),
    .S(_05433_),
    .X(_05445_));
 sky130_fd_sc_hd__clkbuf_1 _10547_ (.A(_05445_),
    .X(_00491_));
 sky130_fd_sc_hd__mux2_1 _10548_ (.A0(net860),
    .A1(_05016_),
    .S(_05433_),
    .X(_05446_));
 sky130_fd_sc_hd__clkbuf_1 _10549_ (.A(_05446_),
    .X(_00492_));
 sky130_fd_sc_hd__mux2_1 _10550_ (.A0(net1368),
    .A1(_05018_),
    .S(_05433_),
    .X(_05447_));
 sky130_fd_sc_hd__clkbuf_1 _10551_ (.A(_05447_),
    .X(_00493_));
 sky130_fd_sc_hd__mux2_1 _10552_ (.A0(net356),
    .A1(_05020_),
    .S(_05433_),
    .X(_05448_));
 sky130_fd_sc_hd__clkbuf_1 _10553_ (.A(_05448_),
    .X(_00494_));
 sky130_fd_sc_hd__mux2_1 _10554_ (.A0(net996),
    .A1(_05022_),
    .S(_05433_),
    .X(_05449_));
 sky130_fd_sc_hd__clkbuf_1 _10555_ (.A(_05449_),
    .X(_00495_));
 sky130_fd_sc_hd__mux2_1 _10556_ (.A0(net793),
    .A1(_05024_),
    .S(_05433_),
    .X(_05450_));
 sky130_fd_sc_hd__clkbuf_1 _10557_ (.A(_05450_),
    .X(_00496_));
 sky130_fd_sc_hd__nor2_4 _10558_ (.A(_04072_),
    .B(_04186_),
    .Y(_05451_));
 sky130_fd_sc_hd__buf_4 _10559_ (.A(_05451_),
    .X(_05452_));
 sky130_fd_sc_hd__mux2_1 _10560_ (.A0(net1353),
    .A1(_04992_),
    .S(_05452_),
    .X(_05453_));
 sky130_fd_sc_hd__clkbuf_1 _10561_ (.A(_05453_),
    .X(_00497_));
 sky130_fd_sc_hd__mux2_1 _10562_ (.A0(net1061),
    .A1(_04996_),
    .S(_05452_),
    .X(_05454_));
 sky130_fd_sc_hd__clkbuf_1 _10563_ (.A(_05454_),
    .X(_00498_));
 sky130_fd_sc_hd__mux2_1 _10564_ (.A0(net642),
    .A1(_04998_),
    .S(_05452_),
    .X(_05455_));
 sky130_fd_sc_hd__clkbuf_1 _10565_ (.A(_05455_),
    .X(_00499_));
 sky130_fd_sc_hd__mux2_1 _10566_ (.A0(net1821),
    .A1(_05000_),
    .S(_05452_),
    .X(_05456_));
 sky130_fd_sc_hd__clkbuf_1 _10567_ (.A(_05456_),
    .X(_00500_));
 sky130_fd_sc_hd__mux2_1 _10568_ (.A0(net834),
    .A1(_05002_),
    .S(_05452_),
    .X(_05457_));
 sky130_fd_sc_hd__clkbuf_1 _10569_ (.A(_05457_),
    .X(_00501_));
 sky130_fd_sc_hd__mux2_1 _10570_ (.A0(net1669),
    .A1(_05004_),
    .S(_05452_),
    .X(_05458_));
 sky130_fd_sc_hd__clkbuf_1 _10571_ (.A(_05458_),
    .X(_00502_));
 sky130_fd_sc_hd__mux2_1 _10572_ (.A0(net988),
    .A1(_05006_),
    .S(_05452_),
    .X(_05459_));
 sky130_fd_sc_hd__clkbuf_1 _10573_ (.A(_05459_),
    .X(_00503_));
 sky130_fd_sc_hd__mux2_1 _10574_ (.A0(net1071),
    .A1(_05008_),
    .S(_05452_),
    .X(_05460_));
 sky130_fd_sc_hd__clkbuf_1 _10575_ (.A(_05460_),
    .X(_00504_));
 sky130_fd_sc_hd__mux2_1 _10576_ (.A0(net1111),
    .A1(_05010_),
    .S(_05452_),
    .X(_05461_));
 sky130_fd_sc_hd__clkbuf_1 _10577_ (.A(_05461_),
    .X(_00505_));
 sky130_fd_sc_hd__mux2_1 _10578_ (.A0(net1129),
    .A1(_05012_),
    .S(_05452_),
    .X(_05462_));
 sky130_fd_sc_hd__clkbuf_1 _10579_ (.A(_05462_),
    .X(_00506_));
 sky130_fd_sc_hd__mux2_1 _10580_ (.A0(net983),
    .A1(_05014_),
    .S(_05451_),
    .X(_05463_));
 sky130_fd_sc_hd__clkbuf_1 _10581_ (.A(_05463_),
    .X(_00507_));
 sky130_fd_sc_hd__mux2_1 _10582_ (.A0(net1878),
    .A1(_05016_),
    .S(_05451_),
    .X(_05464_));
 sky130_fd_sc_hd__clkbuf_1 _10583_ (.A(_05464_),
    .X(_00508_));
 sky130_fd_sc_hd__mux2_1 _10584_ (.A0(net1839),
    .A1(_05018_),
    .S(_05451_),
    .X(_05465_));
 sky130_fd_sc_hd__clkbuf_1 _10585_ (.A(_05465_),
    .X(_00509_));
 sky130_fd_sc_hd__mux2_1 _10586_ (.A0(net1535),
    .A1(_05020_),
    .S(_05451_),
    .X(_05466_));
 sky130_fd_sc_hd__clkbuf_1 _10587_ (.A(_05466_),
    .X(_00510_));
 sky130_fd_sc_hd__mux2_1 _10588_ (.A0(net1480),
    .A1(_05022_),
    .S(_05451_),
    .X(_05467_));
 sky130_fd_sc_hd__clkbuf_1 _10589_ (.A(_05467_),
    .X(_00511_));
 sky130_fd_sc_hd__mux2_1 _10590_ (.A0(net1508),
    .A1(_05024_),
    .S(_05451_),
    .X(_05468_));
 sky130_fd_sc_hd__clkbuf_1 _10591_ (.A(_05468_),
    .X(_00512_));
 sky130_fd_sc_hd__buf_6 _10592_ (.A(_04069_),
    .X(_05469_));
 sky130_fd_sc_hd__nor2_4 _10593_ (.A(_04186_),
    .B(_04501_),
    .Y(_05470_));
 sky130_fd_sc_hd__buf_4 _10594_ (.A(_05470_),
    .X(_05471_));
 sky130_fd_sc_hd__mux2_1 _10595_ (.A0(net1112),
    .A1(_05469_),
    .S(_05471_),
    .X(_05472_));
 sky130_fd_sc_hd__clkbuf_1 _10596_ (.A(_05472_),
    .X(_00513_));
 sky130_fd_sc_hd__clkbuf_4 _10597_ (.A(_04080_),
    .X(_05473_));
 sky130_fd_sc_hd__mux2_1 _10598_ (.A0(net671),
    .A1(_05473_),
    .S(_05471_),
    .X(_05474_));
 sky130_fd_sc_hd__clkbuf_1 _10599_ (.A(_05474_),
    .X(_00514_));
 sky130_fd_sc_hd__buf_6 _10600_ (.A(_04083_),
    .X(_05475_));
 sky130_fd_sc_hd__mux2_1 _10601_ (.A0(net1985),
    .A1(_05475_),
    .S(_05471_),
    .X(_05476_));
 sky130_fd_sc_hd__clkbuf_1 _10602_ (.A(_05476_),
    .X(_00515_));
 sky130_fd_sc_hd__buf_6 _10603_ (.A(_04086_),
    .X(_05477_));
 sky130_fd_sc_hd__mux2_1 _10604_ (.A0(net1455),
    .A1(_05477_),
    .S(_05471_),
    .X(_05478_));
 sky130_fd_sc_hd__clkbuf_1 _10605_ (.A(_05478_),
    .X(_00516_));
 sky130_fd_sc_hd__buf_4 _10606_ (.A(_04089_),
    .X(_05479_));
 sky130_fd_sc_hd__mux2_1 _10607_ (.A0(net1703),
    .A1(_05479_),
    .S(_05471_),
    .X(_05480_));
 sky130_fd_sc_hd__clkbuf_1 _10608_ (.A(_05480_),
    .X(_00517_));
 sky130_fd_sc_hd__clkbuf_4 _10609_ (.A(_04092_),
    .X(_05481_));
 sky130_fd_sc_hd__mux2_1 _10610_ (.A0(net1412),
    .A1(_05481_),
    .S(_05471_),
    .X(_05482_));
 sky130_fd_sc_hd__clkbuf_1 _10611_ (.A(_05482_),
    .X(_00518_));
 sky130_fd_sc_hd__clkbuf_4 _10612_ (.A(_04095_),
    .X(_05483_));
 sky130_fd_sc_hd__mux2_1 _10613_ (.A0(net1802),
    .A1(_05483_),
    .S(_05471_),
    .X(_05484_));
 sky130_fd_sc_hd__clkbuf_1 _10614_ (.A(_05484_),
    .X(_00519_));
 sky130_fd_sc_hd__buf_4 _10615_ (.A(_04098_),
    .X(_05485_));
 sky130_fd_sc_hd__mux2_1 _10616_ (.A0(net1577),
    .A1(_05485_),
    .S(_05471_),
    .X(_05486_));
 sky130_fd_sc_hd__clkbuf_1 _10617_ (.A(_05486_),
    .X(_00520_));
 sky130_fd_sc_hd__buf_4 _10618_ (.A(_04101_),
    .X(_05487_));
 sky130_fd_sc_hd__mux2_1 _10619_ (.A0(net946),
    .A1(_05487_),
    .S(_05471_),
    .X(_05488_));
 sky130_fd_sc_hd__clkbuf_1 _10620_ (.A(_05488_),
    .X(_00521_));
 sky130_fd_sc_hd__buf_4 _10621_ (.A(_04104_),
    .X(_05489_));
 sky130_fd_sc_hd__mux2_1 _10622_ (.A0(net1313),
    .A1(_05489_),
    .S(_05471_),
    .X(_05490_));
 sky130_fd_sc_hd__clkbuf_1 _10623_ (.A(_05490_),
    .X(_00522_));
 sky130_fd_sc_hd__clkbuf_4 _10624_ (.A(_04107_),
    .X(_05491_));
 sky130_fd_sc_hd__mux2_1 _10625_ (.A0(net1358),
    .A1(_05491_),
    .S(_05470_),
    .X(_05492_));
 sky130_fd_sc_hd__clkbuf_1 _10626_ (.A(_05492_),
    .X(_00523_));
 sky130_fd_sc_hd__clkbuf_4 _10627_ (.A(_04110_),
    .X(_05493_));
 sky130_fd_sc_hd__mux2_1 _10628_ (.A0(net890),
    .A1(_05493_),
    .S(_05470_),
    .X(_05494_));
 sky130_fd_sc_hd__clkbuf_1 _10629_ (.A(_05494_),
    .X(_00524_));
 sky130_fd_sc_hd__clkbuf_4 _10630_ (.A(_04113_),
    .X(_05495_));
 sky130_fd_sc_hd__mux2_1 _10631_ (.A0(net479),
    .A1(_05495_),
    .S(_05470_),
    .X(_05496_));
 sky130_fd_sc_hd__clkbuf_1 _10632_ (.A(_05496_),
    .X(_00525_));
 sky130_fd_sc_hd__clkbuf_4 _10633_ (.A(_04116_),
    .X(_05497_));
 sky130_fd_sc_hd__mux2_1 _10634_ (.A0(net780),
    .A1(_05497_),
    .S(_05470_),
    .X(_05498_));
 sky130_fd_sc_hd__clkbuf_1 _10635_ (.A(_05498_),
    .X(_00526_));
 sky130_fd_sc_hd__clkbuf_4 _10636_ (.A(_04119_),
    .X(_05499_));
 sky130_fd_sc_hd__mux2_1 _10637_ (.A0(net1445),
    .A1(_05499_),
    .S(_05470_),
    .X(_05500_));
 sky130_fd_sc_hd__clkbuf_1 _10638_ (.A(_05500_),
    .X(_00527_));
 sky130_fd_sc_hd__clkbuf_4 _10639_ (.A(_04122_),
    .X(_05501_));
 sky130_fd_sc_hd__mux2_1 _10640_ (.A0(net1299),
    .A1(_05501_),
    .S(_05470_),
    .X(_05502_));
 sky130_fd_sc_hd__clkbuf_1 _10641_ (.A(_05502_),
    .X(_00528_));
 sky130_fd_sc_hd__nor2_4 _10642_ (.A(_04186_),
    .B(_04225_),
    .Y(_05503_));
 sky130_fd_sc_hd__buf_4 _10643_ (.A(_05503_),
    .X(_05504_));
 sky130_fd_sc_hd__mux2_1 _10644_ (.A0(net1591),
    .A1(_05469_),
    .S(_05504_),
    .X(_05505_));
 sky130_fd_sc_hd__clkbuf_1 _10645_ (.A(_05505_),
    .X(_00529_));
 sky130_fd_sc_hd__mux2_1 _10646_ (.A0(net1249),
    .A1(_05473_),
    .S(_05504_),
    .X(_05506_));
 sky130_fd_sc_hd__clkbuf_1 _10647_ (.A(_05506_),
    .X(_00530_));
 sky130_fd_sc_hd__mux2_1 _10648_ (.A0(net2055),
    .A1(_05475_),
    .S(_05504_),
    .X(_05507_));
 sky130_fd_sc_hd__clkbuf_1 _10649_ (.A(_05507_),
    .X(_00531_));
 sky130_fd_sc_hd__mux2_1 _10650_ (.A0(net1585),
    .A1(_05477_),
    .S(_05504_),
    .X(_05508_));
 sky130_fd_sc_hd__clkbuf_1 _10651_ (.A(_05508_),
    .X(_00532_));
 sky130_fd_sc_hd__mux2_1 _10652_ (.A0(net1933),
    .A1(_05479_),
    .S(_05504_),
    .X(_05509_));
 sky130_fd_sc_hd__clkbuf_1 _10653_ (.A(_05509_),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_1 _10654_ (.A0(net746),
    .A1(_05481_),
    .S(_05504_),
    .X(_05510_));
 sky130_fd_sc_hd__clkbuf_1 _10655_ (.A(_05510_),
    .X(_00534_));
 sky130_fd_sc_hd__mux2_1 _10656_ (.A0(net1149),
    .A1(_05483_),
    .S(_05504_),
    .X(_05511_));
 sky130_fd_sc_hd__clkbuf_1 _10657_ (.A(_05511_),
    .X(_00535_));
 sky130_fd_sc_hd__mux2_1 _10658_ (.A0(net1987),
    .A1(_05485_),
    .S(_05504_),
    .X(_05512_));
 sky130_fd_sc_hd__clkbuf_1 _10659_ (.A(_05512_),
    .X(_00536_));
 sky130_fd_sc_hd__mux2_1 _10660_ (.A0(net1726),
    .A1(_05487_),
    .S(_05504_),
    .X(_05513_));
 sky130_fd_sc_hd__clkbuf_1 _10661_ (.A(_05513_),
    .X(_00537_));
 sky130_fd_sc_hd__mux2_1 _10662_ (.A0(net1288),
    .A1(_05489_),
    .S(_05504_),
    .X(_05514_));
 sky130_fd_sc_hd__clkbuf_1 _10663_ (.A(_05514_),
    .X(_00538_));
 sky130_fd_sc_hd__mux2_1 _10664_ (.A0(net788),
    .A1(_05491_),
    .S(_05503_),
    .X(_05515_));
 sky130_fd_sc_hd__clkbuf_1 _10665_ (.A(_05515_),
    .X(_00539_));
 sky130_fd_sc_hd__mux2_1 _10666_ (.A0(net577),
    .A1(_05493_),
    .S(_05503_),
    .X(_05516_));
 sky130_fd_sc_hd__clkbuf_1 _10667_ (.A(_05516_),
    .X(_00540_));
 sky130_fd_sc_hd__mux2_1 _10668_ (.A0(net761),
    .A1(_05495_),
    .S(_05503_),
    .X(_05517_));
 sky130_fd_sc_hd__clkbuf_1 _10669_ (.A(_05517_),
    .X(_00541_));
 sky130_fd_sc_hd__mux2_1 _10670_ (.A0(net1259),
    .A1(_05497_),
    .S(_05503_),
    .X(_05518_));
 sky130_fd_sc_hd__clkbuf_1 _10671_ (.A(_05518_),
    .X(_00542_));
 sky130_fd_sc_hd__mux2_1 _10672_ (.A0(net1271),
    .A1(_05499_),
    .S(_05503_),
    .X(_05519_));
 sky130_fd_sc_hd__clkbuf_1 _10673_ (.A(_05519_),
    .X(_00543_));
 sky130_fd_sc_hd__mux2_1 _10674_ (.A0(net809),
    .A1(_05501_),
    .S(_05503_),
    .X(_05520_));
 sky130_fd_sc_hd__clkbuf_1 _10675_ (.A(_05520_),
    .X(_00544_));
 sky130_fd_sc_hd__nor2_4 _10676_ (.A(_04186_),
    .B(_04569_),
    .Y(_05521_));
 sky130_fd_sc_hd__buf_4 _10677_ (.A(_05521_),
    .X(_05522_));
 sky130_fd_sc_hd__mux2_1 _10678_ (.A0(net1722),
    .A1(_05469_),
    .S(_05522_),
    .X(_05523_));
 sky130_fd_sc_hd__clkbuf_1 _10679_ (.A(_05523_),
    .X(_00545_));
 sky130_fd_sc_hd__mux2_1 _10680_ (.A0(net148),
    .A1(_05473_),
    .S(_05522_),
    .X(_05524_));
 sky130_fd_sc_hd__clkbuf_1 _10681_ (.A(_05524_),
    .X(_00546_));
 sky130_fd_sc_hd__mux2_1 _10682_ (.A0(net1584),
    .A1(_05475_),
    .S(_05522_),
    .X(_05525_));
 sky130_fd_sc_hd__clkbuf_1 _10683_ (.A(_05525_),
    .X(_00547_));
 sky130_fd_sc_hd__mux2_1 _10684_ (.A0(net1418),
    .A1(_05477_),
    .S(_05522_),
    .X(_05526_));
 sky130_fd_sc_hd__clkbuf_1 _10685_ (.A(_05526_),
    .X(_00548_));
 sky130_fd_sc_hd__mux2_1 _10686_ (.A0(net55),
    .A1(_05479_),
    .S(_05522_),
    .X(_05527_));
 sky130_fd_sc_hd__clkbuf_1 _10687_ (.A(_05527_),
    .X(_00549_));
 sky130_fd_sc_hd__mux2_1 _10688_ (.A0(net144),
    .A1(_05481_),
    .S(_05522_),
    .X(_05528_));
 sky130_fd_sc_hd__clkbuf_1 _10689_ (.A(_05528_),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_1 _10690_ (.A0(net184),
    .A1(_05483_),
    .S(_05522_),
    .X(_05529_));
 sky130_fd_sc_hd__clkbuf_1 _10691_ (.A(_05529_),
    .X(_00551_));
 sky130_fd_sc_hd__mux2_1 _10692_ (.A0(net406),
    .A1(_05485_),
    .S(_05522_),
    .X(_05530_));
 sky130_fd_sc_hd__clkbuf_1 _10693_ (.A(_05530_),
    .X(_00552_));
 sky130_fd_sc_hd__mux2_1 _10694_ (.A0(net158),
    .A1(_05487_),
    .S(_05522_),
    .X(_05531_));
 sky130_fd_sc_hd__clkbuf_1 _10695_ (.A(_05531_),
    .X(_00553_));
 sky130_fd_sc_hd__mux2_1 _10696_ (.A0(net75),
    .A1(_05489_),
    .S(_05522_),
    .X(_05532_));
 sky130_fd_sc_hd__clkbuf_1 _10697_ (.A(_05532_),
    .X(_00554_));
 sky130_fd_sc_hd__mux2_1 _10698_ (.A0(net69),
    .A1(_05491_),
    .S(_05521_),
    .X(_05533_));
 sky130_fd_sc_hd__clkbuf_1 _10699_ (.A(_05533_),
    .X(_00555_));
 sky130_fd_sc_hd__mux2_1 _10700_ (.A0(net61),
    .A1(_05493_),
    .S(_05521_),
    .X(_05534_));
 sky130_fd_sc_hd__clkbuf_1 _10701_ (.A(_05534_),
    .X(_00556_));
 sky130_fd_sc_hd__mux2_1 _10702_ (.A0(net114),
    .A1(_05495_),
    .S(_05521_),
    .X(_05535_));
 sky130_fd_sc_hd__clkbuf_1 _10703_ (.A(_05535_),
    .X(_00557_));
 sky130_fd_sc_hd__mux2_1 _10704_ (.A0(net195),
    .A1(_05497_),
    .S(_05521_),
    .X(_05536_));
 sky130_fd_sc_hd__clkbuf_1 _10705_ (.A(_05536_),
    .X(_00558_));
 sky130_fd_sc_hd__mux2_1 _10706_ (.A0(net455),
    .A1(_05499_),
    .S(_05521_),
    .X(_05537_));
 sky130_fd_sc_hd__clkbuf_1 _10707_ (.A(_05537_),
    .X(_00559_));
 sky130_fd_sc_hd__mux2_1 _10708_ (.A0(net149),
    .A1(_05501_),
    .S(_05521_),
    .X(_05538_));
 sky130_fd_sc_hd__clkbuf_1 _10709_ (.A(_05538_),
    .X(_00560_));
 sky130_fd_sc_hd__nor2_4 _10710_ (.A(_04368_),
    .B(_04607_),
    .Y(_05539_));
 sky130_fd_sc_hd__buf_4 _10711_ (.A(_05539_),
    .X(_05540_));
 sky130_fd_sc_hd__mux2_1 _10712_ (.A0(net1755),
    .A1(_05469_),
    .S(_05540_),
    .X(_05541_));
 sky130_fd_sc_hd__clkbuf_1 _10713_ (.A(_05541_),
    .X(_00561_));
 sky130_fd_sc_hd__mux2_1 _10714_ (.A0(net343),
    .A1(_05473_),
    .S(_05540_),
    .X(_05542_));
 sky130_fd_sc_hd__clkbuf_1 _10715_ (.A(_05542_),
    .X(_00562_));
 sky130_fd_sc_hd__mux2_1 _10716_ (.A0(net1730),
    .A1(_05475_),
    .S(_05540_),
    .X(_05543_));
 sky130_fd_sc_hd__clkbuf_1 _10717_ (.A(_05543_),
    .X(_00563_));
 sky130_fd_sc_hd__mux2_1 _10718_ (.A0(net1913),
    .A1(_05477_),
    .S(_05540_),
    .X(_05544_));
 sky130_fd_sc_hd__clkbuf_1 _10719_ (.A(_05544_),
    .X(_00564_));
 sky130_fd_sc_hd__mux2_1 _10720_ (.A0(net1639),
    .A1(_05479_),
    .S(_05540_),
    .X(_05545_));
 sky130_fd_sc_hd__clkbuf_1 _10721_ (.A(_05545_),
    .X(_00565_));
 sky130_fd_sc_hd__mux2_1 _10722_ (.A0(net1715),
    .A1(_05481_),
    .S(_05540_),
    .X(_05546_));
 sky130_fd_sc_hd__clkbuf_1 _10723_ (.A(_05546_),
    .X(_00566_));
 sky130_fd_sc_hd__mux2_1 _10724_ (.A0(net1831),
    .A1(_05483_),
    .S(_05540_),
    .X(_05547_));
 sky130_fd_sc_hd__clkbuf_1 _10725_ (.A(_05547_),
    .X(_00567_));
 sky130_fd_sc_hd__mux2_1 _10726_ (.A0(net853),
    .A1(_05485_),
    .S(_05540_),
    .X(_05548_));
 sky130_fd_sc_hd__clkbuf_1 _10727_ (.A(_05548_),
    .X(_00568_));
 sky130_fd_sc_hd__mux2_1 _10728_ (.A0(net1373),
    .A1(_05487_),
    .S(_05540_),
    .X(_05549_));
 sky130_fd_sc_hd__clkbuf_1 _10729_ (.A(_05549_),
    .X(_00569_));
 sky130_fd_sc_hd__mux2_1 _10730_ (.A0(net1293),
    .A1(_05489_),
    .S(_05540_),
    .X(_05550_));
 sky130_fd_sc_hd__clkbuf_1 _10731_ (.A(_05550_),
    .X(_00570_));
 sky130_fd_sc_hd__mux2_1 _10732_ (.A0(net1626),
    .A1(_05491_),
    .S(_05539_),
    .X(_05551_));
 sky130_fd_sc_hd__clkbuf_1 _10733_ (.A(_05551_),
    .X(_00571_));
 sky130_fd_sc_hd__mux2_1 _10734_ (.A0(net1066),
    .A1(_05493_),
    .S(_05539_),
    .X(_05552_));
 sky130_fd_sc_hd__clkbuf_1 _10735_ (.A(_05552_),
    .X(_00572_));
 sky130_fd_sc_hd__mux2_1 _10736_ (.A0(net992),
    .A1(_05495_),
    .S(_05539_),
    .X(_05553_));
 sky130_fd_sc_hd__clkbuf_1 _10737_ (.A(_05553_),
    .X(_00573_));
 sky130_fd_sc_hd__mux2_1 _10738_ (.A0(net1180),
    .A1(_05497_),
    .S(_05539_),
    .X(_05554_));
 sky130_fd_sc_hd__clkbuf_1 _10739_ (.A(_05554_),
    .X(_00574_));
 sky130_fd_sc_hd__mux2_1 _10740_ (.A0(net1351),
    .A1(_05499_),
    .S(_05539_),
    .X(_05555_));
 sky130_fd_sc_hd__clkbuf_1 _10741_ (.A(_05555_),
    .X(_00575_));
 sky130_fd_sc_hd__mux2_1 _10742_ (.A0(net912),
    .A1(_05501_),
    .S(_05539_),
    .X(_05556_));
 sky130_fd_sc_hd__clkbuf_1 _10743_ (.A(_05556_),
    .X(_00576_));
 sky130_fd_sc_hd__nor2_4 _10744_ (.A(_04186_),
    .B(_04607_),
    .Y(_05557_));
 sky130_fd_sc_hd__buf_4 _10745_ (.A(_05557_),
    .X(_05558_));
 sky130_fd_sc_hd__mux2_1 _10746_ (.A0(net1087),
    .A1(_05469_),
    .S(_05558_),
    .X(_05559_));
 sky130_fd_sc_hd__clkbuf_1 _10747_ (.A(_05559_),
    .X(_00577_));
 sky130_fd_sc_hd__mux2_1 _10748_ (.A0(net1128),
    .A1(_05473_),
    .S(_05558_),
    .X(_05560_));
 sky130_fd_sc_hd__clkbuf_1 _10749_ (.A(_05560_),
    .X(_00578_));
 sky130_fd_sc_hd__mux2_1 _10750_ (.A0(net1321),
    .A1(_05475_),
    .S(_05558_),
    .X(_05561_));
 sky130_fd_sc_hd__clkbuf_1 _10751_ (.A(_05561_),
    .X(_00579_));
 sky130_fd_sc_hd__mux2_1 _10752_ (.A0(net1208),
    .A1(_05477_),
    .S(_05558_),
    .X(_05562_));
 sky130_fd_sc_hd__clkbuf_1 _10753_ (.A(_05562_),
    .X(_00580_));
 sky130_fd_sc_hd__mux2_1 _10754_ (.A0(net1072),
    .A1(_05479_),
    .S(_05558_),
    .X(_05563_));
 sky130_fd_sc_hd__clkbuf_1 _10755_ (.A(_05563_),
    .X(_00581_));
 sky130_fd_sc_hd__mux2_1 _10756_ (.A0(net1692),
    .A1(_05481_),
    .S(_05558_),
    .X(_05564_));
 sky130_fd_sc_hd__clkbuf_1 _10757_ (.A(_05564_),
    .X(_00582_));
 sky130_fd_sc_hd__mux2_1 _10758_ (.A0(net1320),
    .A1(_05483_),
    .S(_05558_),
    .X(_05565_));
 sky130_fd_sc_hd__clkbuf_1 _10759_ (.A(_05565_),
    .X(_00583_));
 sky130_fd_sc_hd__mux2_1 _10760_ (.A0(net1166),
    .A1(_05485_),
    .S(_05558_),
    .X(_05566_));
 sky130_fd_sc_hd__clkbuf_1 _10761_ (.A(_05566_),
    .X(_00584_));
 sky130_fd_sc_hd__mux2_1 _10762_ (.A0(net1140),
    .A1(_05487_),
    .S(_05558_),
    .X(_05567_));
 sky130_fd_sc_hd__clkbuf_1 _10763_ (.A(_05567_),
    .X(_00585_));
 sky130_fd_sc_hd__mux2_1 _10764_ (.A0(net1887),
    .A1(_05489_),
    .S(_05558_),
    .X(_05568_));
 sky130_fd_sc_hd__clkbuf_1 _10765_ (.A(_05568_),
    .X(_00586_));
 sky130_fd_sc_hd__mux2_1 _10766_ (.A0(net798),
    .A1(_05491_),
    .S(_05557_),
    .X(_05569_));
 sky130_fd_sc_hd__clkbuf_1 _10767_ (.A(_05569_),
    .X(_00587_));
 sky130_fd_sc_hd__mux2_1 _10768_ (.A0(net968),
    .A1(_05493_),
    .S(_05557_),
    .X(_05570_));
 sky130_fd_sc_hd__clkbuf_1 _10769_ (.A(_05570_),
    .X(_00588_));
 sky130_fd_sc_hd__mux2_1 _10770_ (.A0(net1454),
    .A1(_05495_),
    .S(_05557_),
    .X(_05571_));
 sky130_fd_sc_hd__clkbuf_1 _10771_ (.A(_05571_),
    .X(_00589_));
 sky130_fd_sc_hd__mux2_1 _10772_ (.A0(net673),
    .A1(_05497_),
    .S(_05557_),
    .X(_05572_));
 sky130_fd_sc_hd__clkbuf_1 _10773_ (.A(_05572_),
    .X(_00590_));
 sky130_fd_sc_hd__mux2_1 _10774_ (.A0(net969),
    .A1(_05499_),
    .S(_05557_),
    .X(_05573_));
 sky130_fd_sc_hd__clkbuf_1 _10775_ (.A(_05573_),
    .X(_00591_));
 sky130_fd_sc_hd__mux2_1 _10776_ (.A0(net652),
    .A1(_05501_),
    .S(_05557_),
    .X(_05574_));
 sky130_fd_sc_hd__clkbuf_1 _10777_ (.A(_05574_),
    .X(_00592_));
 sky130_fd_sc_hd__or3_1 _10778_ (.A(_02498_),
    .B(_05026_),
    .C(_04185_),
    .X(_05575_));
 sky130_fd_sc_hd__buf_2 _10779_ (.A(_05575_),
    .X(_05576_));
 sky130_fd_sc_hd__buf_4 _10780_ (.A(_05576_),
    .X(_05577_));
 sky130_fd_sc_hd__mux2_1 _10781_ (.A0(_05211_),
    .A1(net1979),
    .S(_05577_),
    .X(_05578_));
 sky130_fd_sc_hd__clkbuf_1 _10782_ (.A(_05578_),
    .X(_00593_));
 sky130_fd_sc_hd__mux2_1 _10783_ (.A0(_05216_),
    .A1(net1953),
    .S(_05577_),
    .X(_05579_));
 sky130_fd_sc_hd__clkbuf_1 _10784_ (.A(_05579_),
    .X(_00594_));
 sky130_fd_sc_hd__mux2_1 _10785_ (.A0(_05218_),
    .A1(net1983),
    .S(_05577_),
    .X(_05580_));
 sky130_fd_sc_hd__clkbuf_1 _10786_ (.A(_05580_),
    .X(_00595_));
 sky130_fd_sc_hd__mux2_1 _10787_ (.A0(_05220_),
    .A1(net2046),
    .S(_05577_),
    .X(_05581_));
 sky130_fd_sc_hd__clkbuf_1 _10788_ (.A(_05581_),
    .X(_00596_));
 sky130_fd_sc_hd__mux2_1 _10789_ (.A0(_05222_),
    .A1(net1920),
    .S(_05577_),
    .X(_05582_));
 sky130_fd_sc_hd__clkbuf_1 _10790_ (.A(_05582_),
    .X(_00597_));
 sky130_fd_sc_hd__mux2_1 _10791_ (.A0(_05224_),
    .A1(net1972),
    .S(_05577_),
    .X(_05583_));
 sky130_fd_sc_hd__clkbuf_1 _10792_ (.A(_05583_),
    .X(_00598_));
 sky130_fd_sc_hd__mux2_1 _10793_ (.A0(_05226_),
    .A1(net1464),
    .S(_05577_),
    .X(_05584_));
 sky130_fd_sc_hd__clkbuf_1 _10794_ (.A(_05584_),
    .X(_00599_));
 sky130_fd_sc_hd__mux2_1 _10795_ (.A0(_05228_),
    .A1(net2038),
    .S(_05577_),
    .X(_05585_));
 sky130_fd_sc_hd__clkbuf_1 _10796_ (.A(_05585_),
    .X(_00600_));
 sky130_fd_sc_hd__mux2_1 _10797_ (.A0(_05230_),
    .A1(net2029),
    .S(_05577_),
    .X(_05586_));
 sky130_fd_sc_hd__clkbuf_1 _10798_ (.A(_05586_),
    .X(_00601_));
 sky130_fd_sc_hd__mux2_1 _10799_ (.A0(_05232_),
    .A1(net1971),
    .S(_05577_),
    .X(_05587_));
 sky130_fd_sc_hd__clkbuf_1 _10800_ (.A(_05587_),
    .X(_00602_));
 sky130_fd_sc_hd__mux2_1 _10801_ (.A0(_05234_),
    .A1(net2026),
    .S(_05576_),
    .X(_05588_));
 sky130_fd_sc_hd__clkbuf_1 _10802_ (.A(_05588_),
    .X(_00603_));
 sky130_fd_sc_hd__mux2_1 _10803_ (.A0(_05236_),
    .A1(net2058),
    .S(_05576_),
    .X(_05589_));
 sky130_fd_sc_hd__clkbuf_1 _10804_ (.A(_05589_),
    .X(_00604_));
 sky130_fd_sc_hd__mux2_1 _10805_ (.A0(_05238_),
    .A1(net2018),
    .S(_05576_),
    .X(_05590_));
 sky130_fd_sc_hd__clkbuf_1 _10806_ (.A(_05590_),
    .X(_00605_));
 sky130_fd_sc_hd__mux2_1 _10807_ (.A0(_05240_),
    .A1(net2076),
    .S(_05576_),
    .X(_05591_));
 sky130_fd_sc_hd__clkbuf_1 _10808_ (.A(_05591_),
    .X(_00606_));
 sky130_fd_sc_hd__mux2_1 _10809_ (.A0(_05242_),
    .A1(net2003),
    .S(_05576_),
    .X(_05592_));
 sky130_fd_sc_hd__clkbuf_1 _10810_ (.A(_05592_),
    .X(_00607_));
 sky130_fd_sc_hd__mux2_1 _10811_ (.A0(_05244_),
    .A1(net1897),
    .S(_05576_),
    .X(_05593_));
 sky130_fd_sc_hd__clkbuf_1 _10812_ (.A(_05593_),
    .X(_00608_));
 sky130_fd_sc_hd__nor2_4 _10813_ (.A(_04186_),
    .B(_04646_),
    .Y(_05594_));
 sky130_fd_sc_hd__buf_4 _10814_ (.A(_05594_),
    .X(_05595_));
 sky130_fd_sc_hd__mux2_1 _10815_ (.A0(net1924),
    .A1(_05469_),
    .S(_05595_),
    .X(_05596_));
 sky130_fd_sc_hd__clkbuf_1 _10816_ (.A(_05596_),
    .X(_00609_));
 sky130_fd_sc_hd__mux2_1 _10817_ (.A0(net355),
    .A1(_05473_),
    .S(_05595_),
    .X(_05597_));
 sky130_fd_sc_hd__clkbuf_1 _10818_ (.A(_05597_),
    .X(_00610_));
 sky130_fd_sc_hd__mux2_1 _10819_ (.A0(net1918),
    .A1(_05475_),
    .S(_05595_),
    .X(_05598_));
 sky130_fd_sc_hd__clkbuf_1 _10820_ (.A(_05598_),
    .X(_00611_));
 sky130_fd_sc_hd__mux2_1 _10821_ (.A0(net1806),
    .A1(_05477_),
    .S(_05595_),
    .X(_05599_));
 sky130_fd_sc_hd__clkbuf_1 _10822_ (.A(_05599_),
    .X(_00612_));
 sky130_fd_sc_hd__mux2_1 _10823_ (.A0(net110),
    .A1(_05479_),
    .S(_05595_),
    .X(_05600_));
 sky130_fd_sc_hd__clkbuf_1 _10824_ (.A(_05600_),
    .X(_00613_));
 sky130_fd_sc_hd__mux2_1 _10825_ (.A0(net679),
    .A1(_05481_),
    .S(_05595_),
    .X(_05601_));
 sky130_fd_sc_hd__clkbuf_1 _10826_ (.A(_05601_),
    .X(_00614_));
 sky130_fd_sc_hd__mux2_1 _10827_ (.A0(net1608),
    .A1(_05483_),
    .S(_05595_),
    .X(_05602_));
 sky130_fd_sc_hd__clkbuf_1 _10828_ (.A(_05602_),
    .X(_00615_));
 sky130_fd_sc_hd__mux2_1 _10829_ (.A0(net230),
    .A1(_05485_),
    .S(_05595_),
    .X(_05603_));
 sky130_fd_sc_hd__clkbuf_1 _10830_ (.A(_05603_),
    .X(_00616_));
 sky130_fd_sc_hd__mux2_1 _10831_ (.A0(net108),
    .A1(_05487_),
    .S(_05595_),
    .X(_05604_));
 sky130_fd_sc_hd__clkbuf_1 _10832_ (.A(_05604_),
    .X(_00617_));
 sky130_fd_sc_hd__mux2_1 _10833_ (.A0(net187),
    .A1(_05489_),
    .S(_05595_),
    .X(_05605_));
 sky130_fd_sc_hd__clkbuf_1 _10834_ (.A(_05605_),
    .X(_00618_));
 sky130_fd_sc_hd__mux2_1 _10835_ (.A0(net1137),
    .A1(_05491_),
    .S(_05594_),
    .X(_05606_));
 sky130_fd_sc_hd__clkbuf_1 _10836_ (.A(_05606_),
    .X(_00619_));
 sky130_fd_sc_hd__mux2_1 _10837_ (.A0(net244),
    .A1(_05493_),
    .S(_05594_),
    .X(_05607_));
 sky130_fd_sc_hd__clkbuf_1 _10838_ (.A(_05607_),
    .X(_00620_));
 sky130_fd_sc_hd__mux2_1 _10839_ (.A0(net162),
    .A1(_05495_),
    .S(_05594_),
    .X(_05608_));
 sky130_fd_sc_hd__clkbuf_1 _10840_ (.A(_05608_),
    .X(_00621_));
 sky130_fd_sc_hd__mux2_1 _10841_ (.A0(net78),
    .A1(_05497_),
    .S(_05594_),
    .X(_05609_));
 sky130_fd_sc_hd__clkbuf_1 _10842_ (.A(_05609_),
    .X(_00622_));
 sky130_fd_sc_hd__mux2_1 _10843_ (.A0(net182),
    .A1(_05499_),
    .S(_05594_),
    .X(_05610_));
 sky130_fd_sc_hd__clkbuf_1 _10844_ (.A(_05610_),
    .X(_00623_));
 sky130_fd_sc_hd__mux2_1 _10845_ (.A0(net157),
    .A1(_05501_),
    .S(_05594_),
    .X(_05611_));
 sky130_fd_sc_hd__clkbuf_1 _10846_ (.A(_05611_),
    .X(_00624_));
 sky130_fd_sc_hd__nor2_4 _10847_ (.A(_04127_),
    .B(_04186_),
    .Y(_05612_));
 sky130_fd_sc_hd__buf_4 _10848_ (.A(_05612_),
    .X(_05613_));
 sky130_fd_sc_hd__mux2_1 _10849_ (.A0(net409),
    .A1(_05469_),
    .S(_05613_),
    .X(_05614_));
 sky130_fd_sc_hd__clkbuf_1 _10850_ (.A(_05614_),
    .X(_00625_));
 sky130_fd_sc_hd__mux2_1 _10851_ (.A0(net1930),
    .A1(_05473_),
    .S(_05613_),
    .X(_05615_));
 sky130_fd_sc_hd__clkbuf_1 _10852_ (.A(_05615_),
    .X(_00626_));
 sky130_fd_sc_hd__mux2_1 _10853_ (.A0(net1243),
    .A1(_05475_),
    .S(_05613_),
    .X(_05616_));
 sky130_fd_sc_hd__clkbuf_1 _10854_ (.A(_05616_),
    .X(_00627_));
 sky130_fd_sc_hd__mux2_1 _10855_ (.A0(net1069),
    .A1(_05477_),
    .S(_05613_),
    .X(_05617_));
 sky130_fd_sc_hd__clkbuf_1 _10856_ (.A(_05617_),
    .X(_00628_));
 sky130_fd_sc_hd__mux2_1 _10857_ (.A0(net1432),
    .A1(_05479_),
    .S(_05613_),
    .X(_05618_));
 sky130_fd_sc_hd__clkbuf_1 _10858_ (.A(_05618_),
    .X(_00629_));
 sky130_fd_sc_hd__mux2_1 _10859_ (.A0(net1232),
    .A1(_05481_),
    .S(_05613_),
    .X(_05619_));
 sky130_fd_sc_hd__clkbuf_1 _10860_ (.A(_05619_),
    .X(_00630_));
 sky130_fd_sc_hd__mux2_1 _10861_ (.A0(net1322),
    .A1(_05483_),
    .S(_05613_),
    .X(_05620_));
 sky130_fd_sc_hd__clkbuf_1 _10862_ (.A(_05620_),
    .X(_00631_));
 sky130_fd_sc_hd__mux2_1 _10863_ (.A0(net418),
    .A1(_05485_),
    .S(_05613_),
    .X(_05621_));
 sky130_fd_sc_hd__clkbuf_1 _10864_ (.A(_05621_),
    .X(_00632_));
 sky130_fd_sc_hd__mux2_1 _10865_ (.A0(net1757),
    .A1(_05487_),
    .S(_05613_),
    .X(_05622_));
 sky130_fd_sc_hd__clkbuf_1 _10866_ (.A(_05622_),
    .X(_00633_));
 sky130_fd_sc_hd__mux2_1 _10867_ (.A0(net762),
    .A1(_05489_),
    .S(_05613_),
    .X(_05623_));
 sky130_fd_sc_hd__clkbuf_1 _10868_ (.A(_05623_),
    .X(_00634_));
 sky130_fd_sc_hd__mux2_1 _10869_ (.A0(net1119),
    .A1(_05491_),
    .S(_05612_),
    .X(_05624_));
 sky130_fd_sc_hd__clkbuf_1 _10870_ (.A(_05624_),
    .X(_00635_));
 sky130_fd_sc_hd__mux2_1 _10871_ (.A0(net903),
    .A1(_05493_),
    .S(_05612_),
    .X(_05625_));
 sky130_fd_sc_hd__clkbuf_1 _10872_ (.A(_05625_),
    .X(_00636_));
 sky130_fd_sc_hd__mux2_1 _10873_ (.A0(net704),
    .A1(_05495_),
    .S(_05612_),
    .X(_05626_));
 sky130_fd_sc_hd__clkbuf_1 _10874_ (.A(_05626_),
    .X(_00637_));
 sky130_fd_sc_hd__mux2_1 _10875_ (.A0(net594),
    .A1(_05497_),
    .S(_05612_),
    .X(_05627_));
 sky130_fd_sc_hd__clkbuf_1 _10876_ (.A(_05627_),
    .X(_00638_));
 sky130_fd_sc_hd__mux2_1 _10877_ (.A0(net708),
    .A1(_05499_),
    .S(_05612_),
    .X(_05628_));
 sky130_fd_sc_hd__clkbuf_1 _10878_ (.A(_05628_),
    .X(_00639_));
 sky130_fd_sc_hd__mux2_1 _10879_ (.A0(net1074),
    .A1(_05501_),
    .S(_05612_),
    .X(_05629_));
 sky130_fd_sc_hd__clkbuf_1 _10880_ (.A(_05629_),
    .X(_00640_));
 sky130_fd_sc_hd__nor2_4 _10881_ (.A(_04186_),
    .B(_04684_),
    .Y(_05630_));
 sky130_fd_sc_hd__buf_4 _10882_ (.A(_05630_),
    .X(_05631_));
 sky130_fd_sc_hd__mux2_1 _10883_ (.A0(net171),
    .A1(_05469_),
    .S(_05631_),
    .X(_05632_));
 sky130_fd_sc_hd__clkbuf_1 _10884_ (.A(_05632_),
    .X(_00641_));
 sky130_fd_sc_hd__mux2_1 _10885_ (.A0(net1328),
    .A1(_05473_),
    .S(_05631_),
    .X(_05633_));
 sky130_fd_sc_hd__clkbuf_1 _10886_ (.A(_05633_),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _10887_ (.A0(net327),
    .A1(_05475_),
    .S(_05631_),
    .X(_05634_));
 sky130_fd_sc_hd__clkbuf_1 _10888_ (.A(_05634_),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _10889_ (.A0(net242),
    .A1(_05477_),
    .S(_05631_),
    .X(_05635_));
 sky130_fd_sc_hd__clkbuf_1 _10890_ (.A(_05635_),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _10891_ (.A0(net525),
    .A1(_05479_),
    .S(_05631_),
    .X(_05636_));
 sky130_fd_sc_hd__clkbuf_1 _10892_ (.A(_05636_),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_1 _10893_ (.A0(net781),
    .A1(_05481_),
    .S(_05631_),
    .X(_05637_));
 sky130_fd_sc_hd__clkbuf_1 _10894_ (.A(_05637_),
    .X(_00646_));
 sky130_fd_sc_hd__mux2_1 _10895_ (.A0(net260),
    .A1(_05483_),
    .S(_05631_),
    .X(_05638_));
 sky130_fd_sc_hd__clkbuf_1 _10896_ (.A(_05638_),
    .X(_00647_));
 sky130_fd_sc_hd__mux2_1 _10897_ (.A0(net1044),
    .A1(_05485_),
    .S(_05631_),
    .X(_05639_));
 sky130_fd_sc_hd__clkbuf_1 _10898_ (.A(_05639_),
    .X(_00648_));
 sky130_fd_sc_hd__mux2_1 _10899_ (.A0(net1078),
    .A1(_05487_),
    .S(_05631_),
    .X(_05640_));
 sky130_fd_sc_hd__clkbuf_1 _10900_ (.A(_05640_),
    .X(_00649_));
 sky130_fd_sc_hd__mux2_1 _10901_ (.A0(net1217),
    .A1(_05489_),
    .S(_05631_),
    .X(_05641_));
 sky130_fd_sc_hd__clkbuf_1 _10902_ (.A(_05641_),
    .X(_00650_));
 sky130_fd_sc_hd__mux2_1 _10903_ (.A0(net109),
    .A1(_05491_),
    .S(_05630_),
    .X(_05642_));
 sky130_fd_sc_hd__clkbuf_1 _10904_ (.A(_05642_),
    .X(_00651_));
 sky130_fd_sc_hd__mux2_1 _10905_ (.A0(net189),
    .A1(_05493_),
    .S(_05630_),
    .X(_05643_));
 sky130_fd_sc_hd__clkbuf_1 _10906_ (.A(_05643_),
    .X(_00652_));
 sky130_fd_sc_hd__mux2_1 _10907_ (.A0(net821),
    .A1(_05495_),
    .S(_05630_),
    .X(_05644_));
 sky130_fd_sc_hd__clkbuf_1 _10908_ (.A(_05644_),
    .X(_00653_));
 sky130_fd_sc_hd__mux2_1 _10909_ (.A0(net668),
    .A1(_05497_),
    .S(_05630_),
    .X(_05645_));
 sky130_fd_sc_hd__clkbuf_1 _10910_ (.A(_05645_),
    .X(_00654_));
 sky130_fd_sc_hd__mux2_1 _10911_ (.A0(net120),
    .A1(_05499_),
    .S(_05630_),
    .X(_05646_));
 sky130_fd_sc_hd__clkbuf_1 _10912_ (.A(_05646_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _10913_ (.A0(net177),
    .A1(_05501_),
    .S(_05630_),
    .X(_05647_));
 sky130_fd_sc_hd__clkbuf_1 _10914_ (.A(_05647_),
    .X(_00656_));
 sky130_fd_sc_hd__buf_6 _10915_ (.A(_04069_),
    .X(_05648_));
 sky130_fd_sc_hd__or3_1 _10916_ (.A(_02707_),
    .B(_05026_),
    .C(_04185_),
    .X(_05649_));
 sky130_fd_sc_hd__clkbuf_4 _10917_ (.A(_05649_),
    .X(_05650_));
 sky130_fd_sc_hd__buf_4 _10918_ (.A(_05650_),
    .X(_05651_));
 sky130_fd_sc_hd__mux2_1 _10919_ (.A0(_05648_),
    .A1(net1657),
    .S(_05651_),
    .X(_05652_));
 sky130_fd_sc_hd__clkbuf_1 _10920_ (.A(_05652_),
    .X(_00657_));
 sky130_fd_sc_hd__clkbuf_4 _10921_ (.A(_04080_),
    .X(_05653_));
 sky130_fd_sc_hd__mux2_1 _10922_ (.A0(_05653_),
    .A1(net2019),
    .S(_05651_),
    .X(_05654_));
 sky130_fd_sc_hd__clkbuf_1 _10923_ (.A(_05654_),
    .X(_00658_));
 sky130_fd_sc_hd__buf_6 _10924_ (.A(_04083_),
    .X(_05655_));
 sky130_fd_sc_hd__mux2_1 _10925_ (.A0(_05655_),
    .A1(net1820),
    .S(_05651_),
    .X(_05656_));
 sky130_fd_sc_hd__clkbuf_1 _10926_ (.A(_05656_),
    .X(_00659_));
 sky130_fd_sc_hd__buf_6 _10927_ (.A(_04086_),
    .X(_05657_));
 sky130_fd_sc_hd__mux2_1 _10928_ (.A0(_05657_),
    .A1(net1903),
    .S(_05651_),
    .X(_05658_));
 sky130_fd_sc_hd__clkbuf_1 _10929_ (.A(_05658_),
    .X(_00660_));
 sky130_fd_sc_hd__buf_4 _10930_ (.A(_04089_),
    .X(_05659_));
 sky130_fd_sc_hd__mux2_1 _10931_ (.A0(_05659_),
    .A1(net1754),
    .S(_05651_),
    .X(_05660_));
 sky130_fd_sc_hd__clkbuf_1 _10932_ (.A(_05660_),
    .X(_00661_));
 sky130_fd_sc_hd__buf_4 _10933_ (.A(_04092_),
    .X(_05661_));
 sky130_fd_sc_hd__mux2_1 _10934_ (.A0(_05661_),
    .A1(net2042),
    .S(_05651_),
    .X(_05662_));
 sky130_fd_sc_hd__clkbuf_1 _10935_ (.A(_05662_),
    .X(_00662_));
 sky130_fd_sc_hd__buf_4 _10936_ (.A(_04095_),
    .X(_05663_));
 sky130_fd_sc_hd__mux2_1 _10937_ (.A0(_05663_),
    .A1(net1993),
    .S(_05651_),
    .X(_05664_));
 sky130_fd_sc_hd__clkbuf_1 _10938_ (.A(_05664_),
    .X(_00663_));
 sky130_fd_sc_hd__buf_4 _10939_ (.A(_04098_),
    .X(_05665_));
 sky130_fd_sc_hd__mux2_1 _10940_ (.A0(_05665_),
    .A1(net1458),
    .S(_05651_),
    .X(_05666_));
 sky130_fd_sc_hd__clkbuf_1 _10941_ (.A(_05666_),
    .X(_00664_));
 sky130_fd_sc_hd__buf_4 _10942_ (.A(_04101_),
    .X(_05667_));
 sky130_fd_sc_hd__mux2_1 _10943_ (.A0(_05667_),
    .A1(net1416),
    .S(_05651_),
    .X(_05668_));
 sky130_fd_sc_hd__clkbuf_1 _10944_ (.A(_05668_),
    .X(_00665_));
 sky130_fd_sc_hd__buf_4 _10945_ (.A(_04104_),
    .X(_05669_));
 sky130_fd_sc_hd__mux2_1 _10946_ (.A0(_05669_),
    .A1(net1941),
    .S(_05651_),
    .X(_05670_));
 sky130_fd_sc_hd__clkbuf_1 _10947_ (.A(_05670_),
    .X(_00666_));
 sky130_fd_sc_hd__buf_4 _10948_ (.A(_04107_),
    .X(_05671_));
 sky130_fd_sc_hd__mux2_1 _10949_ (.A0(_05671_),
    .A1(net1505),
    .S(_05650_),
    .X(_05672_));
 sky130_fd_sc_hd__clkbuf_1 _10950_ (.A(_05672_),
    .X(_00667_));
 sky130_fd_sc_hd__clkbuf_4 _10951_ (.A(_04110_),
    .X(_05673_));
 sky130_fd_sc_hd__mux2_1 _10952_ (.A0(_05673_),
    .A1(net1808),
    .S(_05650_),
    .X(_05674_));
 sky130_fd_sc_hd__clkbuf_1 _10953_ (.A(_05674_),
    .X(_00668_));
 sky130_fd_sc_hd__buf_4 _10954_ (.A(_04113_),
    .X(_05675_));
 sky130_fd_sc_hd__mux2_1 _10955_ (.A0(_05675_),
    .A1(net1859),
    .S(_05650_),
    .X(_05676_));
 sky130_fd_sc_hd__clkbuf_1 _10956_ (.A(_05676_),
    .X(_00669_));
 sky130_fd_sc_hd__clkbuf_4 _10957_ (.A(_04116_),
    .X(_05677_));
 sky130_fd_sc_hd__mux2_1 _10958_ (.A0(_05677_),
    .A1(net1875),
    .S(_05650_),
    .X(_05678_));
 sky130_fd_sc_hd__clkbuf_1 _10959_ (.A(_05678_),
    .X(_00670_));
 sky130_fd_sc_hd__buf_4 _10960_ (.A(_04119_),
    .X(_05679_));
 sky130_fd_sc_hd__mux2_1 _10961_ (.A0(_05679_),
    .A1(net1736),
    .S(_05650_),
    .X(_05680_));
 sky130_fd_sc_hd__clkbuf_1 _10962_ (.A(_05680_),
    .X(_00671_));
 sky130_fd_sc_hd__buf_4 _10963_ (.A(_04122_),
    .X(_05681_));
 sky130_fd_sc_hd__mux2_1 _10964_ (.A0(_05681_),
    .A1(net1632),
    .S(_05650_),
    .X(_05682_));
 sky130_fd_sc_hd__clkbuf_1 _10965_ (.A(_05682_),
    .X(_00672_));
 sky130_fd_sc_hd__nor2_4 _10966_ (.A(_04185_),
    .B(_04365_),
    .Y(_05683_));
 sky130_fd_sc_hd__buf_4 _10967_ (.A(_05683_),
    .X(_05684_));
 sky130_fd_sc_hd__mux2_1 _10968_ (.A0(net665),
    .A1(_05469_),
    .S(_05684_),
    .X(_05685_));
 sky130_fd_sc_hd__clkbuf_1 _10969_ (.A(_05685_),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_1 _10970_ (.A0(net1211),
    .A1(_05473_),
    .S(_05684_),
    .X(_05686_));
 sky130_fd_sc_hd__clkbuf_1 _10971_ (.A(_05686_),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_1 _10972_ (.A0(net1046),
    .A1(_05475_),
    .S(_05684_),
    .X(_05687_));
 sky130_fd_sc_hd__clkbuf_1 _10973_ (.A(_05687_),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_1 _10974_ (.A0(net422),
    .A1(_05477_),
    .S(_05684_),
    .X(_05688_));
 sky130_fd_sc_hd__clkbuf_1 _10975_ (.A(_05688_),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _10976_ (.A0(net138),
    .A1(_05479_),
    .S(_05684_),
    .X(_05689_));
 sky130_fd_sc_hd__clkbuf_1 _10977_ (.A(_05689_),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _10978_ (.A0(net49),
    .A1(_05481_),
    .S(_05684_),
    .X(_05690_));
 sky130_fd_sc_hd__clkbuf_1 _10979_ (.A(_05690_),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_1 _10980_ (.A0(net373),
    .A1(_05483_),
    .S(_05684_),
    .X(_05691_));
 sky130_fd_sc_hd__clkbuf_1 _10981_ (.A(_05691_),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _10982_ (.A0(net107),
    .A1(_05485_),
    .S(_05684_),
    .X(_05692_));
 sky130_fd_sc_hd__clkbuf_1 _10983_ (.A(_05692_),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_1 _10984_ (.A0(net65),
    .A1(_05487_),
    .S(_05684_),
    .X(_05693_));
 sky130_fd_sc_hd__clkbuf_1 _10985_ (.A(_05693_),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_1 _10986_ (.A0(net91),
    .A1(_05489_),
    .S(_05684_),
    .X(_05694_));
 sky130_fd_sc_hd__clkbuf_1 _10987_ (.A(_05694_),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _10988_ (.A0(net190),
    .A1(_05491_),
    .S(_05683_),
    .X(_05695_));
 sky130_fd_sc_hd__clkbuf_1 _10989_ (.A(_05695_),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _10990_ (.A0(net85),
    .A1(_05493_),
    .S(_05683_),
    .X(_05696_));
 sky130_fd_sc_hd__clkbuf_1 _10991_ (.A(_05696_),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_1 _10992_ (.A0(net105),
    .A1(_05495_),
    .S(_05683_),
    .X(_05697_));
 sky130_fd_sc_hd__clkbuf_1 _10993_ (.A(_05697_),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _10994_ (.A0(net166),
    .A1(_05497_),
    .S(_05683_),
    .X(_05698_));
 sky130_fd_sc_hd__clkbuf_1 _10995_ (.A(_05698_),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_1 _10996_ (.A0(net450),
    .A1(_05499_),
    .S(_05683_),
    .X(_05699_));
 sky130_fd_sc_hd__clkbuf_1 _10997_ (.A(_05699_),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _10998_ (.A0(net67),
    .A1(_05501_),
    .S(_05683_),
    .X(_05700_));
 sky130_fd_sc_hd__clkbuf_1 _10999_ (.A(_05700_),
    .X(_00688_));
 sky130_fd_sc_hd__or3_1 _11000_ (.A(_02484_),
    .B(_02737_),
    .C(_04185_),
    .X(_05701_));
 sky130_fd_sc_hd__buf_2 _11001_ (.A(_05701_),
    .X(_05702_));
 sky130_fd_sc_hd__buf_4 _11002_ (.A(_05702_),
    .X(_05703_));
 sky130_fd_sc_hd__mux2_1 _11003_ (.A0(_05648_),
    .A1(net1743),
    .S(_05703_),
    .X(_05704_));
 sky130_fd_sc_hd__clkbuf_1 _11004_ (.A(_05704_),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _11005_ (.A0(_05653_),
    .A1(net1686),
    .S(_05703_),
    .X(_05705_));
 sky130_fd_sc_hd__clkbuf_1 _11006_ (.A(_05705_),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _11007_ (.A0(_05655_),
    .A1(net1155),
    .S(_05703_),
    .X(_05706_));
 sky130_fd_sc_hd__clkbuf_1 _11008_ (.A(_05706_),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _11009_ (.A0(_05657_),
    .A1(net1536),
    .S(_05703_),
    .X(_05707_));
 sky130_fd_sc_hd__clkbuf_1 _11010_ (.A(_05707_),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _11011_ (.A0(_05659_),
    .A1(net1870),
    .S(_05703_),
    .X(_05708_));
 sky130_fd_sc_hd__clkbuf_1 _11012_ (.A(_05708_),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _11013_ (.A0(_05661_),
    .A1(net1428),
    .S(_05703_),
    .X(_05709_));
 sky130_fd_sc_hd__clkbuf_1 _11014_ (.A(_05709_),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_1 _11015_ (.A0(_05663_),
    .A1(net1033),
    .S(_05703_),
    .X(_05710_));
 sky130_fd_sc_hd__clkbuf_1 _11016_ (.A(_05710_),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _11017_ (.A0(_05665_),
    .A1(net1977),
    .S(_05703_),
    .X(_05711_));
 sky130_fd_sc_hd__clkbuf_1 _11018_ (.A(_05711_),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _11019_ (.A0(_05667_),
    .A1(net1728),
    .S(_05703_),
    .X(_05712_));
 sky130_fd_sc_hd__clkbuf_1 _11020_ (.A(_05712_),
    .X(_00697_));
 sky130_fd_sc_hd__mux2_1 _11021_ (.A0(_05669_),
    .A1(net783),
    .S(_05703_),
    .X(_05713_));
 sky130_fd_sc_hd__clkbuf_1 _11022_ (.A(_05713_),
    .X(_00698_));
 sky130_fd_sc_hd__mux2_1 _11023_ (.A0(_05671_),
    .A1(net1815),
    .S(_05702_),
    .X(_05714_));
 sky130_fd_sc_hd__clkbuf_1 _11024_ (.A(_05714_),
    .X(_00699_));
 sky130_fd_sc_hd__mux2_1 _11025_ (.A0(_05673_),
    .A1(net1619),
    .S(_05702_),
    .X(_05715_));
 sky130_fd_sc_hd__clkbuf_1 _11026_ (.A(_05715_),
    .X(_00700_));
 sky130_fd_sc_hd__mux2_1 _11027_ (.A0(_05675_),
    .A1(net1270),
    .S(_05702_),
    .X(_05716_));
 sky130_fd_sc_hd__clkbuf_1 _11028_ (.A(_05716_),
    .X(_00701_));
 sky130_fd_sc_hd__mux2_1 _11029_ (.A0(_05677_),
    .A1(net939),
    .S(_05702_),
    .X(_05717_));
 sky130_fd_sc_hd__clkbuf_1 _11030_ (.A(_05717_),
    .X(_00702_));
 sky130_fd_sc_hd__mux2_1 _11031_ (.A0(_05679_),
    .A1(net1618),
    .S(_05702_),
    .X(_05718_));
 sky130_fd_sc_hd__clkbuf_1 _11032_ (.A(_05718_),
    .X(_00703_));
 sky130_fd_sc_hd__mux2_1 _11033_ (.A0(_05681_),
    .A1(net838),
    .S(_05702_),
    .X(_05719_));
 sky130_fd_sc_hd__clkbuf_1 _11034_ (.A(_05719_),
    .X(_00704_));
 sky130_fd_sc_hd__nand2b_4 _11035_ (.A_N(_04185_),
    .B(_04408_),
    .Y(_05720_));
 sky130_fd_sc_hd__buf_4 _11036_ (.A(_05720_),
    .X(_05721_));
 sky130_fd_sc_hd__mux2_1 _11037_ (.A0(_05648_),
    .A1(net2033),
    .S(_05721_),
    .X(_05722_));
 sky130_fd_sc_hd__clkbuf_1 _11038_ (.A(_05722_),
    .X(_00705_));
 sky130_fd_sc_hd__mux2_1 _11039_ (.A0(_05653_),
    .A1(net1599),
    .S(_05721_),
    .X(_05723_));
 sky130_fd_sc_hd__clkbuf_1 _11040_ (.A(_05723_),
    .X(_00706_));
 sky130_fd_sc_hd__mux2_1 _11041_ (.A0(_05655_),
    .A1(net2004),
    .S(_05721_),
    .X(_05724_));
 sky130_fd_sc_hd__clkbuf_1 _11042_ (.A(_05724_),
    .X(_00707_));
 sky130_fd_sc_hd__mux2_1 _11043_ (.A0(_05657_),
    .A1(net2036),
    .S(_05721_),
    .X(_05725_));
 sky130_fd_sc_hd__clkbuf_1 _11044_ (.A(_05725_),
    .X(_00708_));
 sky130_fd_sc_hd__mux2_1 _11045_ (.A0(_05659_),
    .A1(net1922),
    .S(_05721_),
    .X(_05726_));
 sky130_fd_sc_hd__clkbuf_1 _11046_ (.A(_05726_),
    .X(_00709_));
 sky130_fd_sc_hd__mux2_1 _11047_ (.A0(_05661_),
    .A1(net1494),
    .S(_05721_),
    .X(_05727_));
 sky130_fd_sc_hd__clkbuf_1 _11048_ (.A(_05727_),
    .X(_00710_));
 sky130_fd_sc_hd__mux2_1 _11049_ (.A0(_05663_),
    .A1(net1622),
    .S(_05721_),
    .X(_05728_));
 sky130_fd_sc_hd__clkbuf_1 _11050_ (.A(_05728_),
    .X(_00711_));
 sky130_fd_sc_hd__mux2_1 _11051_ (.A0(_05665_),
    .A1(net1965),
    .S(_05721_),
    .X(_05729_));
 sky130_fd_sc_hd__clkbuf_1 _11052_ (.A(_05729_),
    .X(_00712_));
 sky130_fd_sc_hd__mux2_1 _11053_ (.A0(_05667_),
    .A1(net1829),
    .S(_05721_),
    .X(_05730_));
 sky130_fd_sc_hd__clkbuf_1 _11054_ (.A(_05730_),
    .X(_00713_));
 sky130_fd_sc_hd__mux2_1 _11055_ (.A0(_05669_),
    .A1(net1837),
    .S(_05721_),
    .X(_05731_));
 sky130_fd_sc_hd__clkbuf_1 _11056_ (.A(_05731_),
    .X(_00714_));
 sky130_fd_sc_hd__mux2_1 _11057_ (.A0(_05671_),
    .A1(net1876),
    .S(_05720_),
    .X(_05732_));
 sky130_fd_sc_hd__clkbuf_1 _11058_ (.A(_05732_),
    .X(_00715_));
 sky130_fd_sc_hd__mux2_1 _11059_ (.A0(_05673_),
    .A1(net1490),
    .S(_05720_),
    .X(_05733_));
 sky130_fd_sc_hd__clkbuf_1 _11060_ (.A(_05733_),
    .X(_00716_));
 sky130_fd_sc_hd__mux2_1 _11061_ (.A0(_05675_),
    .A1(net1275),
    .S(_05720_),
    .X(_05734_));
 sky130_fd_sc_hd__clkbuf_1 _11062_ (.A(_05734_),
    .X(_00717_));
 sky130_fd_sc_hd__mux2_1 _11063_ (.A0(_05677_),
    .A1(net1772),
    .S(_05720_),
    .X(_05735_));
 sky130_fd_sc_hd__clkbuf_1 _11064_ (.A(_05735_),
    .X(_00718_));
 sky130_fd_sc_hd__mux2_1 _11065_ (.A0(_05679_),
    .A1(net1811),
    .S(_05720_),
    .X(_05736_));
 sky130_fd_sc_hd__clkbuf_1 _11066_ (.A(_05736_),
    .X(_00719_));
 sky130_fd_sc_hd__mux2_1 _11067_ (.A0(_05681_),
    .A1(net1277),
    .S(_05720_),
    .X(_05737_));
 sky130_fd_sc_hd__clkbuf_1 _11068_ (.A(_05737_),
    .X(_00720_));
 sky130_fd_sc_hd__or3_1 _11069_ (.A(_02498_),
    .B(_05026_),
    .C(_04367_),
    .X(_05738_));
 sky130_fd_sc_hd__clkbuf_4 _11070_ (.A(_05738_),
    .X(_05739_));
 sky130_fd_sc_hd__buf_4 _11071_ (.A(_05739_),
    .X(_05740_));
 sky130_fd_sc_hd__mux2_1 _11072_ (.A0(_05648_),
    .A1(net1989),
    .S(_05740_),
    .X(_05741_));
 sky130_fd_sc_hd__clkbuf_1 _11073_ (.A(_05741_),
    .X(_00721_));
 sky130_fd_sc_hd__mux2_1 _11074_ (.A0(_05653_),
    .A1(net1803),
    .S(_05740_),
    .X(_05742_));
 sky130_fd_sc_hd__clkbuf_1 _11075_ (.A(_05742_),
    .X(_00722_));
 sky130_fd_sc_hd__mux2_1 _11076_ (.A0(_05655_),
    .A1(net1565),
    .S(_05740_),
    .X(_05743_));
 sky130_fd_sc_hd__clkbuf_1 _11077_ (.A(_05743_),
    .X(_00723_));
 sky130_fd_sc_hd__mux2_1 _11078_ (.A0(_05657_),
    .A1(net1150),
    .S(_05740_),
    .X(_05744_));
 sky130_fd_sc_hd__clkbuf_1 _11079_ (.A(_05744_),
    .X(_00724_));
 sky130_fd_sc_hd__mux2_1 _11080_ (.A0(_05659_),
    .A1(net1334),
    .S(_05740_),
    .X(_05745_));
 sky130_fd_sc_hd__clkbuf_1 _11081_ (.A(_05745_),
    .X(_00725_));
 sky130_fd_sc_hd__mux2_1 _11082_ (.A0(_05661_),
    .A1(net2049),
    .S(_05740_),
    .X(_05746_));
 sky130_fd_sc_hd__clkbuf_1 _11083_ (.A(_05746_),
    .X(_00726_));
 sky130_fd_sc_hd__mux2_1 _11084_ (.A0(_05663_),
    .A1(net1507),
    .S(_05740_),
    .X(_05747_));
 sky130_fd_sc_hd__clkbuf_1 _11085_ (.A(_05747_),
    .X(_00727_));
 sky130_fd_sc_hd__mux2_1 _11086_ (.A0(_05665_),
    .A1(net1886),
    .S(_05740_),
    .X(_05748_));
 sky130_fd_sc_hd__clkbuf_1 _11087_ (.A(_05748_),
    .X(_00728_));
 sky130_fd_sc_hd__mux2_1 _11088_ (.A0(_05667_),
    .A1(net2025),
    .S(_05740_),
    .X(_05749_));
 sky130_fd_sc_hd__clkbuf_1 _11089_ (.A(_05749_),
    .X(_00729_));
 sky130_fd_sc_hd__mux2_1 _11090_ (.A0(_05669_),
    .A1(net1904),
    .S(_05740_),
    .X(_05750_));
 sky130_fd_sc_hd__clkbuf_1 _11091_ (.A(_05750_),
    .X(_00730_));
 sky130_fd_sc_hd__mux2_1 _11092_ (.A0(_05671_),
    .A1(net1928),
    .S(_05739_),
    .X(_05751_));
 sky130_fd_sc_hd__clkbuf_1 _11093_ (.A(_05751_),
    .X(_00731_));
 sky130_fd_sc_hd__mux2_1 _11094_ (.A0(_05673_),
    .A1(net1838),
    .S(_05739_),
    .X(_05752_));
 sky130_fd_sc_hd__clkbuf_1 _11095_ (.A(_05752_),
    .X(_00732_));
 sky130_fd_sc_hd__mux2_1 _11096_ (.A0(_05675_),
    .A1(net1640),
    .S(_05739_),
    .X(_05753_));
 sky130_fd_sc_hd__clkbuf_1 _11097_ (.A(_05753_),
    .X(_00733_));
 sky130_fd_sc_hd__mux2_1 _11098_ (.A0(_05677_),
    .A1(net949),
    .S(_05739_),
    .X(_05754_));
 sky130_fd_sc_hd__clkbuf_1 _11099_ (.A(_05754_),
    .X(_00734_));
 sky130_fd_sc_hd__mux2_1 _11100_ (.A0(_05679_),
    .A1(net1175),
    .S(_05739_),
    .X(_05755_));
 sky130_fd_sc_hd__clkbuf_1 _11101_ (.A(_05755_),
    .X(_00735_));
 sky130_fd_sc_hd__mux2_1 _11102_ (.A0(_05681_),
    .A1(net1641),
    .S(_05739_),
    .X(_05756_));
 sky130_fd_sc_hd__clkbuf_1 _11103_ (.A(_05756_),
    .X(_00736_));
 sky130_fd_sc_hd__buf_4 _11104_ (.A(_04129_),
    .X(_05757_));
 sky130_fd_sc_hd__nor2_4 _11105_ (.A(_05757_),
    .B(_04461_),
    .Y(_05758_));
 sky130_fd_sc_hd__buf_4 _11106_ (.A(_05758_),
    .X(_05759_));
 sky130_fd_sc_hd__mux2_1 _11107_ (.A0(net1209),
    .A1(_05469_),
    .S(_05759_),
    .X(_05760_));
 sky130_fd_sc_hd__clkbuf_1 _11108_ (.A(_05760_),
    .X(_00737_));
 sky130_fd_sc_hd__mux2_1 _11109_ (.A0(net1952),
    .A1(_05473_),
    .S(_05759_),
    .X(_05761_));
 sky130_fd_sc_hd__clkbuf_1 _11110_ (.A(_05761_),
    .X(_00738_));
 sky130_fd_sc_hd__mux2_1 _11111_ (.A0(net1908),
    .A1(_05475_),
    .S(_05759_),
    .X(_05762_));
 sky130_fd_sc_hd__clkbuf_1 _11112_ (.A(_05762_),
    .X(_00739_));
 sky130_fd_sc_hd__mux2_1 _11113_ (.A0(net1153),
    .A1(_05477_),
    .S(_05759_),
    .X(_05763_));
 sky130_fd_sc_hd__clkbuf_1 _11114_ (.A(_05763_),
    .X(_00740_));
 sky130_fd_sc_hd__mux2_1 _11115_ (.A0(net1580),
    .A1(_05479_),
    .S(_05759_),
    .X(_05764_));
 sky130_fd_sc_hd__clkbuf_1 _11116_ (.A(_05764_),
    .X(_00741_));
 sky130_fd_sc_hd__mux2_1 _11117_ (.A0(net929),
    .A1(_05481_),
    .S(_05759_),
    .X(_05765_));
 sky130_fd_sc_hd__clkbuf_1 _11118_ (.A(_05765_),
    .X(_00742_));
 sky130_fd_sc_hd__mux2_1 _11119_ (.A0(net2057),
    .A1(_05483_),
    .S(_05759_),
    .X(_05766_));
 sky130_fd_sc_hd__clkbuf_1 _11120_ (.A(_05766_),
    .X(_00743_));
 sky130_fd_sc_hd__mux2_1 _11121_ (.A0(net1606),
    .A1(_05485_),
    .S(_05759_),
    .X(_05767_));
 sky130_fd_sc_hd__clkbuf_1 _11122_ (.A(_05767_),
    .X(_00744_));
 sky130_fd_sc_hd__mux2_1 _11123_ (.A0(net1961),
    .A1(_05487_),
    .S(_05759_),
    .X(_05768_));
 sky130_fd_sc_hd__clkbuf_1 _11124_ (.A(_05768_),
    .X(_00745_));
 sky130_fd_sc_hd__mux2_1 _11125_ (.A0(net1447),
    .A1(_05489_),
    .S(_05759_),
    .X(_05769_));
 sky130_fd_sc_hd__clkbuf_1 _11126_ (.A(_05769_),
    .X(_00746_));
 sky130_fd_sc_hd__mux2_1 _11127_ (.A0(net2067),
    .A1(_05491_),
    .S(_05758_),
    .X(_05770_));
 sky130_fd_sc_hd__clkbuf_1 _11128_ (.A(_05770_),
    .X(_00747_));
 sky130_fd_sc_hd__mux2_1 _11129_ (.A0(net2039),
    .A1(_05493_),
    .S(_05758_),
    .X(_05771_));
 sky130_fd_sc_hd__clkbuf_1 _11130_ (.A(_05771_),
    .X(_00748_));
 sky130_fd_sc_hd__mux2_1 _11131_ (.A0(net2075),
    .A1(_05495_),
    .S(_05758_),
    .X(_05772_));
 sky130_fd_sc_hd__clkbuf_1 _11132_ (.A(_05772_),
    .X(_00749_));
 sky130_fd_sc_hd__mux2_1 _11133_ (.A0(net1650),
    .A1(_05497_),
    .S(_05758_),
    .X(_05773_));
 sky130_fd_sc_hd__clkbuf_1 _11134_ (.A(_05773_),
    .X(_00750_));
 sky130_fd_sc_hd__mux2_1 _11135_ (.A0(net2068),
    .A1(_05499_),
    .S(_05758_),
    .X(_05774_));
 sky130_fd_sc_hd__clkbuf_1 _11136_ (.A(_05774_),
    .X(_00751_));
 sky130_fd_sc_hd__mux2_1 _11137_ (.A0(net578),
    .A1(_05501_),
    .S(_05758_),
    .X(_05775_));
 sky130_fd_sc_hd__clkbuf_1 _11138_ (.A(_05775_),
    .X(_00752_));
 sky130_fd_sc_hd__buf_8 _11139_ (.A(_04069_),
    .X(_05776_));
 sky130_fd_sc_hd__nor2_4 _11140_ (.A(_04072_),
    .B(_05757_),
    .Y(_05777_));
 sky130_fd_sc_hd__buf_4 _11141_ (.A(_05777_),
    .X(_05778_));
 sky130_fd_sc_hd__mux2_1 _11142_ (.A0(net865),
    .A1(_05776_),
    .S(_05778_),
    .X(_05779_));
 sky130_fd_sc_hd__clkbuf_1 _11143_ (.A(_05779_),
    .X(_00753_));
 sky130_fd_sc_hd__buf_6 _11144_ (.A(_04080_),
    .X(_05780_));
 sky130_fd_sc_hd__mux2_1 _11145_ (.A0(net458),
    .A1(_05780_),
    .S(_05778_),
    .X(_05781_));
 sky130_fd_sc_hd__clkbuf_1 _11146_ (.A(_05781_),
    .X(_00754_));
 sky130_fd_sc_hd__clkbuf_16 _11147_ (.A(_04083_),
    .X(_05782_));
 sky130_fd_sc_hd__mux2_1 _11148_ (.A0(net1117),
    .A1(_05782_),
    .S(_05778_),
    .X(_05783_));
 sky130_fd_sc_hd__clkbuf_1 _11149_ (.A(_05783_),
    .X(_00755_));
 sky130_fd_sc_hd__clkbuf_16 _11150_ (.A(_04086_),
    .X(_05784_));
 sky130_fd_sc_hd__mux2_1 _11151_ (.A0(net1484),
    .A1(_05784_),
    .S(_05778_),
    .X(_05785_));
 sky130_fd_sc_hd__clkbuf_1 _11152_ (.A(_05785_),
    .X(_00756_));
 sky130_fd_sc_hd__buf_8 _11153_ (.A(_04089_),
    .X(_05786_));
 sky130_fd_sc_hd__mux2_1 _11154_ (.A0(net844),
    .A1(_05786_),
    .S(_05778_),
    .X(_05787_));
 sky130_fd_sc_hd__clkbuf_1 _11155_ (.A(_05787_),
    .X(_00757_));
 sky130_fd_sc_hd__buf_6 _11156_ (.A(_04092_),
    .X(_05788_));
 sky130_fd_sc_hd__mux2_1 _11157_ (.A0(net1551),
    .A1(_05788_),
    .S(_05778_),
    .X(_05789_));
 sky130_fd_sc_hd__clkbuf_1 _11158_ (.A(_05789_),
    .X(_00758_));
 sky130_fd_sc_hd__buf_6 _11159_ (.A(_04095_),
    .X(_05790_));
 sky130_fd_sc_hd__mux2_1 _11160_ (.A0(net1691),
    .A1(_05790_),
    .S(_05778_),
    .X(_05791_));
 sky130_fd_sc_hd__clkbuf_1 _11161_ (.A(_05791_),
    .X(_00759_));
 sky130_fd_sc_hd__buf_8 _11162_ (.A(_04098_),
    .X(_05792_));
 sky130_fd_sc_hd__mux2_1 _11163_ (.A0(net694),
    .A1(_05792_),
    .S(_05778_),
    .X(_05793_));
 sky130_fd_sc_hd__clkbuf_1 _11164_ (.A(_05793_),
    .X(_00760_));
 sky130_fd_sc_hd__buf_8 _11165_ (.A(_04101_),
    .X(_05794_));
 sky130_fd_sc_hd__mux2_1 _11166_ (.A0(net636),
    .A1(_05794_),
    .S(_05778_),
    .X(_05795_));
 sky130_fd_sc_hd__clkbuf_1 _11167_ (.A(_05795_),
    .X(_00761_));
 sky130_fd_sc_hd__buf_8 _11168_ (.A(_04104_),
    .X(_05796_));
 sky130_fd_sc_hd__mux2_1 _11169_ (.A0(net1307),
    .A1(_05796_),
    .S(_05778_),
    .X(_05797_));
 sky130_fd_sc_hd__clkbuf_1 _11170_ (.A(_05797_),
    .X(_00762_));
 sky130_fd_sc_hd__buf_6 _11171_ (.A(_04107_),
    .X(_05798_));
 sky130_fd_sc_hd__mux2_1 _11172_ (.A0(net1191),
    .A1(_05798_),
    .S(_05777_),
    .X(_05799_));
 sky130_fd_sc_hd__clkbuf_1 _11173_ (.A(_05799_),
    .X(_00763_));
 sky130_fd_sc_hd__clkbuf_8 _11174_ (.A(_04110_),
    .X(_05800_));
 sky130_fd_sc_hd__mux2_1 _11175_ (.A0(net530),
    .A1(_05800_),
    .S(_05777_),
    .X(_05801_));
 sky130_fd_sc_hd__clkbuf_1 _11176_ (.A(_05801_),
    .X(_00764_));
 sky130_fd_sc_hd__buf_6 _11177_ (.A(_04113_),
    .X(_05802_));
 sky130_fd_sc_hd__mux2_1 _11178_ (.A0(net899),
    .A1(_05802_),
    .S(_05777_),
    .X(_05803_));
 sky130_fd_sc_hd__clkbuf_1 _11179_ (.A(_05803_),
    .X(_00765_));
 sky130_fd_sc_hd__clkbuf_8 _11180_ (.A(_04116_),
    .X(_05804_));
 sky130_fd_sc_hd__mux2_1 _11181_ (.A0(net1718),
    .A1(_05804_),
    .S(_05777_),
    .X(_05805_));
 sky130_fd_sc_hd__clkbuf_1 _11182_ (.A(_05805_),
    .X(_00766_));
 sky130_fd_sc_hd__buf_6 _11183_ (.A(_04119_),
    .X(_05806_));
 sky130_fd_sc_hd__mux2_1 _11184_ (.A0(net1267),
    .A1(_05806_),
    .S(_05777_),
    .X(_05807_));
 sky130_fd_sc_hd__clkbuf_1 _11185_ (.A(_05807_),
    .X(_00767_));
 sky130_fd_sc_hd__buf_6 _11186_ (.A(_04122_),
    .X(_05808_));
 sky130_fd_sc_hd__mux2_1 _11187_ (.A0(net874),
    .A1(_05808_),
    .S(_05777_),
    .X(_05809_));
 sky130_fd_sc_hd__clkbuf_1 _11188_ (.A(_05809_),
    .X(_00768_));
 sky130_fd_sc_hd__nor2_4 _11189_ (.A(_05757_),
    .B(_04501_),
    .Y(_05810_));
 sky130_fd_sc_hd__buf_4 _11190_ (.A(_05810_),
    .X(_05811_));
 sky130_fd_sc_hd__mux2_1 _11191_ (.A0(net268),
    .A1(_05776_),
    .S(_05811_),
    .X(_05812_));
 sky130_fd_sc_hd__clkbuf_1 _11192_ (.A(_05812_),
    .X(_00769_));
 sky130_fd_sc_hd__mux2_1 _11193_ (.A0(net456),
    .A1(_05780_),
    .S(_05811_),
    .X(_05813_));
 sky130_fd_sc_hd__clkbuf_1 _11194_ (.A(_05813_),
    .X(_00770_));
 sky130_fd_sc_hd__mux2_1 _11195_ (.A0(net66),
    .A1(_05782_),
    .S(_05811_),
    .X(_05814_));
 sky130_fd_sc_hd__clkbuf_1 _11196_ (.A(_05814_),
    .X(_00771_));
 sky130_fd_sc_hd__mux2_1 _11197_ (.A0(net136),
    .A1(_05784_),
    .S(_05811_),
    .X(_05815_));
 sky130_fd_sc_hd__clkbuf_1 _11198_ (.A(_05815_),
    .X(_00772_));
 sky130_fd_sc_hd__mux2_1 _11199_ (.A0(net121),
    .A1(_05786_),
    .S(_05811_),
    .X(_05816_));
 sky130_fd_sc_hd__clkbuf_1 _11200_ (.A(_05816_),
    .X(_00773_));
 sky130_fd_sc_hd__mux2_1 _11201_ (.A0(net439),
    .A1(_05788_),
    .S(_05811_),
    .X(_05817_));
 sky130_fd_sc_hd__clkbuf_1 _11202_ (.A(_05817_),
    .X(_00774_));
 sky130_fd_sc_hd__mux2_1 _11203_ (.A0(net1050),
    .A1(_05790_),
    .S(_05811_),
    .X(_05818_));
 sky130_fd_sc_hd__clkbuf_1 _11204_ (.A(_05818_),
    .X(_00775_));
 sky130_fd_sc_hd__mux2_1 _11205_ (.A0(net317),
    .A1(_05792_),
    .S(_05811_),
    .X(_05819_));
 sky130_fd_sc_hd__clkbuf_1 _11206_ (.A(_05819_),
    .X(_00776_));
 sky130_fd_sc_hd__mux2_1 _11207_ (.A0(net446),
    .A1(_05794_),
    .S(_05811_),
    .X(_05820_));
 sky130_fd_sc_hd__clkbuf_1 _11208_ (.A(_05820_),
    .X(_00777_));
 sky130_fd_sc_hd__mux2_1 _11209_ (.A0(net1460),
    .A1(_05796_),
    .S(_05811_),
    .X(_05821_));
 sky130_fd_sc_hd__clkbuf_1 _11210_ (.A(_05821_),
    .X(_00778_));
 sky130_fd_sc_hd__mux2_1 _11211_ (.A0(net204),
    .A1(_05798_),
    .S(_05810_),
    .X(_05822_));
 sky130_fd_sc_hd__clkbuf_1 _11212_ (.A(_05822_),
    .X(_00779_));
 sky130_fd_sc_hd__mux2_1 _11213_ (.A0(net848),
    .A1(_05800_),
    .S(_05810_),
    .X(_05823_));
 sky130_fd_sc_hd__clkbuf_1 _11214_ (.A(_05823_),
    .X(_00780_));
 sky130_fd_sc_hd__mux2_1 _11215_ (.A0(net488),
    .A1(_05802_),
    .S(_05810_),
    .X(_05824_));
 sky130_fd_sc_hd__clkbuf_1 _11216_ (.A(_05824_),
    .X(_00781_));
 sky130_fd_sc_hd__mux2_1 _11217_ (.A0(net495),
    .A1(_05804_),
    .S(_05810_),
    .X(_05825_));
 sky130_fd_sc_hd__clkbuf_1 _11218_ (.A(_05825_),
    .X(_00782_));
 sky130_fd_sc_hd__mux2_1 _11219_ (.A0(net289),
    .A1(_05806_),
    .S(_05810_),
    .X(_05826_));
 sky130_fd_sc_hd__clkbuf_1 _11220_ (.A(_05826_),
    .X(_00783_));
 sky130_fd_sc_hd__mux2_1 _11221_ (.A0(net217),
    .A1(_05808_),
    .S(_05810_),
    .X(_05827_));
 sky130_fd_sc_hd__clkbuf_1 _11222_ (.A(_05827_),
    .X(_00784_));
 sky130_fd_sc_hd__or2_1 _11223_ (.A(_05757_),
    .B(_04225_),
    .X(_05828_));
 sky130_fd_sc_hd__clkbuf_4 _11224_ (.A(_05828_),
    .X(_05829_));
 sky130_fd_sc_hd__buf_4 _11225_ (.A(_05829_),
    .X(_05830_));
 sky130_fd_sc_hd__mux2_1 _11226_ (.A0(_05648_),
    .A1(net1959),
    .S(_05830_),
    .X(_05831_));
 sky130_fd_sc_hd__clkbuf_1 _11227_ (.A(_05831_),
    .X(_00785_));
 sky130_fd_sc_hd__mux2_1 _11228_ (.A0(_05653_),
    .A1(net2053),
    .S(_05830_),
    .X(_05832_));
 sky130_fd_sc_hd__clkbuf_1 _11229_ (.A(_05832_),
    .X(_00786_));
 sky130_fd_sc_hd__mux2_1 _11230_ (.A0(_05655_),
    .A1(net1943),
    .S(_05830_),
    .X(_05833_));
 sky130_fd_sc_hd__clkbuf_1 _11231_ (.A(_05833_),
    .X(_00787_));
 sky130_fd_sc_hd__mux2_1 _11232_ (.A0(_05657_),
    .A1(net1633),
    .S(_05830_),
    .X(_05834_));
 sky130_fd_sc_hd__clkbuf_1 _11233_ (.A(_05834_),
    .X(_00788_));
 sky130_fd_sc_hd__mux2_1 _11234_ (.A0(_05659_),
    .A1(net1796),
    .S(_05830_),
    .X(_05835_));
 sky130_fd_sc_hd__clkbuf_1 _11235_ (.A(_05835_),
    .X(_00789_));
 sky130_fd_sc_hd__mux2_1 _11236_ (.A0(_05661_),
    .A1(net1981),
    .S(_05830_),
    .X(_05836_));
 sky130_fd_sc_hd__clkbuf_1 _11237_ (.A(_05836_),
    .X(_00790_));
 sky130_fd_sc_hd__mux2_1 _11238_ (.A0(_05663_),
    .A1(net2016),
    .S(_05830_),
    .X(_05837_));
 sky130_fd_sc_hd__clkbuf_1 _11239_ (.A(_05837_),
    .X(_00791_));
 sky130_fd_sc_hd__mux2_1 _11240_ (.A0(_05665_),
    .A1(net1896),
    .S(_05830_),
    .X(_05838_));
 sky130_fd_sc_hd__clkbuf_1 _11241_ (.A(_05838_),
    .X(_00792_));
 sky130_fd_sc_hd__mux2_1 _11242_ (.A0(_05667_),
    .A1(net2010),
    .S(_05830_),
    .X(_05839_));
 sky130_fd_sc_hd__clkbuf_1 _11243_ (.A(_05839_),
    .X(_00793_));
 sky130_fd_sc_hd__mux2_1 _11244_ (.A0(_05669_),
    .A1(net1969),
    .S(_05830_),
    .X(_05840_));
 sky130_fd_sc_hd__clkbuf_1 _11245_ (.A(_05840_),
    .X(_00794_));
 sky130_fd_sc_hd__mux2_1 _11246_ (.A0(_05671_),
    .A1(net1766),
    .S(_05829_),
    .X(_05841_));
 sky130_fd_sc_hd__clkbuf_1 _11247_ (.A(_05841_),
    .X(_00795_));
 sky130_fd_sc_hd__mux2_1 _11248_ (.A0(_05673_),
    .A1(net1817),
    .S(_05829_),
    .X(_05842_));
 sky130_fd_sc_hd__clkbuf_1 _11249_ (.A(_05842_),
    .X(_00796_));
 sky130_fd_sc_hd__mux2_1 _11250_ (.A0(_05675_),
    .A1(net2017),
    .S(_05829_),
    .X(_05843_));
 sky130_fd_sc_hd__clkbuf_1 _11251_ (.A(_05843_),
    .X(_00797_));
 sky130_fd_sc_hd__mux2_1 _11252_ (.A0(_05677_),
    .A1(net1786),
    .S(_05829_),
    .X(_05844_));
 sky130_fd_sc_hd__clkbuf_1 _11253_ (.A(_05844_),
    .X(_00798_));
 sky130_fd_sc_hd__mux2_1 _11254_ (.A0(_05679_),
    .A1(net1872),
    .S(_05829_),
    .X(_05845_));
 sky130_fd_sc_hd__clkbuf_1 _11255_ (.A(_05845_),
    .X(_00799_));
 sky130_fd_sc_hd__mux2_1 _11256_ (.A0(_05681_),
    .A1(net1614),
    .S(_05829_),
    .X(_05846_));
 sky130_fd_sc_hd__clkbuf_1 _11257_ (.A(_05846_),
    .X(_00800_));
 sky130_fd_sc_hd__nor2_4 _11258_ (.A(_05757_),
    .B(_04569_),
    .Y(_05847_));
 sky130_fd_sc_hd__buf_4 _11259_ (.A(_05847_),
    .X(_05848_));
 sky130_fd_sc_hd__mux2_1 _11260_ (.A0(net314),
    .A1(_05776_),
    .S(_05848_),
    .X(_05849_));
 sky130_fd_sc_hd__clkbuf_1 _11261_ (.A(_05849_),
    .X(_00801_));
 sky130_fd_sc_hd__mux2_1 _11262_ (.A0(net122),
    .A1(_05780_),
    .S(_05848_),
    .X(_05850_));
 sky130_fd_sc_hd__clkbuf_1 _11263_ (.A(_05850_),
    .X(_00802_));
 sky130_fd_sc_hd__mux2_1 _11264_ (.A0(net839),
    .A1(_05782_),
    .S(_05848_),
    .X(_05851_));
 sky130_fd_sc_hd__clkbuf_1 _11265_ (.A(_05851_),
    .X(_00803_));
 sky130_fd_sc_hd__mux2_1 _11266_ (.A0(net228),
    .A1(_05784_),
    .S(_05848_),
    .X(_05852_));
 sky130_fd_sc_hd__clkbuf_1 _11267_ (.A(_05852_),
    .X(_00804_));
 sky130_fd_sc_hd__mux2_1 _11268_ (.A0(net116),
    .A1(_05786_),
    .S(_05848_),
    .X(_05853_));
 sky130_fd_sc_hd__clkbuf_1 _11269_ (.A(_05853_),
    .X(_00805_));
 sky130_fd_sc_hd__mux2_1 _11270_ (.A0(net1060),
    .A1(_05788_),
    .S(_05848_),
    .X(_05854_));
 sky130_fd_sc_hd__clkbuf_1 _11271_ (.A(_05854_),
    .X(_00806_));
 sky130_fd_sc_hd__mux2_1 _11272_ (.A0(net46),
    .A1(_05790_),
    .S(_05848_),
    .X(_05855_));
 sky130_fd_sc_hd__clkbuf_1 _11273_ (.A(_05855_),
    .X(_00807_));
 sky130_fd_sc_hd__mux2_1 _11274_ (.A0(net71),
    .A1(_05792_),
    .S(_05848_),
    .X(_05856_));
 sky130_fd_sc_hd__clkbuf_1 _11275_ (.A(_05856_),
    .X(_00808_));
 sky130_fd_sc_hd__mux2_1 _11276_ (.A0(net115),
    .A1(_05794_),
    .S(_05848_),
    .X(_05857_));
 sky130_fd_sc_hd__clkbuf_1 _11277_ (.A(_05857_),
    .X(_00809_));
 sky130_fd_sc_hd__mux2_1 _11278_ (.A0(net216),
    .A1(_05796_),
    .S(_05848_),
    .X(_05858_));
 sky130_fd_sc_hd__clkbuf_1 _11279_ (.A(_05858_),
    .X(_00810_));
 sky130_fd_sc_hd__mux2_1 _11280_ (.A0(net500),
    .A1(_05798_),
    .S(_05847_),
    .X(_05859_));
 sky130_fd_sc_hd__clkbuf_1 _11281_ (.A(_05859_),
    .X(_00811_));
 sky130_fd_sc_hd__mux2_1 _11282_ (.A0(net229),
    .A1(_05800_),
    .S(_05847_),
    .X(_05860_));
 sky130_fd_sc_hd__clkbuf_1 _11283_ (.A(_05860_),
    .X(_00812_));
 sky130_fd_sc_hd__mux2_1 _11284_ (.A0(net359),
    .A1(_05802_),
    .S(_05847_),
    .X(_05861_));
 sky130_fd_sc_hd__clkbuf_1 _11285_ (.A(_05861_),
    .X(_00813_));
 sky130_fd_sc_hd__mux2_1 _11286_ (.A0(net127),
    .A1(_05804_),
    .S(_05847_),
    .X(_05862_));
 sky130_fd_sc_hd__clkbuf_1 _11287_ (.A(_05862_),
    .X(_00814_));
 sky130_fd_sc_hd__mux2_1 _11288_ (.A0(net736),
    .A1(_05806_),
    .S(_05847_),
    .X(_05863_));
 sky130_fd_sc_hd__clkbuf_1 _11289_ (.A(_05863_),
    .X(_00815_));
 sky130_fd_sc_hd__mux2_1 _11290_ (.A0(net165),
    .A1(_05808_),
    .S(_05847_),
    .X(_05864_));
 sky130_fd_sc_hd__clkbuf_1 _11291_ (.A(_05864_),
    .X(_00816_));
 sky130_fd_sc_hd__or2_1 _11292_ (.A(_05757_),
    .B(_04184_),
    .X(_05865_));
 sky130_fd_sc_hd__buf_4 _11293_ (.A(_05865_),
    .X(_05866_));
 sky130_fd_sc_hd__buf_4 _11294_ (.A(_05866_),
    .X(_05867_));
 sky130_fd_sc_hd__mux2_1 _11295_ (.A0(_05648_),
    .A1(net1427),
    .S(_05867_),
    .X(_05868_));
 sky130_fd_sc_hd__clkbuf_1 _11296_ (.A(_05868_),
    .X(_00817_));
 sky130_fd_sc_hd__mux2_1 _11297_ (.A0(_05653_),
    .A1(net1988),
    .S(_05867_),
    .X(_05869_));
 sky130_fd_sc_hd__clkbuf_1 _11298_ (.A(_05869_),
    .X(_00818_));
 sky130_fd_sc_hd__mux2_1 _11299_ (.A0(_05655_),
    .A1(net1768),
    .S(_05867_),
    .X(_05870_));
 sky130_fd_sc_hd__clkbuf_1 _11300_ (.A(_05870_),
    .X(_00819_));
 sky130_fd_sc_hd__mux2_1 _11301_ (.A0(_05657_),
    .A1(net1804),
    .S(_05867_),
    .X(_05871_));
 sky130_fd_sc_hd__clkbuf_1 _11302_ (.A(_05871_),
    .X(_00820_));
 sky130_fd_sc_hd__mux2_1 _11303_ (.A0(_05659_),
    .A1(net1830),
    .S(_05867_),
    .X(_05872_));
 sky130_fd_sc_hd__clkbuf_1 _11304_ (.A(_05872_),
    .X(_00821_));
 sky130_fd_sc_hd__mux2_1 _11305_ (.A0(_05661_),
    .A1(net1974),
    .S(_05867_),
    .X(_05873_));
 sky130_fd_sc_hd__clkbuf_1 _11306_ (.A(_05873_),
    .X(_00822_));
 sky130_fd_sc_hd__mux2_1 _11307_ (.A0(_05663_),
    .A1(net2083),
    .S(_05867_),
    .X(_05874_));
 sky130_fd_sc_hd__clkbuf_1 _11308_ (.A(_05874_),
    .X(_00823_));
 sky130_fd_sc_hd__mux2_1 _11309_ (.A0(_05665_),
    .A1(net1216),
    .S(_05867_),
    .X(_05875_));
 sky130_fd_sc_hd__clkbuf_1 _11310_ (.A(_05875_),
    .X(_00824_));
 sky130_fd_sc_hd__mux2_1 _11311_ (.A0(_05667_),
    .A1(net1108),
    .S(_05867_),
    .X(_05876_));
 sky130_fd_sc_hd__clkbuf_1 _11312_ (.A(_05876_),
    .X(_00825_));
 sky130_fd_sc_hd__mux2_1 _11313_ (.A0(_05669_),
    .A1(net1554),
    .S(_05867_),
    .X(_05877_));
 sky130_fd_sc_hd__clkbuf_1 _11314_ (.A(_05877_),
    .X(_00826_));
 sky130_fd_sc_hd__mux2_1 _11315_ (.A0(_05671_),
    .A1(net1801),
    .S(_05866_),
    .X(_05878_));
 sky130_fd_sc_hd__clkbuf_1 _11316_ (.A(_05878_),
    .X(_00827_));
 sky130_fd_sc_hd__mux2_1 _11317_ (.A0(_05673_),
    .A1(net1544),
    .S(_05866_),
    .X(_05879_));
 sky130_fd_sc_hd__clkbuf_1 _11318_ (.A(_05879_),
    .X(_00828_));
 sky130_fd_sc_hd__mux2_1 _11319_ (.A0(_05675_),
    .A1(net1419),
    .S(_05866_),
    .X(_05880_));
 sky130_fd_sc_hd__clkbuf_1 _11320_ (.A(_05880_),
    .X(_00829_));
 sky130_fd_sc_hd__mux2_1 _11321_ (.A0(_05677_),
    .A1(net1889),
    .S(_05866_),
    .X(_05881_));
 sky130_fd_sc_hd__clkbuf_1 _11322_ (.A(_05881_),
    .X(_00830_));
 sky130_fd_sc_hd__mux2_1 _11323_ (.A0(_05679_),
    .A1(net1555),
    .S(_05866_),
    .X(_05882_));
 sky130_fd_sc_hd__clkbuf_1 _11324_ (.A(_05882_),
    .X(_00831_));
 sky130_fd_sc_hd__mux2_1 _11325_ (.A0(_05681_),
    .A1(net1579),
    .S(_05866_),
    .X(_05883_));
 sky130_fd_sc_hd__clkbuf_1 _11326_ (.A(_05883_),
    .X(_00832_));
 sky130_fd_sc_hd__or2_1 _11327_ (.A(_05757_),
    .B(_04607_),
    .X(_05884_));
 sky130_fd_sc_hd__clkbuf_4 _11328_ (.A(_05884_),
    .X(_05885_));
 sky130_fd_sc_hd__buf_4 _11329_ (.A(_05885_),
    .X(_05886_));
 sky130_fd_sc_hd__mux2_1 _11330_ (.A0(_05648_),
    .A1(net1462),
    .S(_05886_),
    .X(_05887_));
 sky130_fd_sc_hd__clkbuf_1 _11331_ (.A(_05887_),
    .X(_00833_));
 sky130_fd_sc_hd__mux2_1 _11332_ (.A0(_05653_),
    .A1(net2045),
    .S(_05886_),
    .X(_05888_));
 sky130_fd_sc_hd__clkbuf_1 _11333_ (.A(_05888_),
    .X(_00834_));
 sky130_fd_sc_hd__mux2_1 _11334_ (.A0(_05655_),
    .A1(net1929),
    .S(_05886_),
    .X(_05889_));
 sky130_fd_sc_hd__clkbuf_1 _11335_ (.A(_05889_),
    .X(_00835_));
 sky130_fd_sc_hd__mux2_1 _11336_ (.A0(_05657_),
    .A1(net1901),
    .S(_05886_),
    .X(_05890_));
 sky130_fd_sc_hd__clkbuf_1 _11337_ (.A(_05890_),
    .X(_00836_));
 sky130_fd_sc_hd__mux2_1 _11338_ (.A0(_05659_),
    .A1(net1842),
    .S(_05886_),
    .X(_05891_));
 sky130_fd_sc_hd__clkbuf_1 _11339_ (.A(_05891_),
    .X(_00837_));
 sky130_fd_sc_hd__mux2_1 _11340_ (.A0(_05661_),
    .A1(net2061),
    .S(_05886_),
    .X(_05892_));
 sky130_fd_sc_hd__clkbuf_1 _11341_ (.A(_05892_),
    .X(_00838_));
 sky130_fd_sc_hd__mux2_1 _11342_ (.A0(_05663_),
    .A1(net2078),
    .S(_05886_),
    .X(_05893_));
 sky130_fd_sc_hd__clkbuf_1 _11343_ (.A(_05893_),
    .X(_00839_));
 sky130_fd_sc_hd__mux2_1 _11344_ (.A0(_05665_),
    .A1(net1784),
    .S(_05886_),
    .X(_05894_));
 sky130_fd_sc_hd__clkbuf_1 _11345_ (.A(_05894_),
    .X(_00840_));
 sky130_fd_sc_hd__mux2_1 _11346_ (.A0(_05667_),
    .A1(net1992),
    .S(_05886_),
    .X(_05895_));
 sky130_fd_sc_hd__clkbuf_1 _11347_ (.A(_05895_),
    .X(_00841_));
 sky130_fd_sc_hd__mux2_1 _11348_ (.A0(_05669_),
    .A1(net1714),
    .S(_05886_),
    .X(_05896_));
 sky130_fd_sc_hd__clkbuf_1 _11349_ (.A(_05896_),
    .X(_00842_));
 sky130_fd_sc_hd__mux2_1 _11350_ (.A0(_05671_),
    .A1(net1390),
    .S(_05885_),
    .X(_05897_));
 sky130_fd_sc_hd__clkbuf_1 _11351_ (.A(_05897_),
    .X(_00843_));
 sky130_fd_sc_hd__mux2_1 _11352_ (.A0(_05673_),
    .A1(net1604),
    .S(_05885_),
    .X(_05898_));
 sky130_fd_sc_hd__clkbuf_1 _11353_ (.A(_05898_),
    .X(_00844_));
 sky130_fd_sc_hd__mux2_1 _11354_ (.A0(_05675_),
    .A1(net1603),
    .S(_05885_),
    .X(_05899_));
 sky130_fd_sc_hd__clkbuf_1 _11355_ (.A(_05899_),
    .X(_00845_));
 sky130_fd_sc_hd__mux2_1 _11356_ (.A0(_05677_),
    .A1(net1597),
    .S(_05885_),
    .X(_05900_));
 sky130_fd_sc_hd__clkbuf_1 _11357_ (.A(_05900_),
    .X(_00846_));
 sky130_fd_sc_hd__mux2_1 _11358_ (.A0(_05679_),
    .A1(net1963),
    .S(_05885_),
    .X(_05901_));
 sky130_fd_sc_hd__clkbuf_1 _11359_ (.A(_05901_),
    .X(_00847_));
 sky130_fd_sc_hd__mux2_1 _11360_ (.A0(_05681_),
    .A1(net1925),
    .S(_05885_),
    .X(_05902_));
 sky130_fd_sc_hd__clkbuf_1 _11361_ (.A(_05902_),
    .X(_00848_));
 sky130_fd_sc_hd__or3_1 _11362_ (.A(_02498_),
    .B(_05026_),
    .C(_04129_),
    .X(_05903_));
 sky130_fd_sc_hd__clkbuf_4 _11363_ (.A(_05903_),
    .X(_05904_));
 sky130_fd_sc_hd__buf_4 _11364_ (.A(_05904_),
    .X(_05905_));
 sky130_fd_sc_hd__mux2_1 _11365_ (.A0(_05648_),
    .A1(net1785),
    .S(_05905_),
    .X(_05906_));
 sky130_fd_sc_hd__clkbuf_1 _11366_ (.A(_05906_),
    .X(_00849_));
 sky130_fd_sc_hd__mux2_1 _11367_ (.A0(_05653_),
    .A1(net2023),
    .S(_05905_),
    .X(_05907_));
 sky130_fd_sc_hd__clkbuf_1 _11368_ (.A(_05907_),
    .X(_00850_));
 sky130_fd_sc_hd__mux2_1 _11369_ (.A0(_05655_),
    .A1(net1973),
    .S(_05905_),
    .X(_05908_));
 sky130_fd_sc_hd__clkbuf_1 _11370_ (.A(_05908_),
    .X(_00851_));
 sky130_fd_sc_hd__mux2_1 _11371_ (.A0(_05657_),
    .A1(net1863),
    .S(_05905_),
    .X(_05909_));
 sky130_fd_sc_hd__clkbuf_1 _11372_ (.A(_05909_),
    .X(_00852_));
 sky130_fd_sc_hd__mux2_1 _11373_ (.A0(_05659_),
    .A1(net1310),
    .S(_05905_),
    .X(_05910_));
 sky130_fd_sc_hd__clkbuf_1 _11374_ (.A(_05910_),
    .X(_00853_));
 sky130_fd_sc_hd__mux2_1 _11375_ (.A0(_05661_),
    .A1(net2050),
    .S(_05905_),
    .X(_05911_));
 sky130_fd_sc_hd__clkbuf_1 _11376_ (.A(_05911_),
    .X(_00854_));
 sky130_fd_sc_hd__mux2_1 _11377_ (.A0(_05663_),
    .A1(net2071),
    .S(_05905_),
    .X(_05912_));
 sky130_fd_sc_hd__clkbuf_1 _11378_ (.A(_05912_),
    .X(_00855_));
 sky130_fd_sc_hd__mux2_1 _11379_ (.A0(_05665_),
    .A1(net1473),
    .S(_05905_),
    .X(_05913_));
 sky130_fd_sc_hd__clkbuf_1 _11380_ (.A(_05913_),
    .X(_00856_));
 sky130_fd_sc_hd__mux2_1 _11381_ (.A0(_05667_),
    .A1(net2007),
    .S(_05905_),
    .X(_05914_));
 sky130_fd_sc_hd__clkbuf_1 _11382_ (.A(_05914_),
    .X(_00857_));
 sky130_fd_sc_hd__mux2_1 _11383_ (.A0(_05669_),
    .A1(net2008),
    .S(_05905_),
    .X(_05915_));
 sky130_fd_sc_hd__clkbuf_1 _11384_ (.A(_05915_),
    .X(_00858_));
 sky130_fd_sc_hd__mux2_1 _11385_ (.A0(_05671_),
    .A1(net1935),
    .S(_05904_),
    .X(_05916_));
 sky130_fd_sc_hd__clkbuf_1 _11386_ (.A(_05916_),
    .X(_00859_));
 sky130_fd_sc_hd__mux2_1 _11387_ (.A0(_05673_),
    .A1(net1362),
    .S(_05904_),
    .X(_05917_));
 sky130_fd_sc_hd__clkbuf_1 _11388_ (.A(_05917_),
    .X(_00860_));
 sky130_fd_sc_hd__mux2_1 _11389_ (.A0(_05675_),
    .A1(net1477),
    .S(_05904_),
    .X(_05918_));
 sky130_fd_sc_hd__clkbuf_1 _11390_ (.A(_05918_),
    .X(_00861_));
 sky130_fd_sc_hd__mux2_1 _11391_ (.A0(_05677_),
    .A1(net1812),
    .S(_05904_),
    .X(_05919_));
 sky130_fd_sc_hd__clkbuf_1 _11392_ (.A(_05919_),
    .X(_00862_));
 sky130_fd_sc_hd__mux2_1 _11393_ (.A0(_05679_),
    .A1(net1524),
    .S(_05904_),
    .X(_05920_));
 sky130_fd_sc_hd__clkbuf_1 _11394_ (.A(_05920_),
    .X(_00863_));
 sky130_fd_sc_hd__mux2_1 _11395_ (.A0(_05681_),
    .A1(net1895),
    .S(_05904_),
    .X(_05921_));
 sky130_fd_sc_hd__clkbuf_1 _11396_ (.A(_05921_),
    .X(_00864_));
 sky130_fd_sc_hd__nor2_4 _11397_ (.A(_05757_),
    .B(_04646_),
    .Y(_05922_));
 sky130_fd_sc_hd__buf_4 _11398_ (.A(_05922_),
    .X(_05923_));
 sky130_fd_sc_hd__mux2_1 _11399_ (.A0(net1170),
    .A1(_05776_),
    .S(_05923_),
    .X(_05924_));
 sky130_fd_sc_hd__clkbuf_1 _11400_ (.A(_05924_),
    .X(_00865_));
 sky130_fd_sc_hd__mux2_1 _11401_ (.A0(net1976),
    .A1(_05780_),
    .S(_05923_),
    .X(_05925_));
 sky130_fd_sc_hd__clkbuf_1 _11402_ (.A(_05925_),
    .X(_00866_));
 sky130_fd_sc_hd__mux2_1 _11403_ (.A0(net1178),
    .A1(_05782_),
    .S(_05923_),
    .X(_05926_));
 sky130_fd_sc_hd__clkbuf_1 _11404_ (.A(_05926_),
    .X(_00867_));
 sky130_fd_sc_hd__mux2_1 _11405_ (.A0(net1200),
    .A1(_05784_),
    .S(_05923_),
    .X(_05927_));
 sky130_fd_sc_hd__clkbuf_1 _11406_ (.A(_05927_),
    .X(_00868_));
 sky130_fd_sc_hd__mux2_1 _11407_ (.A0(net274),
    .A1(_05786_),
    .S(_05923_),
    .X(_05928_));
 sky130_fd_sc_hd__clkbuf_1 _11408_ (.A(_05928_),
    .X(_00869_));
 sky130_fd_sc_hd__mux2_1 _11409_ (.A0(net2051),
    .A1(_05788_),
    .S(_05923_),
    .X(_05929_));
 sky130_fd_sc_hd__clkbuf_1 _11410_ (.A(_05929_),
    .X(_00870_));
 sky130_fd_sc_hd__mux2_1 _11411_ (.A0(net1105),
    .A1(_05790_),
    .S(_05923_),
    .X(_05930_));
 sky130_fd_sc_hd__clkbuf_1 _11412_ (.A(_05930_),
    .X(_00871_));
 sky130_fd_sc_hd__mux2_1 _11413_ (.A0(net724),
    .A1(_05792_),
    .S(_05923_),
    .X(_05931_));
 sky130_fd_sc_hd__clkbuf_1 _11414_ (.A(_05931_),
    .X(_00872_));
 sky130_fd_sc_hd__mux2_1 _11415_ (.A0(net948),
    .A1(_05794_),
    .S(_05923_),
    .X(_05932_));
 sky130_fd_sc_hd__clkbuf_1 _11416_ (.A(_05932_),
    .X(_00873_));
 sky130_fd_sc_hd__mux2_1 _11417_ (.A0(net1527),
    .A1(_05796_),
    .S(_05923_),
    .X(_05933_));
 sky130_fd_sc_hd__clkbuf_1 _11418_ (.A(_05933_),
    .X(_00874_));
 sky130_fd_sc_hd__mux2_1 _11419_ (.A0(net440),
    .A1(_05798_),
    .S(_05922_),
    .X(_05934_));
 sky130_fd_sc_hd__clkbuf_1 _11420_ (.A(_05934_),
    .X(_00875_));
 sky130_fd_sc_hd__mux2_1 _11421_ (.A0(net921),
    .A1(_05800_),
    .S(_05922_),
    .X(_05935_));
 sky130_fd_sc_hd__clkbuf_1 _11422_ (.A(_05935_),
    .X(_00876_));
 sky130_fd_sc_hd__mux2_1 _11423_ (.A0(net442),
    .A1(_05802_),
    .S(_05922_),
    .X(_05936_));
 sky130_fd_sc_hd__clkbuf_1 _11424_ (.A(_05936_),
    .X(_00877_));
 sky130_fd_sc_hd__mux2_1 _11425_ (.A0(net1274),
    .A1(_05804_),
    .S(_05922_),
    .X(_05937_));
 sky130_fd_sc_hd__clkbuf_1 _11426_ (.A(_05937_),
    .X(_00878_));
 sky130_fd_sc_hd__mux2_1 _11427_ (.A0(net1091),
    .A1(_05806_),
    .S(_05922_),
    .X(_05938_));
 sky130_fd_sc_hd__clkbuf_1 _11428_ (.A(_05938_),
    .X(_00879_));
 sky130_fd_sc_hd__mux2_1 _11429_ (.A0(net1264),
    .A1(_05808_),
    .S(_05922_),
    .X(_05939_));
 sky130_fd_sc_hd__clkbuf_1 _11430_ (.A(_05939_),
    .X(_00880_));
 sky130_fd_sc_hd__nor2_4 _11431_ (.A(_04368_),
    .B(_04646_),
    .Y(_05940_));
 sky130_fd_sc_hd__buf_4 _11432_ (.A(_05940_),
    .X(_05941_));
 sky130_fd_sc_hd__mux2_1 _11433_ (.A0(net1248),
    .A1(_05776_),
    .S(_05941_),
    .X(_05942_));
 sky130_fd_sc_hd__clkbuf_1 _11434_ (.A(_05942_),
    .X(_00881_));
 sky130_fd_sc_hd__mux2_1 _11435_ (.A0(net750),
    .A1(_05780_),
    .S(_05941_),
    .X(_05943_));
 sky130_fd_sc_hd__clkbuf_1 _11436_ (.A(_05943_),
    .X(_00882_));
 sky130_fd_sc_hd__mux2_1 _11437_ (.A0(net160),
    .A1(_05782_),
    .S(_05941_),
    .X(_05944_));
 sky130_fd_sc_hd__clkbuf_1 _11438_ (.A(_05944_),
    .X(_00883_));
 sky130_fd_sc_hd__mux2_1 _11439_ (.A0(net1729),
    .A1(_05784_),
    .S(_05941_),
    .X(_05945_));
 sky130_fd_sc_hd__clkbuf_1 _11440_ (.A(_05945_),
    .X(_00884_));
 sky130_fd_sc_hd__mux2_1 _11441_ (.A0(net102),
    .A1(_05786_),
    .S(_05941_),
    .X(_05946_));
 sky130_fd_sc_hd__clkbuf_1 _11442_ (.A(_05946_),
    .X(_00885_));
 sky130_fd_sc_hd__mux2_1 _11443_ (.A0(net248),
    .A1(_05788_),
    .S(_05941_),
    .X(_05947_));
 sky130_fd_sc_hd__clkbuf_1 _11444_ (.A(_05947_),
    .X(_00886_));
 sky130_fd_sc_hd__mux2_1 _11445_ (.A0(net375),
    .A1(_05790_),
    .S(_05941_),
    .X(_05948_));
 sky130_fd_sc_hd__clkbuf_1 _11446_ (.A(_05948_),
    .X(_00887_));
 sky130_fd_sc_hd__mux2_1 _11447_ (.A0(net93),
    .A1(_05792_),
    .S(_05941_),
    .X(_05949_));
 sky130_fd_sc_hd__clkbuf_1 _11448_ (.A(_05949_),
    .X(_00888_));
 sky130_fd_sc_hd__mux2_1 _11449_ (.A0(net305),
    .A1(_05794_),
    .S(_05941_),
    .X(_05950_));
 sky130_fd_sc_hd__clkbuf_1 _11450_ (.A(_05950_),
    .X(_00889_));
 sky130_fd_sc_hd__mux2_1 _11451_ (.A0(net318),
    .A1(_05796_),
    .S(_05941_),
    .X(_05951_));
 sky130_fd_sc_hd__clkbuf_1 _11452_ (.A(_05951_),
    .X(_00890_));
 sky130_fd_sc_hd__mux2_1 _11453_ (.A0(net1345),
    .A1(_05798_),
    .S(_05940_),
    .X(_05952_));
 sky130_fd_sc_hd__clkbuf_1 _11454_ (.A(_05952_),
    .X(_00891_));
 sky130_fd_sc_hd__mux2_1 _11455_ (.A0(net1501),
    .A1(_05800_),
    .S(_05940_),
    .X(_05953_));
 sky130_fd_sc_hd__clkbuf_1 _11456_ (.A(_05953_),
    .X(_00892_));
 sky130_fd_sc_hd__mux2_1 _11457_ (.A0(net1083),
    .A1(_05802_),
    .S(_05940_),
    .X(_05954_));
 sky130_fd_sc_hd__clkbuf_1 _11458_ (.A(_05954_),
    .X(_00893_));
 sky130_fd_sc_hd__mux2_1 _11459_ (.A0(net1968),
    .A1(_05804_),
    .S(_05940_),
    .X(_05955_));
 sky130_fd_sc_hd__clkbuf_1 _11460_ (.A(_05955_),
    .X(_00894_));
 sky130_fd_sc_hd__mux2_1 _11461_ (.A0(net520),
    .A1(_05806_),
    .S(_05940_),
    .X(_05956_));
 sky130_fd_sc_hd__clkbuf_1 _11462_ (.A(_05956_),
    .X(_00895_));
 sky130_fd_sc_hd__mux2_1 _11463_ (.A0(net2065),
    .A1(_05808_),
    .S(_05940_),
    .X(_05957_));
 sky130_fd_sc_hd__clkbuf_1 _11464_ (.A(_05957_),
    .X(_00896_));
 sky130_fd_sc_hd__or2_1 _11465_ (.A(_05757_),
    .B(_04684_),
    .X(_05958_));
 sky130_fd_sc_hd__clkbuf_4 _11466_ (.A(_05958_),
    .X(_05959_));
 sky130_fd_sc_hd__buf_4 _11467_ (.A(_05959_),
    .X(_05960_));
 sky130_fd_sc_hd__mux2_1 _11468_ (.A0(_05648_),
    .A1(net1504),
    .S(_05960_),
    .X(_05961_));
 sky130_fd_sc_hd__clkbuf_1 _11469_ (.A(_05961_),
    .X(_00897_));
 sky130_fd_sc_hd__mux2_1 _11470_ (.A0(_05653_),
    .A1(net1954),
    .S(_05960_),
    .X(_05962_));
 sky130_fd_sc_hd__clkbuf_1 _11471_ (.A(_05962_),
    .X(_00898_));
 sky130_fd_sc_hd__mux2_1 _11472_ (.A0(_05655_),
    .A1(net1799),
    .S(_05960_),
    .X(_05963_));
 sky130_fd_sc_hd__clkbuf_1 _11473_ (.A(_05963_),
    .X(_00899_));
 sky130_fd_sc_hd__mux2_1 _11474_ (.A0(_05657_),
    .A1(net1506),
    .S(_05960_),
    .X(_05964_));
 sky130_fd_sc_hd__clkbuf_1 _11475_ (.A(_05964_),
    .X(_00900_));
 sky130_fd_sc_hd__mux2_1 _11476_ (.A0(_05659_),
    .A1(net1205),
    .S(_05960_),
    .X(_05965_));
 sky130_fd_sc_hd__clkbuf_1 _11477_ (.A(_05965_),
    .X(_00901_));
 sky130_fd_sc_hd__mux2_1 _11478_ (.A0(_05661_),
    .A1(net1665),
    .S(_05960_),
    .X(_05966_));
 sky130_fd_sc_hd__clkbuf_1 _11479_ (.A(_05966_),
    .X(_00902_));
 sky130_fd_sc_hd__mux2_1 _11480_ (.A0(_05663_),
    .A1(net1982),
    .S(_05960_),
    .X(_05967_));
 sky130_fd_sc_hd__clkbuf_1 _11481_ (.A(_05967_),
    .X(_00903_));
 sky130_fd_sc_hd__mux2_1 _11482_ (.A0(_05665_),
    .A1(net782),
    .S(_05960_),
    .X(_05968_));
 sky130_fd_sc_hd__clkbuf_1 _11483_ (.A(_05968_),
    .X(_00904_));
 sky130_fd_sc_hd__mux2_1 _11484_ (.A0(_05667_),
    .A1(net1636),
    .S(_05960_),
    .X(_05969_));
 sky130_fd_sc_hd__clkbuf_1 _11485_ (.A(_05969_),
    .X(_00905_));
 sky130_fd_sc_hd__mux2_1 _11486_ (.A0(_05669_),
    .A1(net1122),
    .S(_05960_),
    .X(_05970_));
 sky130_fd_sc_hd__clkbuf_1 _11487_ (.A(_05970_),
    .X(_00906_));
 sky130_fd_sc_hd__mux2_1 _11488_ (.A0(_05671_),
    .A1(net1285),
    .S(_05959_),
    .X(_05971_));
 sky130_fd_sc_hd__clkbuf_1 _11489_ (.A(_05971_),
    .X(_00907_));
 sky130_fd_sc_hd__mux2_1 _11490_ (.A0(_05673_),
    .A1(net1475),
    .S(_05959_),
    .X(_05972_));
 sky130_fd_sc_hd__clkbuf_1 _11491_ (.A(_05972_),
    .X(_00908_));
 sky130_fd_sc_hd__mux2_1 _11492_ (.A0(_05675_),
    .A1(net1157),
    .S(_05959_),
    .X(_05973_));
 sky130_fd_sc_hd__clkbuf_1 _11493_ (.A(_05973_),
    .X(_00909_));
 sky130_fd_sc_hd__mux2_1 _11494_ (.A0(_05677_),
    .A1(net1704),
    .S(_05959_),
    .X(_05974_));
 sky130_fd_sc_hd__clkbuf_1 _11495_ (.A(_05974_),
    .X(_00910_));
 sky130_fd_sc_hd__mux2_1 _11496_ (.A0(_05679_),
    .A1(net1862),
    .S(_05959_),
    .X(_05975_));
 sky130_fd_sc_hd__clkbuf_1 _11497_ (.A(_05975_),
    .X(_00911_));
 sky130_fd_sc_hd__mux2_1 _11498_ (.A0(_05681_),
    .A1(net1760),
    .S(_05959_),
    .X(_05976_));
 sky130_fd_sc_hd__clkbuf_1 _11499_ (.A(_05976_),
    .X(_00912_));
 sky130_fd_sc_hd__or3_1 _11500_ (.A(_02506_),
    .B(_05026_),
    .C(_04129_),
    .X(_05977_));
 sky130_fd_sc_hd__clkbuf_4 _11501_ (.A(_05977_),
    .X(_05978_));
 sky130_fd_sc_hd__buf_4 _11502_ (.A(_05978_),
    .X(_05979_));
 sky130_fd_sc_hd__mux2_1 _11503_ (.A0(_05648_),
    .A1(net1745),
    .S(_05979_),
    .X(_05980_));
 sky130_fd_sc_hd__clkbuf_1 _11504_ (.A(_05980_),
    .X(_00913_));
 sky130_fd_sc_hd__mux2_1 _11505_ (.A0(_05653_),
    .A1(net1996),
    .S(_05979_),
    .X(_05981_));
 sky130_fd_sc_hd__clkbuf_1 _11506_ (.A(_05981_),
    .X(_00914_));
 sky130_fd_sc_hd__mux2_1 _11507_ (.A0(_05655_),
    .A1(net1835),
    .S(_05979_),
    .X(_05982_));
 sky130_fd_sc_hd__clkbuf_1 _11508_ (.A(_05982_),
    .X(_00915_));
 sky130_fd_sc_hd__mux2_1 _11509_ (.A0(_05657_),
    .A1(net1410),
    .S(_05979_),
    .X(_05983_));
 sky130_fd_sc_hd__clkbuf_1 _11510_ (.A(_05983_),
    .X(_00916_));
 sky130_fd_sc_hd__mux2_1 _11511_ (.A0(_05659_),
    .A1(net1562),
    .S(_05979_),
    .X(_05984_));
 sky130_fd_sc_hd__clkbuf_1 _11512_ (.A(_05984_),
    .X(_00917_));
 sky130_fd_sc_hd__mux2_1 _11513_ (.A0(_05661_),
    .A1(net1939),
    .S(_05979_),
    .X(_05985_));
 sky130_fd_sc_hd__clkbuf_1 _11514_ (.A(_05985_),
    .X(_00918_));
 sky130_fd_sc_hd__mux2_1 _11515_ (.A0(_05663_),
    .A1(net2052),
    .S(_05979_),
    .X(_05986_));
 sky130_fd_sc_hd__clkbuf_1 _11516_ (.A(_05986_),
    .X(_00919_));
 sky130_fd_sc_hd__mux2_1 _11517_ (.A0(_05665_),
    .A1(net1721),
    .S(_05979_),
    .X(_05987_));
 sky130_fd_sc_hd__clkbuf_1 _11518_ (.A(_05987_),
    .X(_00920_));
 sky130_fd_sc_hd__mux2_1 _11519_ (.A0(_05667_),
    .A1(net1980),
    .S(_05979_),
    .X(_05988_));
 sky130_fd_sc_hd__clkbuf_1 _11520_ (.A(_05988_),
    .X(_00921_));
 sky130_fd_sc_hd__mux2_1 _11521_ (.A0(_05669_),
    .A1(net1915),
    .S(_05979_),
    .X(_05989_));
 sky130_fd_sc_hd__clkbuf_1 _11522_ (.A(_05989_),
    .X(_00922_));
 sky130_fd_sc_hd__mux2_1 _11523_ (.A0(_05671_),
    .A1(net1956),
    .S(_05978_),
    .X(_05990_));
 sky130_fd_sc_hd__clkbuf_1 _11524_ (.A(_05990_),
    .X(_00923_));
 sky130_fd_sc_hd__mux2_1 _11525_ (.A0(_05673_),
    .A1(net1695),
    .S(_05978_),
    .X(_05991_));
 sky130_fd_sc_hd__clkbuf_1 _11526_ (.A(_05991_),
    .X(_00924_));
 sky130_fd_sc_hd__mux2_1 _11527_ (.A0(_05675_),
    .A1(net1966),
    .S(_05978_),
    .X(_05992_));
 sky130_fd_sc_hd__clkbuf_1 _11528_ (.A(_05992_),
    .X(_00925_));
 sky130_fd_sc_hd__mux2_1 _11529_ (.A0(_05677_),
    .A1(net1546),
    .S(_05978_),
    .X(_05993_));
 sky130_fd_sc_hd__clkbuf_1 _11530_ (.A(_05993_),
    .X(_00926_));
 sky130_fd_sc_hd__mux2_1 _11531_ (.A0(_05679_),
    .A1(net1882),
    .S(_05978_),
    .X(_05994_));
 sky130_fd_sc_hd__clkbuf_1 _11532_ (.A(_05994_),
    .X(_00927_));
 sky130_fd_sc_hd__mux2_1 _11533_ (.A0(_05681_),
    .A1(net1316),
    .S(_05978_),
    .X(_05995_));
 sky130_fd_sc_hd__clkbuf_1 _11534_ (.A(_05995_),
    .X(_00928_));
 sky130_fd_sc_hd__buf_6 _11535_ (.A(_04069_),
    .X(_05996_));
 sky130_fd_sc_hd__or2_1 _11536_ (.A(_04129_),
    .B(_04365_),
    .X(_05997_));
 sky130_fd_sc_hd__clkbuf_4 _11537_ (.A(_05997_),
    .X(_05998_));
 sky130_fd_sc_hd__buf_4 _11538_ (.A(_05998_),
    .X(_05999_));
 sky130_fd_sc_hd__mux2_1 _11539_ (.A0(_05996_),
    .A1(net1550),
    .S(_05999_),
    .X(_06000_));
 sky130_fd_sc_hd__clkbuf_1 _11540_ (.A(_06000_),
    .X(_00929_));
 sky130_fd_sc_hd__buf_4 _11541_ (.A(_04080_),
    .X(_06001_));
 sky130_fd_sc_hd__mux2_1 _11542_ (.A0(_06001_),
    .A1(net632),
    .S(_05999_),
    .X(_06002_));
 sky130_fd_sc_hd__clkbuf_1 _11543_ (.A(_06002_),
    .X(_00930_));
 sky130_fd_sc_hd__buf_6 _11544_ (.A(_04083_),
    .X(_06003_));
 sky130_fd_sc_hd__mux2_1 _11545_ (.A0(_06003_),
    .A1(net346),
    .S(_05999_),
    .X(_06004_));
 sky130_fd_sc_hd__clkbuf_1 _11546_ (.A(_06004_),
    .X(_00931_));
 sky130_fd_sc_hd__buf_6 _11547_ (.A(_04086_),
    .X(_06005_));
 sky130_fd_sc_hd__mux2_1 _11548_ (.A0(_06005_),
    .A1(net425),
    .S(_05999_),
    .X(_06006_));
 sky130_fd_sc_hd__clkbuf_1 _11549_ (.A(_06006_),
    .X(_00932_));
 sky130_fd_sc_hd__buf_6 _11550_ (.A(_04089_),
    .X(_06007_));
 sky130_fd_sc_hd__mux2_1 _11551_ (.A0(_06007_),
    .A1(net608),
    .S(_05999_),
    .X(_06008_));
 sky130_fd_sc_hd__clkbuf_1 _11552_ (.A(_06008_),
    .X(_00933_));
 sky130_fd_sc_hd__buf_4 _11553_ (.A(_04092_),
    .X(_06009_));
 sky130_fd_sc_hd__mux2_1 _11554_ (.A0(_06009_),
    .A1(net737),
    .S(_05999_),
    .X(_06010_));
 sky130_fd_sc_hd__clkbuf_1 _11555_ (.A(_06010_),
    .X(_00934_));
 sky130_fd_sc_hd__buf_4 _11556_ (.A(_04095_),
    .X(_06011_));
 sky130_fd_sc_hd__mux2_1 _11557_ (.A0(_06011_),
    .A1(net703),
    .S(_05999_),
    .X(_06012_));
 sky130_fd_sc_hd__clkbuf_1 _11558_ (.A(_06012_),
    .X(_00935_));
 sky130_fd_sc_hd__buf_6 _11559_ (.A(_04098_),
    .X(_06013_));
 sky130_fd_sc_hd__mux2_1 _11560_ (.A0(_06013_),
    .A1(net1103),
    .S(_05999_),
    .X(_06014_));
 sky130_fd_sc_hd__clkbuf_1 _11561_ (.A(_06014_),
    .X(_00936_));
 sky130_fd_sc_hd__buf_6 _11562_ (.A(_04101_),
    .X(_06015_));
 sky130_fd_sc_hd__mux2_1 _11563_ (.A0(_06015_),
    .A1(net1231),
    .S(_05999_),
    .X(_06016_));
 sky130_fd_sc_hd__clkbuf_1 _11564_ (.A(_06016_),
    .X(_00937_));
 sky130_fd_sc_hd__buf_6 _11565_ (.A(_04104_),
    .X(_06017_));
 sky130_fd_sc_hd__mux2_1 _11566_ (.A0(_06017_),
    .A1(net915),
    .S(_05999_),
    .X(_06018_));
 sky130_fd_sc_hd__clkbuf_1 _11567_ (.A(_06018_),
    .X(_00938_));
 sky130_fd_sc_hd__buf_6 _11568_ (.A(_04107_),
    .X(_06019_));
 sky130_fd_sc_hd__mux2_1 _11569_ (.A0(_06019_),
    .A1(net501),
    .S(_05998_),
    .X(_06020_));
 sky130_fd_sc_hd__clkbuf_1 _11570_ (.A(_06020_),
    .X(_00939_));
 sky130_fd_sc_hd__buf_4 _11571_ (.A(_04110_),
    .X(_06021_));
 sky130_fd_sc_hd__mux2_1 _11572_ (.A0(_06021_),
    .A1(net1654),
    .S(_05998_),
    .X(_06022_));
 sky130_fd_sc_hd__clkbuf_1 _11573_ (.A(_06022_),
    .X(_00940_));
 sky130_fd_sc_hd__buf_6 _11574_ (.A(_04113_),
    .X(_06023_));
 sky130_fd_sc_hd__mux2_1 _11575_ (.A0(_06023_),
    .A1(net963),
    .S(_05998_),
    .X(_06024_));
 sky130_fd_sc_hd__clkbuf_1 _11576_ (.A(_06024_),
    .X(_00941_));
 sky130_fd_sc_hd__buf_4 _11577_ (.A(_04116_),
    .X(_06025_));
 sky130_fd_sc_hd__mux2_1 _11578_ (.A0(_06025_),
    .A1(net291),
    .S(_05998_),
    .X(_06026_));
 sky130_fd_sc_hd__clkbuf_1 _11579_ (.A(_06026_),
    .X(_00942_));
 sky130_fd_sc_hd__clkbuf_8 _11580_ (.A(_04119_),
    .X(_06027_));
 sky130_fd_sc_hd__mux2_1 _11581_ (.A0(_06027_),
    .A1(net733),
    .S(_05998_),
    .X(_06028_));
 sky130_fd_sc_hd__clkbuf_1 _11582_ (.A(_06028_),
    .X(_00943_));
 sky130_fd_sc_hd__buf_6 _11583_ (.A(_04122_),
    .X(_06029_));
 sky130_fd_sc_hd__mux2_1 _11584_ (.A0(_06029_),
    .A1(net664),
    .S(_05998_),
    .X(_06030_));
 sky130_fd_sc_hd__clkbuf_1 _11585_ (.A(_06030_),
    .X(_00944_));
 sky130_fd_sc_hd__or3_1 _11586_ (.A(_02484_),
    .B(_02737_),
    .C(_04129_),
    .X(_06031_));
 sky130_fd_sc_hd__clkbuf_4 _11587_ (.A(_06031_),
    .X(_06032_));
 sky130_fd_sc_hd__buf_4 _11588_ (.A(_06032_),
    .X(_06033_));
 sky130_fd_sc_hd__mux2_1 _11589_ (.A0(_05996_),
    .A1(net1885),
    .S(_06033_),
    .X(_06034_));
 sky130_fd_sc_hd__clkbuf_1 _11590_ (.A(_06034_),
    .X(_00945_));
 sky130_fd_sc_hd__mux2_1 _11591_ (.A0(_06001_),
    .A1(net2006),
    .S(_06033_),
    .X(_06035_));
 sky130_fd_sc_hd__clkbuf_1 _11592_ (.A(_06035_),
    .X(_00946_));
 sky130_fd_sc_hd__mux2_1 _11593_ (.A0(_06003_),
    .A1(net1378),
    .S(_06033_),
    .X(_06036_));
 sky130_fd_sc_hd__clkbuf_1 _11594_ (.A(_06036_),
    .X(_00947_));
 sky130_fd_sc_hd__mux2_1 _11595_ (.A0(_06005_),
    .A1(net1556),
    .S(_06033_),
    .X(_06037_));
 sky130_fd_sc_hd__clkbuf_1 _11596_ (.A(_06037_),
    .X(_00948_));
 sky130_fd_sc_hd__mux2_1 _11597_ (.A0(_06007_),
    .A1(net1720),
    .S(_06033_),
    .X(_06038_));
 sky130_fd_sc_hd__clkbuf_1 _11598_ (.A(_06038_),
    .X(_00949_));
 sky130_fd_sc_hd__mux2_1 _11599_ (.A0(_06009_),
    .A1(net1502),
    .S(_06033_),
    .X(_06039_));
 sky130_fd_sc_hd__clkbuf_1 _11600_ (.A(_06039_),
    .X(_00950_));
 sky130_fd_sc_hd__mux2_1 _11601_ (.A0(_06011_),
    .A1(net1238),
    .S(_06033_),
    .X(_06040_));
 sky130_fd_sc_hd__clkbuf_1 _11602_ (.A(_06040_),
    .X(_00951_));
 sky130_fd_sc_hd__mux2_1 _11603_ (.A0(_06013_),
    .A1(net1241),
    .S(_06033_),
    .X(_06041_));
 sky130_fd_sc_hd__clkbuf_1 _11604_ (.A(_06041_),
    .X(_00952_));
 sky130_fd_sc_hd__mux2_1 _11605_ (.A0(_06015_),
    .A1(net1533),
    .S(_06033_),
    .X(_06042_));
 sky130_fd_sc_hd__clkbuf_1 _11606_ (.A(_06042_),
    .X(_00953_));
 sky130_fd_sc_hd__mux2_1 _11607_ (.A0(_06017_),
    .A1(net1690),
    .S(_06033_),
    .X(_06043_));
 sky130_fd_sc_hd__clkbuf_1 _11608_ (.A(_06043_),
    .X(_00954_));
 sky130_fd_sc_hd__mux2_1 _11609_ (.A0(_06019_),
    .A1(net2037),
    .S(_06032_),
    .X(_06044_));
 sky130_fd_sc_hd__clkbuf_1 _11610_ (.A(_06044_),
    .X(_00955_));
 sky130_fd_sc_hd__mux2_1 _11611_ (.A0(_06021_),
    .A1(net1857),
    .S(_06032_),
    .X(_06045_));
 sky130_fd_sc_hd__clkbuf_1 _11612_ (.A(_06045_),
    .X(_00956_));
 sky130_fd_sc_hd__mux2_1 _11613_ (.A0(_06023_),
    .A1(net1909),
    .S(_06032_),
    .X(_06046_));
 sky130_fd_sc_hd__clkbuf_1 _11614_ (.A(_06046_),
    .X(_00957_));
 sky130_fd_sc_hd__mux2_1 _11615_ (.A0(_06025_),
    .A1(net1375),
    .S(_06032_),
    .X(_06047_));
 sky130_fd_sc_hd__clkbuf_1 _11616_ (.A(_06047_),
    .X(_00958_));
 sky130_fd_sc_hd__mux2_1 _11617_ (.A0(_06027_),
    .A1(net1787),
    .S(_06032_),
    .X(_06048_));
 sky130_fd_sc_hd__clkbuf_1 _11618_ (.A(_06048_),
    .X(_00959_));
 sky130_fd_sc_hd__mux2_1 _11619_ (.A0(_06029_),
    .A1(net1474),
    .S(_06032_),
    .X(_06049_));
 sky130_fd_sc_hd__clkbuf_1 _11620_ (.A(_06049_),
    .X(_00960_));
 sky130_fd_sc_hd__nand2b_4 _11621_ (.A_N(_05757_),
    .B(_04408_),
    .Y(_06050_));
 sky130_fd_sc_hd__buf_4 _11622_ (.A(_06050_),
    .X(_06051_));
 sky130_fd_sc_hd__mux2_1 _11623_ (.A0(_05996_),
    .A1(net1986),
    .S(_06051_),
    .X(_06052_));
 sky130_fd_sc_hd__clkbuf_1 _11624_ (.A(_06052_),
    .X(_00961_));
 sky130_fd_sc_hd__mux2_1 _11625_ (.A0(_06001_),
    .A1(net1679),
    .S(_06051_),
    .X(_06053_));
 sky130_fd_sc_hd__clkbuf_1 _11626_ (.A(_06053_),
    .X(_00962_));
 sky130_fd_sc_hd__mux2_1 _11627_ (.A0(_06003_),
    .A1(net1881),
    .S(_06051_),
    .X(_06054_));
 sky130_fd_sc_hd__clkbuf_1 _11628_ (.A(_06054_),
    .X(_00963_));
 sky130_fd_sc_hd__mux2_1 _11629_ (.A0(_06005_),
    .A1(net1674),
    .S(_06051_),
    .X(_06055_));
 sky130_fd_sc_hd__clkbuf_1 _11630_ (.A(_06055_),
    .X(_00964_));
 sky130_fd_sc_hd__mux2_1 _11631_ (.A0(_06007_),
    .A1(net1752),
    .S(_06051_),
    .X(_06056_));
 sky130_fd_sc_hd__clkbuf_1 _11632_ (.A(_06056_),
    .X(_00965_));
 sky130_fd_sc_hd__mux2_1 _11633_ (.A0(_06009_),
    .A1(net1167),
    .S(_06051_),
    .X(_06057_));
 sky130_fd_sc_hd__clkbuf_1 _11634_ (.A(_06057_),
    .X(_00966_));
 sky130_fd_sc_hd__mux2_1 _11635_ (.A0(_06011_),
    .A1(net1648),
    .S(_06051_),
    .X(_06058_));
 sky130_fd_sc_hd__clkbuf_1 _11636_ (.A(_06058_),
    .X(_00967_));
 sky130_fd_sc_hd__mux2_1 _11637_ (.A0(_06013_),
    .A1(net1659),
    .S(_06051_),
    .X(_06059_));
 sky130_fd_sc_hd__clkbuf_1 _11638_ (.A(_06059_),
    .X(_00968_));
 sky130_fd_sc_hd__mux2_1 _11639_ (.A0(_06015_),
    .A1(net1814),
    .S(_06051_),
    .X(_06060_));
 sky130_fd_sc_hd__clkbuf_1 _11640_ (.A(_06060_),
    .X(_00969_));
 sky130_fd_sc_hd__mux2_1 _11641_ (.A0(_06017_),
    .A1(net1950),
    .S(_06051_),
    .X(_06061_));
 sky130_fd_sc_hd__clkbuf_1 _11642_ (.A(_06061_),
    .X(_00970_));
 sky130_fd_sc_hd__mux2_1 _11643_ (.A0(_06019_),
    .A1(net1767),
    .S(_06050_),
    .X(_06062_));
 sky130_fd_sc_hd__clkbuf_1 _11644_ (.A(_06062_),
    .X(_00971_));
 sky130_fd_sc_hd__mux2_1 _11645_ (.A0(_06021_),
    .A1(net1849),
    .S(_06050_),
    .X(_06063_));
 sky130_fd_sc_hd__clkbuf_1 _11646_ (.A(_06063_),
    .X(_00972_));
 sky130_fd_sc_hd__mux2_1 _11647_ (.A0(_06023_),
    .A1(net1911),
    .S(_06050_),
    .X(_06064_));
 sky130_fd_sc_hd__clkbuf_1 _11648_ (.A(_06064_),
    .X(_00973_));
 sky130_fd_sc_hd__mux2_1 _11649_ (.A0(_06025_),
    .A1(net1877),
    .S(_06050_),
    .X(_06065_));
 sky130_fd_sc_hd__clkbuf_1 _11650_ (.A(_06065_),
    .X(_00974_));
 sky130_fd_sc_hd__mux2_1 _11651_ (.A0(_06027_),
    .A1(net831),
    .S(_06050_),
    .X(_06066_));
 sky130_fd_sc_hd__clkbuf_1 _11652_ (.A(_06066_),
    .X(_00975_));
 sky130_fd_sc_hd__mux2_1 _11653_ (.A0(_06029_),
    .A1(net1892),
    .S(_06050_),
    .X(_06067_));
 sky130_fd_sc_hd__clkbuf_1 _11654_ (.A(_06067_),
    .X(_00976_));
 sky130_fd_sc_hd__or3_1 _11655_ (.A(_02484_),
    .B(_05026_),
    .C(_04129_),
    .X(_06068_));
 sky130_fd_sc_hd__clkbuf_4 _11656_ (.A(_06068_),
    .X(_06069_));
 sky130_fd_sc_hd__buf_4 _11657_ (.A(_06069_),
    .X(_06070_));
 sky130_fd_sc_hd__mux2_1 _11658_ (.A0(_05996_),
    .A1(net1343),
    .S(_06070_),
    .X(_06071_));
 sky130_fd_sc_hd__clkbuf_1 _11659_ (.A(_06071_),
    .X(_00977_));
 sky130_fd_sc_hd__mux2_1 _11660_ (.A0(_06001_),
    .A1(net1997),
    .S(_06070_),
    .X(_06072_));
 sky130_fd_sc_hd__clkbuf_1 _11661_ (.A(_06072_),
    .X(_00978_));
 sky130_fd_sc_hd__mux2_1 _11662_ (.A0(_06003_),
    .A1(net1734),
    .S(_06070_),
    .X(_06073_));
 sky130_fd_sc_hd__clkbuf_1 _11663_ (.A(_06073_),
    .X(_00979_));
 sky130_fd_sc_hd__mux2_1 _11664_ (.A0(_06005_),
    .A1(net1781),
    .S(_06070_),
    .X(_06074_));
 sky130_fd_sc_hd__clkbuf_1 _11665_ (.A(_06074_),
    .X(_00980_));
 sky130_fd_sc_hd__mux2_1 _11666_ (.A0(_06007_),
    .A1(net1609),
    .S(_06070_),
    .X(_06075_));
 sky130_fd_sc_hd__clkbuf_1 _11667_ (.A(_06075_),
    .X(_00981_));
 sky130_fd_sc_hd__mux2_1 _11668_ (.A0(_06009_),
    .A1(net1845),
    .S(_06070_),
    .X(_06076_));
 sky130_fd_sc_hd__clkbuf_1 _11669_ (.A(_06076_),
    .X(_00982_));
 sky130_fd_sc_hd__mux2_1 _11670_ (.A0(_06011_),
    .A1(net1800),
    .S(_06070_),
    .X(_06077_));
 sky130_fd_sc_hd__clkbuf_1 _11671_ (.A(_06077_),
    .X(_00983_));
 sky130_fd_sc_hd__mux2_1 _11672_ (.A0(_06013_),
    .A1(net1479),
    .S(_06070_),
    .X(_06078_));
 sky130_fd_sc_hd__clkbuf_1 _11673_ (.A(_06078_),
    .X(_00984_));
 sky130_fd_sc_hd__mux2_1 _11674_ (.A0(_06015_),
    .A1(net1683),
    .S(_06070_),
    .X(_06079_));
 sky130_fd_sc_hd__clkbuf_1 _11675_ (.A(_06079_),
    .X(_00985_));
 sky130_fd_sc_hd__mux2_1 _11676_ (.A0(_06017_),
    .A1(net1696),
    .S(_06070_),
    .X(_06080_));
 sky130_fd_sc_hd__clkbuf_1 _11677_ (.A(_06080_),
    .X(_00986_));
 sky130_fd_sc_hd__mux2_1 _11678_ (.A0(_06019_),
    .A1(net1854),
    .S(_06069_),
    .X(_06081_));
 sky130_fd_sc_hd__clkbuf_1 _11679_ (.A(_06081_),
    .X(_00987_));
 sky130_fd_sc_hd__mux2_1 _11680_ (.A0(_06021_),
    .A1(net1433),
    .S(_06069_),
    .X(_06082_));
 sky130_fd_sc_hd__clkbuf_1 _11681_ (.A(_06082_),
    .X(_00988_));
 sky130_fd_sc_hd__mux2_1 _11682_ (.A0(_06023_),
    .A1(net1713),
    .S(_06069_),
    .X(_06083_));
 sky130_fd_sc_hd__clkbuf_1 _11683_ (.A(_06083_),
    .X(_00989_));
 sky130_fd_sc_hd__mux2_1 _11684_ (.A0(_06025_),
    .A1(net1174),
    .S(_06069_),
    .X(_06084_));
 sky130_fd_sc_hd__clkbuf_1 _11685_ (.A(_06084_),
    .X(_00990_));
 sky130_fd_sc_hd__mux2_1 _11686_ (.A0(_06027_),
    .A1(net1441),
    .S(_06069_),
    .X(_06085_));
 sky130_fd_sc_hd__clkbuf_1 _11687_ (.A(_06085_),
    .X(_00991_));
 sky130_fd_sc_hd__mux2_1 _11688_ (.A0(_06029_),
    .A1(net2014),
    .S(_06069_),
    .X(_06086_));
 sky130_fd_sc_hd__clkbuf_1 _11689_ (.A(_06086_),
    .X(_00992_));
 sky130_fd_sc_hd__nor2_4 _11690_ (.A(_04286_),
    .B(_04461_),
    .Y(_06087_));
 sky130_fd_sc_hd__buf_4 _11691_ (.A(_06087_),
    .X(_06088_));
 sky130_fd_sc_hd__mux2_1 _11692_ (.A0(net621),
    .A1(_05776_),
    .S(_06088_),
    .X(_06089_));
 sky130_fd_sc_hd__clkbuf_1 _11693_ (.A(_06089_),
    .X(_00993_));
 sky130_fd_sc_hd__mux2_1 _11694_ (.A0(net672),
    .A1(_05780_),
    .S(_06088_),
    .X(_06090_));
 sky130_fd_sc_hd__clkbuf_1 _11695_ (.A(_06090_),
    .X(_00994_));
 sky130_fd_sc_hd__mux2_1 _11696_ (.A0(net582),
    .A1(_05782_),
    .S(_06088_),
    .X(_06091_));
 sky130_fd_sc_hd__clkbuf_1 _11697_ (.A(_06091_),
    .X(_00995_));
 sky130_fd_sc_hd__mux2_1 _11698_ (.A0(net259),
    .A1(_05784_),
    .S(_06088_),
    .X(_06092_));
 sky130_fd_sc_hd__clkbuf_1 _11699_ (.A(_06092_),
    .X(_00996_));
 sky130_fd_sc_hd__mux2_1 _11700_ (.A0(net405),
    .A1(_05786_),
    .S(_06088_),
    .X(_06093_));
 sky130_fd_sc_hd__clkbuf_1 _11701_ (.A(_06093_),
    .X(_00997_));
 sky130_fd_sc_hd__mux2_1 _11702_ (.A0(net1014),
    .A1(_05788_),
    .S(_06088_),
    .X(_06094_));
 sky130_fd_sc_hd__clkbuf_1 _11703_ (.A(_06094_),
    .X(_00998_));
 sky130_fd_sc_hd__mux2_1 _11704_ (.A0(net543),
    .A1(_05790_),
    .S(_06088_),
    .X(_06095_));
 sky130_fd_sc_hd__clkbuf_1 _11705_ (.A(_06095_),
    .X(_00999_));
 sky130_fd_sc_hd__mux2_1 _11706_ (.A0(net628),
    .A1(_05792_),
    .S(_06088_),
    .X(_06096_));
 sky130_fd_sc_hd__clkbuf_1 _11707_ (.A(_06096_),
    .X(_01000_));
 sky130_fd_sc_hd__mux2_1 _11708_ (.A0(net429),
    .A1(_05794_),
    .S(_06088_),
    .X(_06097_));
 sky130_fd_sc_hd__clkbuf_1 _11709_ (.A(_06097_),
    .X(_01001_));
 sky130_fd_sc_hd__mux2_1 _11710_ (.A0(net83),
    .A1(_05796_),
    .S(_06088_),
    .X(_06098_));
 sky130_fd_sc_hd__clkbuf_1 _11711_ (.A(_06098_),
    .X(_01002_));
 sky130_fd_sc_hd__mux2_1 _11712_ (.A0(net512),
    .A1(_05798_),
    .S(_06087_),
    .X(_06099_));
 sky130_fd_sc_hd__clkbuf_1 _11713_ (.A(_06099_),
    .X(_01003_));
 sky130_fd_sc_hd__mux2_1 _11714_ (.A0(net153),
    .A1(_05800_),
    .S(_06087_),
    .X(_06100_));
 sky130_fd_sc_hd__clkbuf_1 _11715_ (.A(_06100_),
    .X(_01004_));
 sky130_fd_sc_hd__mux2_1 _11716_ (.A0(net928),
    .A1(_05802_),
    .S(_06087_),
    .X(_06101_));
 sky130_fd_sc_hd__clkbuf_1 _11717_ (.A(_06101_),
    .X(_01005_));
 sky130_fd_sc_hd__mux2_1 _11718_ (.A0(net541),
    .A1(_05804_),
    .S(_06087_),
    .X(_06102_));
 sky130_fd_sc_hd__clkbuf_1 _11719_ (.A(_06102_),
    .X(_01006_));
 sky130_fd_sc_hd__mux2_1 _11720_ (.A0(net773),
    .A1(_05806_),
    .S(_06087_),
    .X(_06103_));
 sky130_fd_sc_hd__clkbuf_1 _11721_ (.A(_06103_),
    .X(_01007_));
 sky130_fd_sc_hd__mux2_1 _11722_ (.A0(net597),
    .A1(_05808_),
    .S(_06087_),
    .X(_06104_));
 sky130_fd_sc_hd__clkbuf_1 _11723_ (.A(_06104_),
    .X(_01008_));
 sky130_fd_sc_hd__nor2_4 _11724_ (.A(_04072_),
    .B(_04286_),
    .Y(_06105_));
 sky130_fd_sc_hd__buf_6 _11725_ (.A(_06105_),
    .X(_06106_));
 sky130_fd_sc_hd__mux2_1 _11726_ (.A0(net358),
    .A1(_05776_),
    .S(_06106_),
    .X(_06107_));
 sky130_fd_sc_hd__clkbuf_1 _11727_ (.A(_06107_),
    .X(_01009_));
 sky130_fd_sc_hd__mux2_1 _11728_ (.A0(net155),
    .A1(_05780_),
    .S(_06106_),
    .X(_06108_));
 sky130_fd_sc_hd__clkbuf_1 _11729_ (.A(_06108_),
    .X(_01010_));
 sky130_fd_sc_hd__mux2_1 _11730_ (.A0(net1092),
    .A1(_05782_),
    .S(_06106_),
    .X(_06109_));
 sky130_fd_sc_hd__clkbuf_1 _11731_ (.A(_06109_),
    .X(_01011_));
 sky130_fd_sc_hd__mux2_1 _11732_ (.A0(net1121),
    .A1(_05784_),
    .S(_06106_),
    .X(_06110_));
 sky130_fd_sc_hd__clkbuf_1 _11733_ (.A(_06110_),
    .X(_01012_));
 sky130_fd_sc_hd__mux2_1 _11734_ (.A0(net130),
    .A1(_05786_),
    .S(_06106_),
    .X(_06111_));
 sky130_fd_sc_hd__clkbuf_1 _11735_ (.A(_06111_),
    .X(_01013_));
 sky130_fd_sc_hd__mux2_1 _11736_ (.A0(net1906),
    .A1(_05788_),
    .S(_06106_),
    .X(_06112_));
 sky130_fd_sc_hd__clkbuf_1 _11737_ (.A(_06112_),
    .X(_01014_));
 sky130_fd_sc_hd__mux2_1 _11738_ (.A0(net1156),
    .A1(_05790_),
    .S(_06106_),
    .X(_06113_));
 sky130_fd_sc_hd__clkbuf_1 _11739_ (.A(_06113_),
    .X(_01015_));
 sky130_fd_sc_hd__mux2_1 _11740_ (.A0(net50),
    .A1(_05792_),
    .S(_06106_),
    .X(_06114_));
 sky130_fd_sc_hd__clkbuf_1 _11741_ (.A(_06114_),
    .X(_01016_));
 sky130_fd_sc_hd__mux2_1 _11742_ (.A0(net427),
    .A1(_05794_),
    .S(_06106_),
    .X(_06115_));
 sky130_fd_sc_hd__clkbuf_1 _11743_ (.A(_06115_),
    .X(_01017_));
 sky130_fd_sc_hd__mux2_1 _11744_ (.A0(net391),
    .A1(_05796_),
    .S(_06106_),
    .X(_06116_));
 sky130_fd_sc_hd__clkbuf_1 _11745_ (.A(_06116_),
    .X(_01018_));
 sky130_fd_sc_hd__mux2_1 _11746_ (.A0(net1181),
    .A1(_05798_),
    .S(_06105_),
    .X(_06117_));
 sky130_fd_sc_hd__clkbuf_1 _11747_ (.A(_06117_),
    .X(_01019_));
 sky130_fd_sc_hd__mux2_1 _11748_ (.A0(net57),
    .A1(_05800_),
    .S(_06105_),
    .X(_06118_));
 sky130_fd_sc_hd__clkbuf_1 _11749_ (.A(_06118_),
    .X(_01020_));
 sky130_fd_sc_hd__mux2_1 _11750_ (.A0(net47),
    .A1(_05802_),
    .S(_06105_),
    .X(_06119_));
 sky130_fd_sc_hd__clkbuf_1 _11751_ (.A(_06119_),
    .X(_01021_));
 sky130_fd_sc_hd__mux2_1 _11752_ (.A0(net231),
    .A1(_05804_),
    .S(_06105_),
    .X(_06120_));
 sky130_fd_sc_hd__clkbuf_1 _11753_ (.A(_06120_),
    .X(_01022_));
 sky130_fd_sc_hd__mux2_1 _11754_ (.A0(net168),
    .A1(_05806_),
    .S(_06105_),
    .X(_06121_));
 sky130_fd_sc_hd__clkbuf_1 _11755_ (.A(_06121_),
    .X(_01023_));
 sky130_fd_sc_hd__mux2_1 _11756_ (.A0(net353),
    .A1(_05808_),
    .S(_06105_),
    .X(_06122_));
 sky130_fd_sc_hd__clkbuf_1 _11757_ (.A(_06122_),
    .X(_01024_));
 sky130_fd_sc_hd__nor2_4 _11758_ (.A(_04286_),
    .B(_04501_),
    .Y(_06123_));
 sky130_fd_sc_hd__buf_4 _11759_ (.A(_06123_),
    .X(_06124_));
 sky130_fd_sc_hd__mux2_1 _11760_ (.A0(net522),
    .A1(_05776_),
    .S(_06124_),
    .X(_06125_));
 sky130_fd_sc_hd__clkbuf_1 _11761_ (.A(_06125_),
    .X(_01025_));
 sky130_fd_sc_hd__mux2_1 _11762_ (.A0(net478),
    .A1(_05780_),
    .S(_06124_),
    .X(_06126_));
 sky130_fd_sc_hd__clkbuf_1 _11763_ (.A(_06126_),
    .X(_01026_));
 sky130_fd_sc_hd__mux2_1 _11764_ (.A0(net175),
    .A1(_05782_),
    .S(_06124_),
    .X(_06127_));
 sky130_fd_sc_hd__clkbuf_1 _11765_ (.A(_06127_),
    .X(_01027_));
 sky130_fd_sc_hd__mux2_1 _11766_ (.A0(net386),
    .A1(_05784_),
    .S(_06124_),
    .X(_06128_));
 sky130_fd_sc_hd__clkbuf_1 _11767_ (.A(_06128_),
    .X(_01028_));
 sky130_fd_sc_hd__mux2_1 _11768_ (.A0(net154),
    .A1(_05786_),
    .S(_06124_),
    .X(_06129_));
 sky130_fd_sc_hd__clkbuf_1 _11769_ (.A(_06129_),
    .X(_01029_));
 sky130_fd_sc_hd__mux2_1 _11770_ (.A0(net1456),
    .A1(_05788_),
    .S(_06124_),
    .X(_06130_));
 sky130_fd_sc_hd__clkbuf_1 _11771_ (.A(_06130_),
    .X(_01030_));
 sky130_fd_sc_hd__mux2_1 _11772_ (.A0(net431),
    .A1(_05790_),
    .S(_06124_),
    .X(_06131_));
 sky130_fd_sc_hd__clkbuf_1 _11773_ (.A(_06131_),
    .X(_01031_));
 sky130_fd_sc_hd__mux2_1 _11774_ (.A0(net861),
    .A1(_05792_),
    .S(_06124_),
    .X(_06132_));
 sky130_fd_sc_hd__clkbuf_1 _11775_ (.A(_06132_),
    .X(_01032_));
 sky130_fd_sc_hd__mux2_1 _11776_ (.A0(net710),
    .A1(_05794_),
    .S(_06124_),
    .X(_06133_));
 sky130_fd_sc_hd__clkbuf_1 _11777_ (.A(_06133_),
    .X(_01033_));
 sky130_fd_sc_hd__mux2_1 _11778_ (.A0(net251),
    .A1(_05796_),
    .S(_06124_),
    .X(_06134_));
 sky130_fd_sc_hd__clkbuf_1 _11779_ (.A(_06134_),
    .X(_01034_));
 sky130_fd_sc_hd__mux2_1 _11780_ (.A0(net1068),
    .A1(_05798_),
    .S(_06123_),
    .X(_06135_));
 sky130_fd_sc_hd__clkbuf_1 _11781_ (.A(_06135_),
    .X(_01035_));
 sky130_fd_sc_hd__mux2_1 _11782_ (.A0(net617),
    .A1(_05800_),
    .S(_06123_),
    .X(_06136_));
 sky130_fd_sc_hd__clkbuf_1 _11783_ (.A(_06136_),
    .X(_01036_));
 sky130_fd_sc_hd__mux2_1 _11784_ (.A0(net1245),
    .A1(_05802_),
    .S(_06123_),
    .X(_06137_));
 sky130_fd_sc_hd__clkbuf_1 _11785_ (.A(_06137_),
    .X(_01037_));
 sky130_fd_sc_hd__mux2_1 _11786_ (.A0(net1642),
    .A1(_05804_),
    .S(_06123_),
    .X(_06138_));
 sky130_fd_sc_hd__clkbuf_1 _11787_ (.A(_06138_),
    .X(_01038_));
 sky130_fd_sc_hd__mux2_1 _11788_ (.A0(net510),
    .A1(_05806_),
    .S(_06123_),
    .X(_06139_));
 sky130_fd_sc_hd__clkbuf_1 _11789_ (.A(_06139_),
    .X(_01039_));
 sky130_fd_sc_hd__mux2_1 _11790_ (.A0(net210),
    .A1(_05808_),
    .S(_06123_),
    .X(_06140_));
 sky130_fd_sc_hd__clkbuf_1 _11791_ (.A(_06140_),
    .X(_01040_));
 sky130_fd_sc_hd__nor2_4 _11792_ (.A(_04368_),
    .B(_04461_),
    .Y(_06141_));
 sky130_fd_sc_hd__buf_4 _11793_ (.A(_06141_),
    .X(_06142_));
 sky130_fd_sc_hd__mux2_1 _11794_ (.A0(net896),
    .A1(_05776_),
    .S(_06142_),
    .X(_06143_));
 sky130_fd_sc_hd__clkbuf_1 _11795_ (.A(_06143_),
    .X(_01041_));
 sky130_fd_sc_hd__mux2_1 _11796_ (.A0(net379),
    .A1(_05780_),
    .S(_06142_),
    .X(_06144_));
 sky130_fd_sc_hd__clkbuf_1 _11797_ (.A(_06144_),
    .X(_01042_));
 sky130_fd_sc_hd__mux2_1 _11798_ (.A0(net698),
    .A1(_05782_),
    .S(_06142_),
    .X(_06145_));
 sky130_fd_sc_hd__clkbuf_1 _11799_ (.A(_06145_),
    .X(_01043_));
 sky130_fd_sc_hd__mux2_1 _11800_ (.A0(net461),
    .A1(_05784_),
    .S(_06142_),
    .X(_06146_));
 sky130_fd_sc_hd__clkbuf_1 _11801_ (.A(_06146_),
    .X(_01044_));
 sky130_fd_sc_hd__mux2_1 _11802_ (.A0(net521),
    .A1(_05786_),
    .S(_06142_),
    .X(_06147_));
 sky130_fd_sc_hd__clkbuf_1 _11803_ (.A(_06147_),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _11804_ (.A0(net719),
    .A1(_05788_),
    .S(_06142_),
    .X(_06148_));
 sky130_fd_sc_hd__clkbuf_1 _11805_ (.A(_06148_),
    .X(_01046_));
 sky130_fd_sc_hd__mux2_1 _11806_ (.A0(net1036),
    .A1(_05790_),
    .S(_06142_),
    .X(_06149_));
 sky130_fd_sc_hd__clkbuf_1 _11807_ (.A(_06149_),
    .X(_01047_));
 sky130_fd_sc_hd__mux2_1 _11808_ (.A0(net1290),
    .A1(_05792_),
    .S(_06142_),
    .X(_06150_));
 sky130_fd_sc_hd__clkbuf_1 _11809_ (.A(_06150_),
    .X(_01048_));
 sky130_fd_sc_hd__mux2_1 _11810_ (.A0(net1620),
    .A1(_05794_),
    .S(_06142_),
    .X(_06151_));
 sky130_fd_sc_hd__clkbuf_1 _11811_ (.A(_06151_),
    .X(_01049_));
 sky130_fd_sc_hd__mux2_1 _11812_ (.A0(net938),
    .A1(_05796_),
    .S(_06142_),
    .X(_06152_));
 sky130_fd_sc_hd__clkbuf_1 _11813_ (.A(_06152_),
    .X(_01050_));
 sky130_fd_sc_hd__mux2_1 _11814_ (.A0(net682),
    .A1(_05798_),
    .S(_06141_),
    .X(_06153_));
 sky130_fd_sc_hd__clkbuf_1 _11815_ (.A(_06153_),
    .X(_01051_));
 sky130_fd_sc_hd__mux2_1 _11816_ (.A0(net1429),
    .A1(_05800_),
    .S(_06141_),
    .X(_06154_));
 sky130_fd_sc_hd__clkbuf_1 _11817_ (.A(_06154_),
    .X(_01052_));
 sky130_fd_sc_hd__mux2_1 _11818_ (.A0(net1026),
    .A1(_05802_),
    .S(_06141_),
    .X(_06155_));
 sky130_fd_sc_hd__clkbuf_1 _11819_ (.A(_06155_),
    .X(_01053_));
 sky130_fd_sc_hd__mux2_1 _11820_ (.A0(net222),
    .A1(_05804_),
    .S(_06141_),
    .X(_06156_));
 sky130_fd_sc_hd__clkbuf_1 _11821_ (.A(_06156_),
    .X(_01054_));
 sky130_fd_sc_hd__mux2_1 _11822_ (.A0(net550),
    .A1(_05806_),
    .S(_06141_),
    .X(_06157_));
 sky130_fd_sc_hd__clkbuf_1 _11823_ (.A(_06157_),
    .X(_01055_));
 sky130_fd_sc_hd__mux2_1 _11824_ (.A0(net607),
    .A1(_05808_),
    .S(_06141_),
    .X(_06158_));
 sky130_fd_sc_hd__clkbuf_1 _11825_ (.A(_06158_),
    .X(_01056_));
 sky130_fd_sc_hd__nor2_4 _11826_ (.A(_04286_),
    .B(_04569_),
    .Y(_06159_));
 sky130_fd_sc_hd__buf_4 _11827_ (.A(_06159_),
    .X(_06160_));
 sky130_fd_sc_hd__mux2_1 _11828_ (.A0(net438),
    .A1(_05776_),
    .S(_06160_),
    .X(_06161_));
 sky130_fd_sc_hd__clkbuf_1 _11829_ (.A(_06161_),
    .X(_01057_));
 sky130_fd_sc_hd__mux2_1 _11830_ (.A0(net94),
    .A1(_05780_),
    .S(_06160_),
    .X(_06162_));
 sky130_fd_sc_hd__clkbuf_1 _11831_ (.A(_06162_),
    .X(_01058_));
 sky130_fd_sc_hd__mux2_1 _11832_ (.A0(net345),
    .A1(_05782_),
    .S(_06160_),
    .X(_06163_));
 sky130_fd_sc_hd__clkbuf_1 _11833_ (.A(_06163_),
    .X(_01059_));
 sky130_fd_sc_hd__mux2_1 _11834_ (.A0(net476),
    .A1(_05784_),
    .S(_06160_),
    .X(_06164_));
 sky130_fd_sc_hd__clkbuf_1 _11835_ (.A(_06164_),
    .X(_01060_));
 sky130_fd_sc_hd__mux2_1 _11836_ (.A0(net79),
    .A1(_05786_),
    .S(_06160_),
    .X(_06165_));
 sky130_fd_sc_hd__clkbuf_1 _11837_ (.A(_06165_),
    .X(_01061_));
 sky130_fd_sc_hd__mux2_1 _11838_ (.A0(net1349),
    .A1(_05788_),
    .S(_06160_),
    .X(_06166_));
 sky130_fd_sc_hd__clkbuf_1 _11839_ (.A(_06166_),
    .X(_01062_));
 sky130_fd_sc_hd__mux2_1 _11840_ (.A0(net560),
    .A1(_05790_),
    .S(_06160_),
    .X(_06167_));
 sky130_fd_sc_hd__clkbuf_1 _11841_ (.A(_06167_),
    .X(_01063_));
 sky130_fd_sc_hd__mux2_1 _11842_ (.A0(net619),
    .A1(_05792_),
    .S(_06160_),
    .X(_06168_));
 sky130_fd_sc_hd__clkbuf_1 _11843_ (.A(_06168_),
    .X(_01064_));
 sky130_fd_sc_hd__mux2_1 _11844_ (.A0(net294),
    .A1(_05794_),
    .S(_06160_),
    .X(_06169_));
 sky130_fd_sc_hd__clkbuf_1 _11845_ (.A(_06169_),
    .X(_01065_));
 sky130_fd_sc_hd__mux2_1 _11846_ (.A0(net760),
    .A1(_05796_),
    .S(_06160_),
    .X(_06170_));
 sky130_fd_sc_hd__clkbuf_1 _11847_ (.A(_06170_),
    .X(_01066_));
 sky130_fd_sc_hd__mux2_1 _11848_ (.A0(net833),
    .A1(_05798_),
    .S(_06159_),
    .X(_06171_));
 sky130_fd_sc_hd__clkbuf_1 _11849_ (.A(_06171_),
    .X(_01067_));
 sky130_fd_sc_hd__mux2_1 _11850_ (.A0(net218),
    .A1(_05800_),
    .S(_06159_),
    .X(_06172_));
 sky130_fd_sc_hd__clkbuf_1 _11851_ (.A(_06172_),
    .X(_01068_));
 sky130_fd_sc_hd__mux2_1 _11852_ (.A0(net684),
    .A1(_05802_),
    .S(_06159_),
    .X(_06173_));
 sky130_fd_sc_hd__clkbuf_1 _11853_ (.A(_06173_),
    .X(_01069_));
 sky130_fd_sc_hd__mux2_1 _11854_ (.A0(net920),
    .A1(_05804_),
    .S(_06159_),
    .X(_06174_));
 sky130_fd_sc_hd__clkbuf_1 _11855_ (.A(_06174_),
    .X(_01070_));
 sky130_fd_sc_hd__mux2_1 _11856_ (.A0(net591),
    .A1(_05806_),
    .S(_06159_),
    .X(_06175_));
 sky130_fd_sc_hd__clkbuf_1 _11857_ (.A(_06175_),
    .X(_01071_));
 sky130_fd_sc_hd__mux2_1 _11858_ (.A0(net593),
    .A1(_05808_),
    .S(_06159_),
    .X(_06176_));
 sky130_fd_sc_hd__clkbuf_1 _11859_ (.A(_06176_),
    .X(_01072_));
 sky130_fd_sc_hd__or2_1 _11860_ (.A(_04184_),
    .B(_04285_),
    .X(_06177_));
 sky130_fd_sc_hd__clkbuf_4 _11861_ (.A(_06177_),
    .X(_06178_));
 sky130_fd_sc_hd__buf_4 _11862_ (.A(_06178_),
    .X(_06179_));
 sky130_fd_sc_hd__mux2_1 _11863_ (.A0(_05996_),
    .A1(net1561),
    .S(_06179_),
    .X(_06180_));
 sky130_fd_sc_hd__clkbuf_1 _11864_ (.A(_06180_),
    .X(_01073_));
 sky130_fd_sc_hd__mux2_1 _11865_ (.A0(_06001_),
    .A1(net1568),
    .S(_06179_),
    .X(_06181_));
 sky130_fd_sc_hd__clkbuf_1 _11866_ (.A(_06181_),
    .X(_01074_));
 sky130_fd_sc_hd__mux2_1 _11867_ (.A0(_06003_),
    .A1(net1635),
    .S(_06179_),
    .X(_06182_));
 sky130_fd_sc_hd__clkbuf_1 _11868_ (.A(_06182_),
    .X(_01075_));
 sky130_fd_sc_hd__mux2_1 _11869_ (.A0(_06005_),
    .A1(net467),
    .S(_06179_),
    .X(_06183_));
 sky130_fd_sc_hd__clkbuf_1 _11870_ (.A(_06183_),
    .X(_01076_));
 sky130_fd_sc_hd__mux2_1 _11871_ (.A0(_06007_),
    .A1(net790),
    .S(_06179_),
    .X(_06184_));
 sky130_fd_sc_hd__clkbuf_1 _11872_ (.A(_06184_),
    .X(_01077_));
 sky130_fd_sc_hd__mux2_1 _11873_ (.A0(_06009_),
    .A1(net1733),
    .S(_06179_),
    .X(_06185_));
 sky130_fd_sc_hd__clkbuf_1 _11874_ (.A(_06185_),
    .X(_01078_));
 sky130_fd_sc_hd__mux2_1 _11875_ (.A0(_06011_),
    .A1(net1964),
    .S(_06179_),
    .X(_06186_));
 sky130_fd_sc_hd__clkbuf_1 _11876_ (.A(_06186_),
    .X(_01079_));
 sky130_fd_sc_hd__mux2_1 _11877_ (.A0(_06013_),
    .A1(net1374),
    .S(_06179_),
    .X(_06187_));
 sky130_fd_sc_hd__clkbuf_1 _11878_ (.A(_06187_),
    .X(_01080_));
 sky130_fd_sc_hd__mux2_1 _11879_ (.A0(_06015_),
    .A1(net1187),
    .S(_06179_),
    .X(_06188_));
 sky130_fd_sc_hd__clkbuf_1 _11880_ (.A(_06188_),
    .X(_01081_));
 sky130_fd_sc_hd__mux2_1 _11881_ (.A0(_06017_),
    .A1(net662),
    .S(_06179_),
    .X(_06189_));
 sky130_fd_sc_hd__clkbuf_1 _11882_ (.A(_06189_),
    .X(_01082_));
 sky130_fd_sc_hd__mux2_1 _11883_ (.A0(_06019_),
    .A1(net1278),
    .S(_06178_),
    .X(_06190_));
 sky130_fd_sc_hd__clkbuf_1 _11884_ (.A(_06190_),
    .X(_01083_));
 sky130_fd_sc_hd__mux2_1 _11885_ (.A0(_06021_),
    .A1(net600),
    .S(_06178_),
    .X(_06191_));
 sky130_fd_sc_hd__clkbuf_1 _11886_ (.A(_06191_),
    .X(_01084_));
 sky130_fd_sc_hd__mux2_1 _11887_ (.A0(_06023_),
    .A1(net1280),
    .S(_06178_),
    .X(_06192_));
 sky130_fd_sc_hd__clkbuf_1 _11888_ (.A(_06192_),
    .X(_01085_));
 sky130_fd_sc_hd__mux2_1 _11889_ (.A0(_06025_),
    .A1(net611),
    .S(_06178_),
    .X(_06193_));
 sky130_fd_sc_hd__clkbuf_1 _11890_ (.A(_06193_),
    .X(_01086_));
 sky130_fd_sc_hd__mux2_1 _11891_ (.A0(_06027_),
    .A1(net854),
    .S(_06178_),
    .X(_06194_));
 sky130_fd_sc_hd__clkbuf_1 _11892_ (.A(_06194_),
    .X(_01087_));
 sky130_fd_sc_hd__mux2_1 _11893_ (.A0(_06029_),
    .A1(net962),
    .S(_06178_),
    .X(_06195_));
 sky130_fd_sc_hd__clkbuf_1 _11894_ (.A(_06195_),
    .X(_01088_));
 sky130_fd_sc_hd__or2_1 _11895_ (.A(_04286_),
    .B(_04607_),
    .X(_06196_));
 sky130_fd_sc_hd__clkbuf_4 _11896_ (.A(_06196_),
    .X(_06197_));
 sky130_fd_sc_hd__buf_4 _11897_ (.A(_06197_),
    .X(_06198_));
 sky130_fd_sc_hd__mux2_1 _11898_ (.A0(_05996_),
    .A1(net310),
    .S(_06198_),
    .X(_06199_));
 sky130_fd_sc_hd__clkbuf_1 _11899_ (.A(_06199_),
    .X(_01089_));
 sky130_fd_sc_hd__mux2_1 _11900_ (.A0(_06001_),
    .A1(net1631),
    .S(_06198_),
    .X(_06200_));
 sky130_fd_sc_hd__clkbuf_1 _11901_ (.A(_06200_),
    .X(_01090_));
 sky130_fd_sc_hd__mux2_1 _11902_ (.A0(_06003_),
    .A1(net278),
    .S(_06198_),
    .X(_06201_));
 sky130_fd_sc_hd__clkbuf_1 _11903_ (.A(_06201_),
    .X(_01091_));
 sky130_fd_sc_hd__mux2_1 _11904_ (.A0(_06005_),
    .A1(net1463),
    .S(_06198_),
    .X(_06202_));
 sky130_fd_sc_hd__clkbuf_1 _11905_ (.A(_06202_),
    .X(_01092_));
 sky130_fd_sc_hd__mux2_1 _11906_ (.A0(_06007_),
    .A1(net1000),
    .S(_06198_),
    .X(_06203_));
 sky130_fd_sc_hd__clkbuf_1 _11907_ (.A(_06203_),
    .X(_01093_));
 sky130_fd_sc_hd__mux2_1 _11908_ (.A0(_06009_),
    .A1(net1694),
    .S(_06198_),
    .X(_06204_));
 sky130_fd_sc_hd__clkbuf_1 _11909_ (.A(_06204_),
    .X(_01094_));
 sky130_fd_sc_hd__mux2_1 _11910_ (.A0(_06011_),
    .A1(net1600),
    .S(_06198_),
    .X(_06205_));
 sky130_fd_sc_hd__clkbuf_1 _11911_ (.A(_06205_),
    .X(_01095_));
 sky130_fd_sc_hd__mux2_1 _11912_ (.A0(_06013_),
    .A1(net445),
    .S(_06198_),
    .X(_06206_));
 sky130_fd_sc_hd__clkbuf_1 _11913_ (.A(_06206_),
    .X(_01096_));
 sky130_fd_sc_hd__mux2_1 _11914_ (.A0(_06015_),
    .A1(net1142),
    .S(_06198_),
    .X(_06207_));
 sky130_fd_sc_hd__clkbuf_1 _11915_ (.A(_06207_),
    .X(_01097_));
 sky130_fd_sc_hd__mux2_1 _11916_ (.A0(_06017_),
    .A1(net1566),
    .S(_06198_),
    .X(_06208_));
 sky130_fd_sc_hd__clkbuf_1 _11917_ (.A(_06208_),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_1 _11918_ (.A0(_06019_),
    .A1(net754),
    .S(_06197_),
    .X(_06209_));
 sky130_fd_sc_hd__clkbuf_1 _11919_ (.A(_06209_),
    .X(_01099_));
 sky130_fd_sc_hd__mux2_1 _11920_ (.A0(_06021_),
    .A1(net1098),
    .S(_06197_),
    .X(_06210_));
 sky130_fd_sc_hd__clkbuf_1 _11921_ (.A(_06210_),
    .X(_01100_));
 sky130_fd_sc_hd__mux2_1 _11922_ (.A0(_06023_),
    .A1(net701),
    .S(_06197_),
    .X(_06211_));
 sky130_fd_sc_hd__clkbuf_1 _11923_ (.A(_06211_),
    .X(_01101_));
 sky130_fd_sc_hd__mux2_1 _11924_ (.A0(_06025_),
    .A1(net881),
    .S(_06197_),
    .X(_06212_));
 sky130_fd_sc_hd__clkbuf_1 _11925_ (.A(_06212_),
    .X(_01102_));
 sky130_fd_sc_hd__mux2_1 _11926_ (.A0(_06027_),
    .A1(net1574),
    .S(_06197_),
    .X(_06213_));
 sky130_fd_sc_hd__clkbuf_1 _11927_ (.A(_06213_),
    .X(_01103_));
 sky130_fd_sc_hd__mux2_1 _11928_ (.A0(_06029_),
    .A1(net1080),
    .S(_06197_),
    .X(_06214_));
 sky130_fd_sc_hd__clkbuf_1 _11929_ (.A(_06214_),
    .X(_01104_));
 sky130_fd_sc_hd__or3_1 _11930_ (.A(_02498_),
    .B(_02644_),
    .C(_04285_),
    .X(_06215_));
 sky130_fd_sc_hd__clkbuf_4 _11931_ (.A(_06215_),
    .X(_06216_));
 sky130_fd_sc_hd__buf_4 _11932_ (.A(_06216_),
    .X(_06217_));
 sky130_fd_sc_hd__mux2_1 _11933_ (.A0(_05996_),
    .A1(net984),
    .S(_06217_),
    .X(_06218_));
 sky130_fd_sc_hd__clkbuf_1 _11934_ (.A(_06218_),
    .X(_01105_));
 sky130_fd_sc_hd__mux2_1 _11935_ (.A0(_06001_),
    .A1(net1030),
    .S(_06217_),
    .X(_06219_));
 sky130_fd_sc_hd__clkbuf_1 _11936_ (.A(_06219_),
    .X(_01106_));
 sky130_fd_sc_hd__mux2_1 _11937_ (.A0(_06003_),
    .A1(net383),
    .S(_06217_),
    .X(_06220_));
 sky130_fd_sc_hd__clkbuf_1 _11938_ (.A(_06220_),
    .X(_01107_));
 sky130_fd_sc_hd__mux2_1 _11939_ (.A0(_06005_),
    .A1(net1282),
    .S(_06217_),
    .X(_06221_));
 sky130_fd_sc_hd__clkbuf_1 _11940_ (.A(_06221_),
    .X(_01108_));
 sky130_fd_sc_hd__mux2_1 _11941_ (.A0(_06007_),
    .A1(net884),
    .S(_06217_),
    .X(_06222_));
 sky130_fd_sc_hd__clkbuf_1 _11942_ (.A(_06222_),
    .X(_01109_));
 sky130_fd_sc_hd__mux2_1 _11943_ (.A0(_06009_),
    .A1(net964),
    .S(_06217_),
    .X(_06223_));
 sky130_fd_sc_hd__clkbuf_1 _11944_ (.A(_06223_),
    .X(_01110_));
 sky130_fd_sc_hd__mux2_1 _11945_ (.A0(_06011_),
    .A1(net505),
    .S(_06217_),
    .X(_06224_));
 sky130_fd_sc_hd__clkbuf_1 _11946_ (.A(_06224_),
    .X(_01111_));
 sky130_fd_sc_hd__mux2_1 _11947_ (.A0(_06013_),
    .A1(net1144),
    .S(_06217_),
    .X(_06225_));
 sky130_fd_sc_hd__clkbuf_1 _11948_ (.A(_06225_),
    .X(_01112_));
 sky130_fd_sc_hd__mux2_1 _11949_ (.A0(_06015_),
    .A1(net1323),
    .S(_06217_),
    .X(_06226_));
 sky130_fd_sc_hd__clkbuf_1 _11950_ (.A(_06226_),
    .X(_01113_));
 sky130_fd_sc_hd__mux2_1 _11951_ (.A0(_06017_),
    .A1(net1242),
    .S(_06217_),
    .X(_06227_));
 sky130_fd_sc_hd__clkbuf_1 _11952_ (.A(_06227_),
    .X(_01114_));
 sky130_fd_sc_hd__mux2_1 _11953_ (.A0(_06019_),
    .A1(net869),
    .S(_06216_),
    .X(_06228_));
 sky130_fd_sc_hd__clkbuf_1 _11954_ (.A(_06228_),
    .X(_01115_));
 sky130_fd_sc_hd__mux2_1 _11955_ (.A0(_06021_),
    .A1(net1401),
    .S(_06216_),
    .X(_06229_));
 sky130_fd_sc_hd__clkbuf_1 _11956_ (.A(_06229_),
    .X(_01116_));
 sky130_fd_sc_hd__mux2_1 _11957_ (.A0(_06023_),
    .A1(net931),
    .S(_06216_),
    .X(_06230_));
 sky130_fd_sc_hd__clkbuf_1 _11958_ (.A(_06230_),
    .X(_01117_));
 sky130_fd_sc_hd__mux2_1 _11959_ (.A0(_06025_),
    .A1(net823),
    .S(_06216_),
    .X(_06231_));
 sky130_fd_sc_hd__clkbuf_1 _11960_ (.A(_06231_),
    .X(_01118_));
 sky130_fd_sc_hd__mux2_1 _11961_ (.A0(_06027_),
    .A1(net702),
    .S(_06216_),
    .X(_06232_));
 sky130_fd_sc_hd__clkbuf_1 _11962_ (.A(_06232_),
    .X(_01119_));
 sky130_fd_sc_hd__mux2_1 _11963_ (.A0(_06029_),
    .A1(net777),
    .S(_06216_),
    .X(_06233_));
 sky130_fd_sc_hd__clkbuf_1 _11964_ (.A(_06233_),
    .X(_01120_));
 sky130_fd_sc_hd__nor2_4 _11965_ (.A(_04286_),
    .B(_04646_),
    .Y(_06234_));
 sky130_fd_sc_hd__buf_4 _11966_ (.A(_06234_),
    .X(_06235_));
 sky130_fd_sc_hd__mux2_1 _11967_ (.A0(net2031),
    .A1(_04498_),
    .S(_06235_),
    .X(_06236_));
 sky130_fd_sc_hd__clkbuf_1 _11968_ (.A(_06236_),
    .X(_01121_));
 sky130_fd_sc_hd__mux2_1 _11969_ (.A0(net312),
    .A1(_04505_),
    .S(_06235_),
    .X(_06237_));
 sky130_fd_sc_hd__clkbuf_1 _11970_ (.A(_06237_),
    .X(_01122_));
 sky130_fd_sc_hd__mux2_1 _11971_ (.A0(net2044),
    .A1(_04508_),
    .S(_06235_),
    .X(_06238_));
 sky130_fd_sc_hd__clkbuf_1 _11972_ (.A(_06238_),
    .X(_01123_));
 sky130_fd_sc_hd__mux2_1 _11973_ (.A0(net1363),
    .A1(_04511_),
    .S(_06235_),
    .X(_06239_));
 sky130_fd_sc_hd__clkbuf_1 _11974_ (.A(_06239_),
    .X(_01124_));
 sky130_fd_sc_hd__mux2_1 _11975_ (.A0(net131),
    .A1(_04514_),
    .S(_06235_),
    .X(_06240_));
 sky130_fd_sc_hd__clkbuf_1 _11976_ (.A(_06240_),
    .X(_01125_));
 sky130_fd_sc_hd__mux2_1 _11977_ (.A0(net97),
    .A1(_04517_),
    .S(_06235_),
    .X(_06241_));
 sky130_fd_sc_hd__clkbuf_1 _11978_ (.A(_06241_),
    .X(_01126_));
 sky130_fd_sc_hd__mux2_1 _11979_ (.A0(net1549),
    .A1(_04520_),
    .S(_06235_),
    .X(_06242_));
 sky130_fd_sc_hd__clkbuf_1 _11980_ (.A(_06242_),
    .X(_01127_));
 sky130_fd_sc_hd__mux2_1 _11981_ (.A0(net1866),
    .A1(_04523_),
    .S(_06235_),
    .X(_06243_));
 sky130_fd_sc_hd__clkbuf_1 _11982_ (.A(_06243_),
    .X(_01128_));
 sky130_fd_sc_hd__mux2_1 _11983_ (.A0(net1921),
    .A1(_04526_),
    .S(_06235_),
    .X(_06244_));
 sky130_fd_sc_hd__clkbuf_1 _11984_ (.A(_06244_),
    .X(_01129_));
 sky130_fd_sc_hd__mux2_1 _11985_ (.A0(net643),
    .A1(_04529_),
    .S(_06235_),
    .X(_06245_));
 sky130_fd_sc_hd__clkbuf_1 _11986_ (.A(_06245_),
    .X(_01130_));
 sky130_fd_sc_hd__mux2_1 _11987_ (.A0(net1332),
    .A1(_04532_),
    .S(_06234_),
    .X(_06246_));
 sky130_fd_sc_hd__clkbuf_1 _11988_ (.A(_06246_),
    .X(_01131_));
 sky130_fd_sc_hd__mux2_1 _11989_ (.A0(net313),
    .A1(_04535_),
    .S(_06234_),
    .X(_06247_));
 sky130_fd_sc_hd__clkbuf_1 _11990_ (.A(_06247_),
    .X(_01132_));
 sky130_fd_sc_hd__mux2_1 _11991_ (.A0(net1067),
    .A1(_04538_),
    .S(_06234_),
    .X(_06248_));
 sky130_fd_sc_hd__clkbuf_1 _11992_ (.A(_06248_),
    .X(_01133_));
 sky130_fd_sc_hd__mux2_1 _11993_ (.A0(net1936),
    .A1(_04541_),
    .S(_06234_),
    .X(_06249_));
 sky130_fd_sc_hd__clkbuf_1 _11994_ (.A(_06249_),
    .X(_01134_));
 sky130_fd_sc_hd__mux2_1 _11995_ (.A0(net1724),
    .A1(_04544_),
    .S(_06234_),
    .X(_06250_));
 sky130_fd_sc_hd__clkbuf_1 _11996_ (.A(_06250_),
    .X(_01135_));
 sky130_fd_sc_hd__mux2_1 _11997_ (.A0(net2041),
    .A1(_04547_),
    .S(_06234_),
    .X(_06251_));
 sky130_fd_sc_hd__clkbuf_1 _11998_ (.A(_06251_),
    .X(_01136_));
 sky130_fd_sc_hd__or2_1 _11999_ (.A(_04127_),
    .B(_04285_),
    .X(_06252_));
 sky130_fd_sc_hd__clkbuf_4 _12000_ (.A(_06252_),
    .X(_06253_));
 sky130_fd_sc_hd__buf_4 _12001_ (.A(_06253_),
    .X(_06254_));
 sky130_fd_sc_hd__mux2_1 _12002_ (.A0(_05996_),
    .A1(net645),
    .S(_06254_),
    .X(_06255_));
 sky130_fd_sc_hd__clkbuf_1 _12003_ (.A(_06255_),
    .X(_01137_));
 sky130_fd_sc_hd__mux2_1 _12004_ (.A0(_06001_),
    .A1(net1143),
    .S(_06254_),
    .X(_06256_));
 sky130_fd_sc_hd__clkbuf_1 _12005_ (.A(_06256_),
    .X(_01138_));
 sky130_fd_sc_hd__mux2_1 _12006_ (.A0(_06003_),
    .A1(net1007),
    .S(_06254_),
    .X(_06257_));
 sky130_fd_sc_hd__clkbuf_1 _12007_ (.A(_06257_),
    .X(_01139_));
 sky130_fd_sc_hd__mux2_1 _12008_ (.A0(_06005_),
    .A1(net1503),
    .S(_06254_),
    .X(_06258_));
 sky130_fd_sc_hd__clkbuf_1 _12009_ (.A(_06258_),
    .X(_01140_));
 sky130_fd_sc_hd__mux2_1 _12010_ (.A0(_06007_),
    .A1(net1563),
    .S(_06254_),
    .X(_06259_));
 sky130_fd_sc_hd__clkbuf_1 _12011_ (.A(_06259_),
    .X(_01141_));
 sky130_fd_sc_hd__mux2_1 _12012_ (.A0(_06009_),
    .A1(net325),
    .S(_06254_),
    .X(_06260_));
 sky130_fd_sc_hd__clkbuf_1 _12013_ (.A(_06260_),
    .X(_01142_));
 sky130_fd_sc_hd__mux2_1 _12014_ (.A0(_06011_),
    .A1(net972),
    .S(_06254_),
    .X(_06261_));
 sky130_fd_sc_hd__clkbuf_1 _12015_ (.A(_06261_),
    .X(_01143_));
 sky130_fd_sc_hd__mux2_1 _12016_ (.A0(_06013_),
    .A1(net1256),
    .S(_06254_),
    .X(_06262_));
 sky130_fd_sc_hd__clkbuf_1 _12017_ (.A(_06262_),
    .X(_01144_));
 sky130_fd_sc_hd__mux2_1 _12018_ (.A0(_06015_),
    .A1(net1338),
    .S(_06254_),
    .X(_06263_));
 sky130_fd_sc_hd__clkbuf_1 _12019_ (.A(_06263_),
    .X(_01145_));
 sky130_fd_sc_hd__mux2_1 _12020_ (.A0(_06017_),
    .A1(net891),
    .S(_06254_),
    .X(_06264_));
 sky130_fd_sc_hd__clkbuf_1 _12021_ (.A(_06264_),
    .X(_01146_));
 sky130_fd_sc_hd__mux2_1 _12022_ (.A0(_06019_),
    .A1(net1095),
    .S(_06253_),
    .X(_06265_));
 sky130_fd_sc_hd__clkbuf_1 _12023_ (.A(_06265_),
    .X(_01147_));
 sky130_fd_sc_hd__mux2_1 _12024_ (.A0(_06021_),
    .A1(net486),
    .S(_06253_),
    .X(_06266_));
 sky130_fd_sc_hd__clkbuf_1 _12025_ (.A(_06266_),
    .X(_01148_));
 sky130_fd_sc_hd__mux2_1 _12026_ (.A0(_06023_),
    .A1(net842),
    .S(_06253_),
    .X(_06267_));
 sky130_fd_sc_hd__clkbuf_1 _12027_ (.A(_06267_),
    .X(_01149_));
 sky130_fd_sc_hd__mux2_1 _12028_ (.A0(_06025_),
    .A1(net1206),
    .S(_06253_),
    .X(_06268_));
 sky130_fd_sc_hd__clkbuf_1 _12029_ (.A(_06268_),
    .X(_01150_));
 sky130_fd_sc_hd__mux2_1 _12030_ (.A0(_06027_),
    .A1(net214),
    .S(_06253_),
    .X(_06269_));
 sky130_fd_sc_hd__clkbuf_1 _12031_ (.A(_06269_),
    .X(_01151_));
 sky130_fd_sc_hd__mux2_1 _12032_ (.A0(_06029_),
    .A1(net797),
    .S(_06253_),
    .X(_06270_));
 sky130_fd_sc_hd__clkbuf_1 _12033_ (.A(_06270_),
    .X(_01152_));
 sky130_fd_sc_hd__or2_1 _12034_ (.A(_04286_),
    .B(_04684_),
    .X(_06271_));
 sky130_fd_sc_hd__buf_2 _12035_ (.A(_06271_),
    .X(_06272_));
 sky130_fd_sc_hd__buf_4 _12036_ (.A(_06272_),
    .X(_06273_));
 sky130_fd_sc_hd__mux2_1 _12037_ (.A0(_05996_),
    .A1(net1638),
    .S(_06273_),
    .X(_06274_));
 sky130_fd_sc_hd__clkbuf_1 _12038_ (.A(_06274_),
    .X(_01153_));
 sky130_fd_sc_hd__mux2_1 _12039_ (.A0(_06001_),
    .A1(net319),
    .S(_06273_),
    .X(_06275_));
 sky130_fd_sc_hd__clkbuf_1 _12040_ (.A(_06275_),
    .X(_01154_));
 sky130_fd_sc_hd__mux2_1 _12041_ (.A0(_06003_),
    .A1(net1408),
    .S(_06273_),
    .X(_06276_));
 sky130_fd_sc_hd__clkbuf_1 _12042_ (.A(_06276_),
    .X(_01155_));
 sky130_fd_sc_hd__mux2_1 _12043_ (.A0(_06005_),
    .A1(net625),
    .S(_06273_),
    .X(_06277_));
 sky130_fd_sc_hd__clkbuf_1 _12044_ (.A(_06277_),
    .X(_01156_));
 sky130_fd_sc_hd__mux2_1 _12045_ (.A0(_06007_),
    .A1(net1912),
    .S(_06273_),
    .X(_06278_));
 sky130_fd_sc_hd__clkbuf_1 _12046_ (.A(_06278_),
    .X(_01157_));
 sky130_fd_sc_hd__mux2_1 _12047_ (.A0(_06009_),
    .A1(net257),
    .S(_06273_),
    .X(_06279_));
 sky130_fd_sc_hd__clkbuf_1 _12048_ (.A(_06279_),
    .X(_01158_));
 sky130_fd_sc_hd__mux2_1 _12049_ (.A0(_06011_),
    .A1(net1160),
    .S(_06273_),
    .X(_06280_));
 sky130_fd_sc_hd__clkbuf_1 _12050_ (.A(_06280_),
    .X(_01159_));
 sky130_fd_sc_hd__mux2_1 _12051_ (.A0(_06013_),
    .A1(net1346),
    .S(_06273_),
    .X(_06281_));
 sky130_fd_sc_hd__clkbuf_1 _12052_ (.A(_06281_),
    .X(_01160_));
 sky130_fd_sc_hd__mux2_1 _12053_ (.A0(_06015_),
    .A1(net1415),
    .S(_06273_),
    .X(_06282_));
 sky130_fd_sc_hd__clkbuf_1 _12054_ (.A(_06282_),
    .X(_01161_));
 sky130_fd_sc_hd__mux2_1 _12055_ (.A0(_06017_),
    .A1(net707),
    .S(_06273_),
    .X(_06283_));
 sky130_fd_sc_hd__clkbuf_1 _12056_ (.A(_06283_),
    .X(_01162_));
 sky130_fd_sc_hd__mux2_1 _12057_ (.A0(_06019_),
    .A1(net1070),
    .S(_06272_),
    .X(_06284_));
 sky130_fd_sc_hd__clkbuf_1 _12058_ (.A(_06284_),
    .X(_01163_));
 sky130_fd_sc_hd__mux2_1 _12059_ (.A0(_06021_),
    .A1(net877),
    .S(_06272_),
    .X(_06285_));
 sky130_fd_sc_hd__clkbuf_1 _12060_ (.A(_06285_),
    .X(_01164_));
 sky130_fd_sc_hd__mux2_1 _12061_ (.A0(_06023_),
    .A1(net564),
    .S(_06272_),
    .X(_06286_));
 sky130_fd_sc_hd__clkbuf_1 _12062_ (.A(_06286_),
    .X(_01165_));
 sky130_fd_sc_hd__mux2_1 _12063_ (.A0(_06025_),
    .A1(net1529),
    .S(_06272_),
    .X(_06287_));
 sky130_fd_sc_hd__clkbuf_1 _12064_ (.A(_06287_),
    .X(_01166_));
 sky130_fd_sc_hd__mux2_1 _12065_ (.A0(_06027_),
    .A1(net1224),
    .S(_06272_),
    .X(_06288_));
 sky130_fd_sc_hd__clkbuf_1 _12066_ (.A(_06288_),
    .X(_01167_));
 sky130_fd_sc_hd__mux2_1 _12067_ (.A0(_06029_),
    .A1(net1039),
    .S(_06272_),
    .X(_06289_));
 sky130_fd_sc_hd__clkbuf_1 _12068_ (.A(_06289_),
    .X(_01168_));
 sky130_fd_sc_hd__or3_1 _12069_ (.A(_02506_),
    .B(_02644_),
    .C(_04285_),
    .X(_06290_));
 sky130_fd_sc_hd__clkbuf_4 _12070_ (.A(_06290_),
    .X(_06291_));
 sky130_fd_sc_hd__buf_4 _12071_ (.A(_06291_),
    .X(_06292_));
 sky130_fd_sc_hd__mux2_1 _12072_ (.A0(_05996_),
    .A1(net1309),
    .S(_06292_),
    .X(_06293_));
 sky130_fd_sc_hd__clkbuf_1 _12073_ (.A(_06293_),
    .X(_01169_));
 sky130_fd_sc_hd__mux2_1 _12074_ (.A0(_06001_),
    .A1(net494),
    .S(_06292_),
    .X(_06294_));
 sky130_fd_sc_hd__clkbuf_1 _12075_ (.A(_06294_),
    .X(_01170_));
 sky130_fd_sc_hd__mux2_1 _12076_ (.A0(_06003_),
    .A1(net1016),
    .S(_06292_),
    .X(_06295_));
 sky130_fd_sc_hd__clkbuf_1 _12077_ (.A(_06295_),
    .X(_01171_));
 sky130_fd_sc_hd__mux2_1 _12078_ (.A0(_06005_),
    .A1(net697),
    .S(_06292_),
    .X(_06296_));
 sky130_fd_sc_hd__clkbuf_1 _12079_ (.A(_06296_),
    .X(_01172_));
 sky130_fd_sc_hd__mux2_1 _12080_ (.A0(_06007_),
    .A1(net421),
    .S(_06292_),
    .X(_06297_));
 sky130_fd_sc_hd__clkbuf_1 _12081_ (.A(_06297_),
    .X(_01173_));
 sky130_fd_sc_hd__mux2_1 _12082_ (.A0(_06009_),
    .A1(net545),
    .S(_06292_),
    .X(_06298_));
 sky130_fd_sc_hd__clkbuf_1 _12083_ (.A(_06298_),
    .X(_01174_));
 sky130_fd_sc_hd__mux2_1 _12084_ (.A0(_06011_),
    .A1(net918),
    .S(_06292_),
    .X(_06299_));
 sky130_fd_sc_hd__clkbuf_1 _12085_ (.A(_06299_),
    .X(_01175_));
 sky130_fd_sc_hd__mux2_1 _12086_ (.A0(_06013_),
    .A1(net900),
    .S(_06292_),
    .X(_06300_));
 sky130_fd_sc_hd__clkbuf_1 _12087_ (.A(_06300_),
    .X(_01176_));
 sky130_fd_sc_hd__mux2_1 _12088_ (.A0(_06015_),
    .A1(net1198),
    .S(_06292_),
    .X(_06301_));
 sky130_fd_sc_hd__clkbuf_1 _12089_ (.A(_06301_),
    .X(_01177_));
 sky130_fd_sc_hd__mux2_1 _12090_ (.A0(_06017_),
    .A1(net586),
    .S(_06292_),
    .X(_06302_));
 sky130_fd_sc_hd__clkbuf_1 _12091_ (.A(_06302_),
    .X(_01178_));
 sky130_fd_sc_hd__mux2_1 _12092_ (.A0(_06019_),
    .A1(net784),
    .S(_06291_),
    .X(_06303_));
 sky130_fd_sc_hd__clkbuf_1 _12093_ (.A(_06303_),
    .X(_01179_));
 sky130_fd_sc_hd__mux2_1 _12094_ (.A0(_06021_),
    .A1(net627),
    .S(_06291_),
    .X(_06304_));
 sky130_fd_sc_hd__clkbuf_1 _12095_ (.A(_06304_),
    .X(_01180_));
 sky130_fd_sc_hd__mux2_1 _12096_ (.A0(_06023_),
    .A1(net537),
    .S(_06291_),
    .X(_06305_));
 sky130_fd_sc_hd__clkbuf_1 _12097_ (.A(_06305_),
    .X(_01181_));
 sky130_fd_sc_hd__mux2_1 _12098_ (.A0(_06025_),
    .A1(net1326),
    .S(_06291_),
    .X(_06306_));
 sky130_fd_sc_hd__clkbuf_1 _12099_ (.A(_06306_),
    .X(_01182_));
 sky130_fd_sc_hd__mux2_1 _12100_ (.A0(_06027_),
    .A1(net1409),
    .S(_06291_),
    .X(_06307_));
 sky130_fd_sc_hd__clkbuf_1 _12101_ (.A(_06307_),
    .X(_01183_));
 sky130_fd_sc_hd__mux2_1 _12102_ (.A0(_06029_),
    .A1(net1304),
    .S(_06291_),
    .X(_06308_));
 sky130_fd_sc_hd__clkbuf_1 _12103_ (.A(_06308_),
    .X(_01184_));
 sky130_fd_sc_hd__buf_6 _12104_ (.A(_04069_),
    .X(_06309_));
 sky130_fd_sc_hd__or2_1 _12105_ (.A(_04286_),
    .B(_04365_),
    .X(_06310_));
 sky130_fd_sc_hd__buf_2 _12106_ (.A(_06310_),
    .X(_06311_));
 sky130_fd_sc_hd__buf_4 _12107_ (.A(_06311_),
    .X(_06312_));
 sky130_fd_sc_hd__mux2_1 _12108_ (.A0(_06309_),
    .A1(net1540),
    .S(_06312_),
    .X(_06313_));
 sky130_fd_sc_hd__clkbuf_1 _12109_ (.A(_06313_),
    .X(_01185_));
 sky130_fd_sc_hd__clkbuf_4 _12110_ (.A(_04080_),
    .X(_06314_));
 sky130_fd_sc_hd__mux2_1 _12111_ (.A0(_06314_),
    .A1(net1235),
    .S(_06312_),
    .X(_06315_));
 sky130_fd_sc_hd__clkbuf_1 _12112_ (.A(_06315_),
    .X(_01186_));
 sky130_fd_sc_hd__clkbuf_8 _12113_ (.A(_04083_),
    .X(_06316_));
 sky130_fd_sc_hd__mux2_1 _12114_ (.A0(_06316_),
    .A1(net1244),
    .S(_06312_),
    .X(_06317_));
 sky130_fd_sc_hd__clkbuf_1 _12115_ (.A(_06317_),
    .X(_01187_));
 sky130_fd_sc_hd__buf_4 _12116_ (.A(_04086_),
    .X(_06318_));
 sky130_fd_sc_hd__mux2_1 _12117_ (.A0(_06318_),
    .A1(net965),
    .S(_06312_),
    .X(_06319_));
 sky130_fd_sc_hd__clkbuf_1 _12118_ (.A(_06319_),
    .X(_01188_));
 sky130_fd_sc_hd__buf_4 _12119_ (.A(_04089_),
    .X(_06320_));
 sky130_fd_sc_hd__mux2_1 _12120_ (.A0(_06320_),
    .A1(net1281),
    .S(_06312_),
    .X(_06321_));
 sky130_fd_sc_hd__clkbuf_1 _12121_ (.A(_06321_),
    .X(_01189_));
 sky130_fd_sc_hd__clkbuf_4 _12122_ (.A(_04092_),
    .X(_06322_));
 sky130_fd_sc_hd__mux2_1 _12123_ (.A0(_06322_),
    .A1(net688),
    .S(_06312_),
    .X(_06323_));
 sky130_fd_sc_hd__clkbuf_1 _12124_ (.A(_06323_),
    .X(_01190_));
 sky130_fd_sc_hd__buf_4 _12125_ (.A(_04095_),
    .X(_06324_));
 sky130_fd_sc_hd__mux2_1 _12126_ (.A0(_06324_),
    .A1(net2013),
    .S(_06312_),
    .X(_06325_));
 sky130_fd_sc_hd__clkbuf_1 _12127_ (.A(_06325_),
    .X(_01191_));
 sky130_fd_sc_hd__buf_4 _12128_ (.A(_04098_),
    .X(_06326_));
 sky130_fd_sc_hd__mux2_1 _12129_ (.A0(_06326_),
    .A1(net693),
    .S(_06312_),
    .X(_06327_));
 sky130_fd_sc_hd__clkbuf_1 _12130_ (.A(_06327_),
    .X(_01192_));
 sky130_fd_sc_hd__buf_4 _12131_ (.A(_04101_),
    .X(_06328_));
 sky130_fd_sc_hd__mux2_1 _12132_ (.A0(_06328_),
    .A1(net332),
    .S(_06312_),
    .X(_06329_));
 sky130_fd_sc_hd__clkbuf_1 _12133_ (.A(_06329_),
    .X(_01193_));
 sky130_fd_sc_hd__buf_4 _12134_ (.A(_04104_),
    .X(_06330_));
 sky130_fd_sc_hd__mux2_1 _12135_ (.A0(_06330_),
    .A1(net847),
    .S(_06312_),
    .X(_06331_));
 sky130_fd_sc_hd__clkbuf_1 _12136_ (.A(_06331_),
    .X(_01194_));
 sky130_fd_sc_hd__buf_6 _12137_ (.A(_04107_),
    .X(_06332_));
 sky130_fd_sc_hd__mux2_1 _12138_ (.A0(_06332_),
    .A1(net1955),
    .S(_06311_),
    .X(_06333_));
 sky130_fd_sc_hd__clkbuf_1 _12139_ (.A(_06333_),
    .X(_01195_));
 sky130_fd_sc_hd__buf_4 _12140_ (.A(_04110_),
    .X(_06334_));
 sky130_fd_sc_hd__mux2_1 _12141_ (.A0(_06334_),
    .A1(net1846),
    .S(_06311_),
    .X(_06335_));
 sky130_fd_sc_hd__clkbuf_1 _12142_ (.A(_06335_),
    .X(_01196_));
 sky130_fd_sc_hd__clkbuf_8 _12143_ (.A(_04113_),
    .X(_06336_));
 sky130_fd_sc_hd__mux2_1 _12144_ (.A0(_06336_),
    .A1(net1287),
    .S(_06311_),
    .X(_06337_));
 sky130_fd_sc_hd__clkbuf_1 _12145_ (.A(_06337_),
    .X(_01197_));
 sky130_fd_sc_hd__clkbuf_4 _12146_ (.A(_04116_),
    .X(_06338_));
 sky130_fd_sc_hd__mux2_1 _12147_ (.A0(_06338_),
    .A1(net596),
    .S(_06311_),
    .X(_06339_));
 sky130_fd_sc_hd__clkbuf_1 _12148_ (.A(_06339_),
    .X(_01198_));
 sky130_fd_sc_hd__buf_6 _12149_ (.A(_04119_),
    .X(_06340_));
 sky130_fd_sc_hd__mux2_1 _12150_ (.A0(_06340_),
    .A1(net1193),
    .S(_06311_),
    .X(_06341_));
 sky130_fd_sc_hd__clkbuf_1 _12151_ (.A(_06341_),
    .X(_01199_));
 sky130_fd_sc_hd__buf_4 _12152_ (.A(_04122_),
    .X(_06342_));
 sky130_fd_sc_hd__mux2_1 _12153_ (.A0(_06342_),
    .A1(net935),
    .S(_06311_),
    .X(_06343_));
 sky130_fd_sc_hd__clkbuf_1 _12154_ (.A(_06343_),
    .X(_01200_));
 sky130_fd_sc_hd__nor2_4 _12155_ (.A(_04367_),
    .B(_04684_),
    .Y(_06344_));
 sky130_fd_sc_hd__buf_4 _12156_ (.A(_06344_),
    .X(_06345_));
 sky130_fd_sc_hd__mux2_1 _12157_ (.A0(net2032),
    .A1(_04498_),
    .S(_06345_),
    .X(_06346_));
 sky130_fd_sc_hd__clkbuf_1 _12158_ (.A(_06346_),
    .X(_01201_));
 sky130_fd_sc_hd__mux2_1 _12159_ (.A0(net52),
    .A1(_04505_),
    .S(_06345_),
    .X(_06347_));
 sky130_fd_sc_hd__clkbuf_1 _12160_ (.A(_06347_),
    .X(_01202_));
 sky130_fd_sc_hd__mux2_1 _12161_ (.A0(net285),
    .A1(_04508_),
    .S(_06345_),
    .X(_06348_));
 sky130_fd_sc_hd__clkbuf_1 _12162_ (.A(_06348_),
    .X(_01203_));
 sky130_fd_sc_hd__mux2_1 _12163_ (.A0(net585),
    .A1(_04511_),
    .S(_06345_),
    .X(_06349_));
 sky130_fd_sc_hd__clkbuf_1 _12164_ (.A(_06349_),
    .X(_01204_));
 sky130_fd_sc_hd__mux2_1 _12165_ (.A0(net209),
    .A1(_04514_),
    .S(_06345_),
    .X(_06350_));
 sky130_fd_sc_hd__clkbuf_1 _12166_ (.A(_06350_),
    .X(_01205_));
 sky130_fd_sc_hd__mux2_1 _12167_ (.A0(net62),
    .A1(_04517_),
    .S(_06345_),
    .X(_06351_));
 sky130_fd_sc_hd__clkbuf_1 _12168_ (.A(_06351_),
    .X(_01206_));
 sky130_fd_sc_hd__mux2_1 _12169_ (.A0(net180),
    .A1(_04520_),
    .S(_06345_),
    .X(_06352_));
 sky130_fd_sc_hd__clkbuf_1 _12170_ (.A(_06352_),
    .X(_01207_));
 sky130_fd_sc_hd__mux2_1 _12171_ (.A0(net401),
    .A1(_04523_),
    .S(_06345_),
    .X(_06353_));
 sky130_fd_sc_hd__clkbuf_1 _12172_ (.A(_06353_),
    .X(_01208_));
 sky130_fd_sc_hd__mux2_1 _12173_ (.A0(net252),
    .A1(_04526_),
    .S(_06345_),
    .X(_06354_));
 sky130_fd_sc_hd__clkbuf_1 _12174_ (.A(_06354_),
    .X(_01209_));
 sky130_fd_sc_hd__mux2_1 _12175_ (.A0(net555),
    .A1(_04529_),
    .S(_06345_),
    .X(_06355_));
 sky130_fd_sc_hd__clkbuf_1 _12176_ (.A(_06355_),
    .X(_01210_));
 sky130_fd_sc_hd__mux2_1 _12177_ (.A0(net328),
    .A1(_04532_),
    .S(_06344_),
    .X(_06356_));
 sky130_fd_sc_hd__clkbuf_1 _12178_ (.A(_06356_),
    .X(_01211_));
 sky130_fd_sc_hd__mux2_1 _12179_ (.A0(net199),
    .A1(_04535_),
    .S(_06344_),
    .X(_06357_));
 sky130_fd_sc_hd__clkbuf_1 _12180_ (.A(_06357_),
    .X(_01212_));
 sky130_fd_sc_hd__mux2_1 _12181_ (.A0(net249),
    .A1(_04538_),
    .S(_06344_),
    .X(_06358_));
 sky130_fd_sc_hd__clkbuf_1 _12182_ (.A(_06358_),
    .X(_01213_));
 sky130_fd_sc_hd__mux2_1 _12183_ (.A0(net1312),
    .A1(_04541_),
    .S(_06344_),
    .X(_06359_));
 sky130_fd_sc_hd__clkbuf_1 _12184_ (.A(_06359_),
    .X(_01214_));
 sky130_fd_sc_hd__mux2_1 _12185_ (.A0(net914),
    .A1(_04544_),
    .S(_06344_),
    .X(_06360_));
 sky130_fd_sc_hd__clkbuf_1 _12186_ (.A(_06360_),
    .X(_01215_));
 sky130_fd_sc_hd__mux2_1 _12187_ (.A0(net1011),
    .A1(_04547_),
    .S(_06344_),
    .X(_06361_));
 sky130_fd_sc_hd__clkbuf_1 _12188_ (.A(_06361_),
    .X(_01216_));
 sky130_fd_sc_hd__nand2b_4 _12189_ (.A_N(_04286_),
    .B(_04408_),
    .Y(_06362_));
 sky130_fd_sc_hd__buf_4 _12190_ (.A(_06362_),
    .X(_06363_));
 sky130_fd_sc_hd__mux2_1 _12191_ (.A0(_06309_),
    .A1(net1984),
    .S(_06363_),
    .X(_06364_));
 sky130_fd_sc_hd__clkbuf_1 _12192_ (.A(_06364_),
    .X(_01217_));
 sky130_fd_sc_hd__mux2_1 _12193_ (.A0(_06314_),
    .A1(net1251),
    .S(_06363_),
    .X(_06365_));
 sky130_fd_sc_hd__clkbuf_1 _12194_ (.A(_06365_),
    .X(_01218_));
 sky130_fd_sc_hd__mux2_1 _12195_ (.A0(_06316_),
    .A1(net584),
    .S(_06363_),
    .X(_06366_));
 sky130_fd_sc_hd__clkbuf_1 _12196_ (.A(_06366_),
    .X(_01219_));
 sky130_fd_sc_hd__mux2_1 _12197_ (.A0(_06318_),
    .A1(net768),
    .S(_06363_),
    .X(_06367_));
 sky130_fd_sc_hd__clkbuf_1 _12198_ (.A(_06367_),
    .X(_01220_));
 sky130_fd_sc_hd__mux2_1 _12199_ (.A0(_06320_),
    .A1(net1017),
    .S(_06363_),
    .X(_06368_));
 sky130_fd_sc_hd__clkbuf_1 _12200_ (.A(_06368_),
    .X(_01221_));
 sky130_fd_sc_hd__mux2_1 _12201_ (.A0(_06322_),
    .A1(net1266),
    .S(_06363_),
    .X(_06369_));
 sky130_fd_sc_hd__clkbuf_1 _12202_ (.A(_06369_),
    .X(_01222_));
 sky130_fd_sc_hd__mux2_1 _12203_ (.A0(_06324_),
    .A1(net1698),
    .S(_06363_),
    .X(_06370_));
 sky130_fd_sc_hd__clkbuf_1 _12204_ (.A(_06370_),
    .X(_01223_));
 sky130_fd_sc_hd__mux2_1 _12205_ (.A0(_06326_),
    .A1(net1442),
    .S(_06363_),
    .X(_06371_));
 sky130_fd_sc_hd__clkbuf_1 _12206_ (.A(_06371_),
    .X(_01224_));
 sky130_fd_sc_hd__mux2_1 _12207_ (.A0(_06328_),
    .A1(net511),
    .S(_06363_),
    .X(_06372_));
 sky130_fd_sc_hd__clkbuf_1 _12208_ (.A(_06372_),
    .X(_01225_));
 sky130_fd_sc_hd__mux2_1 _12209_ (.A0(_06330_),
    .A1(net872),
    .S(_06363_),
    .X(_06373_));
 sky130_fd_sc_hd__clkbuf_1 _12210_ (.A(_06373_),
    .X(_01226_));
 sky130_fd_sc_hd__mux2_1 _12211_ (.A0(_06332_),
    .A1(net150),
    .S(_06362_),
    .X(_06374_));
 sky130_fd_sc_hd__clkbuf_1 _12212_ (.A(_06374_),
    .X(_01227_));
 sky130_fd_sc_hd__mux2_1 _12213_ (.A0(_06334_),
    .A1(net1006),
    .S(_06362_),
    .X(_06375_));
 sky130_fd_sc_hd__clkbuf_1 _12214_ (.A(_06375_),
    .X(_01228_));
 sky130_fd_sc_hd__mux2_1 _12215_ (.A0(_06336_),
    .A1(net1020),
    .S(_06362_),
    .X(_06376_));
 sky130_fd_sc_hd__clkbuf_1 _12216_ (.A(_06376_),
    .X(_01229_));
 sky130_fd_sc_hd__mux2_1 _12217_ (.A0(_06338_),
    .A1(net857),
    .S(_06362_),
    .X(_06377_));
 sky130_fd_sc_hd__clkbuf_1 _12218_ (.A(_06377_),
    .X(_01230_));
 sky130_fd_sc_hd__mux2_1 _12219_ (.A0(_06340_),
    .A1(net614),
    .S(_06362_),
    .X(_06378_));
 sky130_fd_sc_hd__clkbuf_1 _12220_ (.A(_06378_),
    .X(_01231_));
 sky130_fd_sc_hd__mux2_1 _12221_ (.A0(_06342_),
    .A1(net1738),
    .S(_06362_),
    .X(_06379_));
 sky130_fd_sc_hd__clkbuf_1 _12222_ (.A(_06379_),
    .X(_01232_));
 sky130_fd_sc_hd__or3_1 _12223_ (.A(_02484_),
    .B(_02644_),
    .C(_04285_),
    .X(_06380_));
 sky130_fd_sc_hd__clkbuf_4 _12224_ (.A(_06380_),
    .X(_06381_));
 sky130_fd_sc_hd__buf_4 _12225_ (.A(_06381_),
    .X(_06382_));
 sky130_fd_sc_hd__mux2_1 _12226_ (.A0(_06309_),
    .A1(net1737),
    .S(_06382_),
    .X(_06383_));
 sky130_fd_sc_hd__clkbuf_1 _12227_ (.A(_06383_),
    .X(_01233_));
 sky130_fd_sc_hd__mux2_1 _12228_ (.A0(_06314_),
    .A1(net898),
    .S(_06382_),
    .X(_06384_));
 sky130_fd_sc_hd__clkbuf_1 _12229_ (.A(_06384_),
    .X(_01234_));
 sky130_fd_sc_hd__mux2_1 _12230_ (.A0(_06316_),
    .A1(net1816),
    .S(_06382_),
    .X(_06385_));
 sky130_fd_sc_hd__clkbuf_1 _12231_ (.A(_06385_),
    .X(_01235_));
 sky130_fd_sc_hd__mux2_1 _12232_ (.A0(_06318_),
    .A1(net922),
    .S(_06382_),
    .X(_06386_));
 sky130_fd_sc_hd__clkbuf_1 _12233_ (.A(_06386_),
    .X(_01236_));
 sky130_fd_sc_hd__mux2_1 _12234_ (.A0(_06320_),
    .A1(net771),
    .S(_06382_),
    .X(_06387_));
 sky130_fd_sc_hd__clkbuf_1 _12235_ (.A(_06387_),
    .X(_01237_));
 sky130_fd_sc_hd__mux2_1 _12236_ (.A0(_06322_),
    .A1(net1701),
    .S(_06382_),
    .X(_06388_));
 sky130_fd_sc_hd__clkbuf_1 _12237_ (.A(_06388_),
    .X(_01238_));
 sky130_fd_sc_hd__mux2_1 _12238_ (.A0(_06324_),
    .A1(net1942),
    .S(_06382_),
    .X(_06389_));
 sky130_fd_sc_hd__clkbuf_1 _12239_ (.A(_06389_),
    .X(_01239_));
 sky130_fd_sc_hd__mux2_1 _12240_ (.A0(_06326_),
    .A1(net1379),
    .S(_06382_),
    .X(_06390_));
 sky130_fd_sc_hd__clkbuf_1 _12241_ (.A(_06390_),
    .X(_01240_));
 sky130_fd_sc_hd__mux2_1 _12242_ (.A0(_06328_),
    .A1(net1680),
    .S(_06382_),
    .X(_06391_));
 sky130_fd_sc_hd__clkbuf_1 _12243_ (.A(_06391_),
    .X(_01241_));
 sky130_fd_sc_hd__mux2_1 _12244_ (.A0(_06330_),
    .A1(net1159),
    .S(_06382_),
    .X(_06392_));
 sky130_fd_sc_hd__clkbuf_1 _12245_ (.A(_06392_),
    .X(_01242_));
 sky130_fd_sc_hd__mux2_1 _12246_ (.A0(_06332_),
    .A1(net1120),
    .S(_06381_),
    .X(_06393_));
 sky130_fd_sc_hd__clkbuf_1 _12247_ (.A(_06393_),
    .X(_01243_));
 sky130_fd_sc_hd__mux2_1 _12248_ (.A0(_06334_),
    .A1(net867),
    .S(_06381_),
    .X(_06394_));
 sky130_fd_sc_hd__clkbuf_1 _12249_ (.A(_06394_),
    .X(_01244_));
 sky130_fd_sc_hd__mux2_1 _12250_ (.A0(_06336_),
    .A1(net751),
    .S(_06381_),
    .X(_06395_));
 sky130_fd_sc_hd__clkbuf_1 _12251_ (.A(_06395_),
    .X(_01245_));
 sky130_fd_sc_hd__mux2_1 _12252_ (.A0(_06338_),
    .A1(net1552),
    .S(_06381_),
    .X(_06396_));
 sky130_fd_sc_hd__clkbuf_1 _12253_ (.A(_06396_),
    .X(_01246_));
 sky130_fd_sc_hd__mux2_1 _12254_ (.A0(_06340_),
    .A1(net1261),
    .S(_06381_),
    .X(_06397_));
 sky130_fd_sc_hd__clkbuf_1 _12255_ (.A(_06397_),
    .X(_01247_));
 sky130_fd_sc_hd__mux2_1 _12256_ (.A0(_06342_),
    .A1(net944),
    .S(_06381_),
    .X(_06398_));
 sky130_fd_sc_hd__clkbuf_1 _12257_ (.A(_06398_),
    .X(_01248_));
 sky130_fd_sc_hd__buf_6 _12258_ (.A(_04325_),
    .X(_06399_));
 sky130_fd_sc_hd__nor2_4 _12259_ (.A(_06399_),
    .B(_04461_),
    .Y(_06400_));
 sky130_fd_sc_hd__buf_4 _12260_ (.A(_06400_),
    .X(_06401_));
 sky130_fd_sc_hd__mux2_1 _12261_ (.A0(net529),
    .A1(_04498_),
    .S(_06401_),
    .X(_06402_));
 sky130_fd_sc_hd__clkbuf_1 _12262_ (.A(_06402_),
    .X(_01249_));
 sky130_fd_sc_hd__mux2_1 _12263_ (.A0(net77),
    .A1(_04505_),
    .S(_06401_),
    .X(_06403_));
 sky130_fd_sc_hd__clkbuf_1 _12264_ (.A(_06403_),
    .X(_01250_));
 sky130_fd_sc_hd__mux2_1 _12265_ (.A0(net380),
    .A1(_04508_),
    .S(_06401_),
    .X(_06404_));
 sky130_fd_sc_hd__clkbuf_1 _12266_ (.A(_06404_),
    .X(_01251_));
 sky130_fd_sc_hd__mux2_1 _12267_ (.A0(net147),
    .A1(_04511_),
    .S(_06401_),
    .X(_06405_));
 sky130_fd_sc_hd__clkbuf_1 _12268_ (.A(_06405_),
    .X(_01252_));
 sky130_fd_sc_hd__mux2_1 _12269_ (.A0(net169),
    .A1(_04514_),
    .S(_06401_),
    .X(_02064_));
 sky130_fd_sc_hd__clkbuf_1 _12270_ (.A(_02064_),
    .X(_01253_));
 sky130_fd_sc_hd__mux2_1 _12271_ (.A0(net80),
    .A1(_04517_),
    .S(_06401_),
    .X(_02065_));
 sky130_fd_sc_hd__clkbuf_1 _12272_ (.A(_02065_),
    .X(_01254_));
 sky130_fd_sc_hd__mux2_1 _12273_ (.A0(net81),
    .A1(_04520_),
    .S(_06401_),
    .X(_02066_));
 sky130_fd_sc_hd__clkbuf_1 _12274_ (.A(_02066_),
    .X(_01255_));
 sky130_fd_sc_hd__mux2_1 _12275_ (.A0(net430),
    .A1(_04523_),
    .S(_06401_),
    .X(_02067_));
 sky130_fd_sc_hd__clkbuf_1 _12276_ (.A(_02067_),
    .X(_01256_));
 sky130_fd_sc_hd__mux2_1 _12277_ (.A0(net297),
    .A1(_04526_),
    .S(_06401_),
    .X(_02068_));
 sky130_fd_sc_hd__clkbuf_1 _12278_ (.A(_02068_),
    .X(_01257_));
 sky130_fd_sc_hd__mux2_1 _12279_ (.A0(net255),
    .A1(_04529_),
    .S(_06401_),
    .X(_02069_));
 sky130_fd_sc_hd__clkbuf_1 _12280_ (.A(_02069_),
    .X(_01258_));
 sky130_fd_sc_hd__mux2_1 _12281_ (.A0(net98),
    .A1(_04532_),
    .S(_06400_),
    .X(_02070_));
 sky130_fd_sc_hd__clkbuf_1 _12282_ (.A(_02070_),
    .X(_01259_));
 sky130_fd_sc_hd__mux2_1 _12283_ (.A0(net635),
    .A1(_04535_),
    .S(_06400_),
    .X(_02071_));
 sky130_fd_sc_hd__clkbuf_1 _12284_ (.A(_02071_),
    .X(_01260_));
 sky130_fd_sc_hd__mux2_1 _12285_ (.A0(net669),
    .A1(_04538_),
    .S(_06400_),
    .X(_02072_));
 sky130_fd_sc_hd__clkbuf_1 _12286_ (.A(_02072_),
    .X(_01261_));
 sky130_fd_sc_hd__mux2_1 _12287_ (.A0(net623),
    .A1(_04541_),
    .S(_06400_),
    .X(_02073_));
 sky130_fd_sc_hd__clkbuf_1 _12288_ (.A(_02073_),
    .X(_01262_));
 sky130_fd_sc_hd__mux2_1 _12289_ (.A0(net473),
    .A1(_04544_),
    .S(_06400_),
    .X(_02074_));
 sky130_fd_sc_hd__clkbuf_1 _12290_ (.A(_02074_),
    .X(_01263_));
 sky130_fd_sc_hd__mux2_1 _12291_ (.A0(net499),
    .A1(_04547_),
    .S(_06400_),
    .X(_02075_));
 sky130_fd_sc_hd__clkbuf_1 _12292_ (.A(_02075_),
    .X(_01264_));
 sky130_fd_sc_hd__nor2_8 _12293_ (.A(_04072_),
    .B(_06399_),
    .Y(_02076_));
 sky130_fd_sc_hd__buf_4 _12294_ (.A(_02076_),
    .X(_02077_));
 sky130_fd_sc_hd__mux2_1 _12295_ (.A0(net408),
    .A1(_04498_),
    .S(_02077_),
    .X(_02078_));
 sky130_fd_sc_hd__clkbuf_1 _12296_ (.A(_02078_),
    .X(_01265_));
 sky130_fd_sc_hd__mux2_1 _12297_ (.A0(net76),
    .A1(_04505_),
    .S(_02077_),
    .X(_02079_));
 sky130_fd_sc_hd__clkbuf_1 _12298_ (.A(_02079_),
    .X(_01266_));
 sky130_fd_sc_hd__mux2_1 _12299_ (.A0(net141),
    .A1(_04508_),
    .S(_02077_),
    .X(_02080_));
 sky130_fd_sc_hd__clkbuf_1 _12300_ (.A(_02080_),
    .X(_01267_));
 sky130_fd_sc_hd__mux2_1 _12301_ (.A0(net360),
    .A1(_04511_),
    .S(_02077_),
    .X(_02081_));
 sky130_fd_sc_hd__clkbuf_1 _12302_ (.A(_02081_),
    .X(_01268_));
 sky130_fd_sc_hd__mux2_1 _12303_ (.A0(net237),
    .A1(_04514_),
    .S(_02077_),
    .X(_02082_));
 sky130_fd_sc_hd__clkbuf_1 _12304_ (.A(_02082_),
    .X(_01269_));
 sky130_fd_sc_hd__mux2_1 _12305_ (.A0(net540),
    .A1(_04517_),
    .S(_02077_),
    .X(_02083_));
 sky130_fd_sc_hd__clkbuf_1 _12306_ (.A(_02083_),
    .X(_01270_));
 sky130_fd_sc_hd__mux2_1 _12307_ (.A0(net315),
    .A1(_04520_),
    .S(_02077_),
    .X(_02084_));
 sky130_fd_sc_hd__clkbuf_1 _12308_ (.A(_02084_),
    .X(_01271_));
 sky130_fd_sc_hd__mux2_1 _12309_ (.A0(net173),
    .A1(_04523_),
    .S(_02077_),
    .X(_02085_));
 sky130_fd_sc_hd__clkbuf_1 _12310_ (.A(_02085_),
    .X(_01272_));
 sky130_fd_sc_hd__mux2_1 _12311_ (.A0(net656),
    .A1(_04526_),
    .S(_02077_),
    .X(_02086_));
 sky130_fd_sc_hd__clkbuf_1 _12312_ (.A(_02086_),
    .X(_01273_));
 sky130_fd_sc_hd__mux2_1 _12313_ (.A0(net215),
    .A1(_04529_),
    .S(_02077_),
    .X(_02087_));
 sky130_fd_sc_hd__clkbuf_1 _12314_ (.A(_02087_),
    .X(_01274_));
 sky130_fd_sc_hd__mux2_1 _12315_ (.A0(net111),
    .A1(_04532_),
    .S(_02076_),
    .X(_02088_));
 sky130_fd_sc_hd__clkbuf_1 _12316_ (.A(_02088_),
    .X(_01275_));
 sky130_fd_sc_hd__mux2_1 _12317_ (.A0(net420),
    .A1(_04535_),
    .S(_02076_),
    .X(_02089_));
 sky130_fd_sc_hd__clkbuf_1 _12318_ (.A(_02089_),
    .X(_01276_));
 sky130_fd_sc_hd__mux2_1 _12319_ (.A0(net295),
    .A1(_04538_),
    .S(_02076_),
    .X(_02090_));
 sky130_fd_sc_hd__clkbuf_1 _12320_ (.A(_02090_),
    .X(_01277_));
 sky130_fd_sc_hd__mux2_1 _12321_ (.A0(net414),
    .A1(_04541_),
    .S(_02076_),
    .X(_02091_));
 sky130_fd_sc_hd__clkbuf_1 _12322_ (.A(_02091_),
    .X(_01278_));
 sky130_fd_sc_hd__mux2_1 _12323_ (.A0(net368),
    .A1(_04544_),
    .S(_02076_),
    .X(_02092_));
 sky130_fd_sc_hd__clkbuf_1 _12324_ (.A(_02092_),
    .X(_01279_));
 sky130_fd_sc_hd__mux2_1 _12325_ (.A0(net448),
    .A1(_04547_),
    .S(_02076_),
    .X(_02093_));
 sky130_fd_sc_hd__clkbuf_1 _12326_ (.A(_02093_),
    .X(_01280_));
 sky130_fd_sc_hd__nor2_4 _12327_ (.A(_06399_),
    .B(_04501_),
    .Y(_02094_));
 sky130_fd_sc_hd__buf_4 _12328_ (.A(_02094_),
    .X(_02095_));
 sky130_fd_sc_hd__mux2_1 _12329_ (.A0(net365),
    .A1(_04498_),
    .S(_02095_),
    .X(_02096_));
 sky130_fd_sc_hd__clkbuf_1 _12330_ (.A(_02096_),
    .X(_01281_));
 sky130_fd_sc_hd__mux2_1 _12331_ (.A0(net674),
    .A1(_04505_),
    .S(_02095_),
    .X(_02097_));
 sky130_fd_sc_hd__clkbuf_1 _12332_ (.A(_02097_),
    .X(_01282_));
 sky130_fd_sc_hd__mux2_1 _12333_ (.A0(net286),
    .A1(_04508_),
    .S(_02095_),
    .X(_02098_));
 sky130_fd_sc_hd__clkbuf_1 _12334_ (.A(_02098_),
    .X(_01283_));
 sky130_fd_sc_hd__mux2_1 _12335_ (.A0(net480),
    .A1(_04511_),
    .S(_02095_),
    .X(_02099_));
 sky130_fd_sc_hd__clkbuf_1 _12336_ (.A(_02099_),
    .X(_01284_));
 sky130_fd_sc_hd__mux2_1 _12337_ (.A0(net329),
    .A1(_04514_),
    .S(_02095_),
    .X(_02100_));
 sky130_fd_sc_hd__clkbuf_1 _12338_ (.A(_02100_),
    .X(_01285_));
 sky130_fd_sc_hd__mux2_1 _12339_ (.A0(net735),
    .A1(_04517_),
    .S(_02095_),
    .X(_02101_));
 sky130_fd_sc_hd__clkbuf_1 _12340_ (.A(_02101_),
    .X(_01286_));
 sky130_fd_sc_hd__mux2_1 _12341_ (.A0(net602),
    .A1(_04520_),
    .S(_02095_),
    .X(_02102_));
 sky130_fd_sc_hd__clkbuf_1 _12342_ (.A(_02102_),
    .X(_01287_));
 sky130_fd_sc_hd__mux2_1 _12343_ (.A0(net240),
    .A1(_04523_),
    .S(_02095_),
    .X(_02103_));
 sky130_fd_sc_hd__clkbuf_1 _12344_ (.A(_02103_),
    .X(_01288_));
 sky130_fd_sc_hd__mux2_1 _12345_ (.A0(net264),
    .A1(_04526_),
    .S(_02095_),
    .X(_02104_));
 sky130_fd_sc_hd__clkbuf_1 _12346_ (.A(_02104_),
    .X(_01289_));
 sky130_fd_sc_hd__mux2_1 _12347_ (.A0(net308),
    .A1(_04529_),
    .S(_02095_),
    .X(_02105_));
 sky130_fd_sc_hd__clkbuf_1 _12348_ (.A(_02105_),
    .X(_01290_));
 sky130_fd_sc_hd__mux2_1 _12349_ (.A0(net601),
    .A1(_04532_),
    .S(_02094_),
    .X(_02106_));
 sky130_fd_sc_hd__clkbuf_1 _12350_ (.A(_02106_),
    .X(_01291_));
 sky130_fd_sc_hd__mux2_1 _12351_ (.A0(net413),
    .A1(_04535_),
    .S(_02094_),
    .X(_02107_));
 sky130_fd_sc_hd__clkbuf_1 _12352_ (.A(_02107_),
    .X(_01292_));
 sky130_fd_sc_hd__mux2_1 _12353_ (.A0(net145),
    .A1(_04538_),
    .S(_02094_),
    .X(_02108_));
 sky130_fd_sc_hd__clkbuf_1 _12354_ (.A(_02108_),
    .X(_01293_));
 sky130_fd_sc_hd__mux2_1 _12355_ (.A0(net90),
    .A1(_04541_),
    .S(_02094_),
    .X(_02109_));
 sky130_fd_sc_hd__clkbuf_1 _12356_ (.A(_02109_),
    .X(_01294_));
 sky130_fd_sc_hd__mux2_1 _12357_ (.A0(net203),
    .A1(_04544_),
    .S(_02094_),
    .X(_02110_));
 sky130_fd_sc_hd__clkbuf_1 _12358_ (.A(_02110_),
    .X(_01295_));
 sky130_fd_sc_hd__mux2_1 _12359_ (.A0(net201),
    .A1(_04547_),
    .S(_02094_),
    .X(_02111_));
 sky130_fd_sc_hd__clkbuf_1 _12360_ (.A(_02111_),
    .X(_01296_));
 sky130_fd_sc_hd__or2_1 _12361_ (.A(_04225_),
    .B(_06399_),
    .X(_02112_));
 sky130_fd_sc_hd__buf_4 _12362_ (.A(_02112_),
    .X(_02113_));
 sky130_fd_sc_hd__buf_4 _12363_ (.A(_02113_),
    .X(_02114_));
 sky130_fd_sc_hd__mux2_1 _12364_ (.A0(_06309_),
    .A1(net836),
    .S(_02114_),
    .X(_02115_));
 sky130_fd_sc_hd__clkbuf_1 _12365_ (.A(_02115_),
    .X(_01297_));
 sky130_fd_sc_hd__mux2_1 _12366_ (.A0(_06314_),
    .A1(net502),
    .S(_02114_),
    .X(_02116_));
 sky130_fd_sc_hd__clkbuf_1 _12367_ (.A(_02116_),
    .X(_01298_));
 sky130_fd_sc_hd__mux2_1 _12368_ (.A0(_06316_),
    .A1(net958),
    .S(_02114_),
    .X(_02117_));
 sky130_fd_sc_hd__clkbuf_1 _12369_ (.A(_02117_),
    .X(_01299_));
 sky130_fd_sc_hd__mux2_1 _12370_ (.A0(_06318_),
    .A1(net970),
    .S(_02114_),
    .X(_02118_));
 sky130_fd_sc_hd__clkbuf_1 _12371_ (.A(_02118_),
    .X(_01300_));
 sky130_fd_sc_hd__mux2_1 _12372_ (.A0(_06320_),
    .A1(net1999),
    .S(_02114_),
    .X(_02119_));
 sky130_fd_sc_hd__clkbuf_1 _12373_ (.A(_02119_),
    .X(_01301_));
 sky130_fd_sc_hd__mux2_1 _12374_ (.A0(_06322_),
    .A1(net186),
    .S(_02114_),
    .X(_02120_));
 sky130_fd_sc_hd__clkbuf_1 _12375_ (.A(_02120_),
    .X(_01302_));
 sky130_fd_sc_hd__mux2_1 _12376_ (.A0(_06324_),
    .A1(net686),
    .S(_02114_),
    .X(_02121_));
 sky130_fd_sc_hd__clkbuf_1 _12377_ (.A(_02121_),
    .X(_01303_));
 sky130_fd_sc_hd__mux2_1 _12378_ (.A0(_06326_),
    .A1(net1075),
    .S(_02114_),
    .X(_02122_));
 sky130_fd_sc_hd__clkbuf_1 _12379_ (.A(_02122_),
    .X(_01304_));
 sky130_fd_sc_hd__mux2_1 _12380_ (.A0(_06328_),
    .A1(net1037),
    .S(_02114_),
    .X(_02123_));
 sky130_fd_sc_hd__clkbuf_1 _12381_ (.A(_02123_),
    .X(_01305_));
 sky130_fd_sc_hd__mux2_1 _12382_ (.A0(_06330_),
    .A1(net1643),
    .S(_02114_),
    .X(_02124_));
 sky130_fd_sc_hd__clkbuf_1 _12383_ (.A(_02124_),
    .X(_01306_));
 sky130_fd_sc_hd__mux2_1 _12384_ (.A0(_06332_),
    .A1(net792),
    .S(_02113_),
    .X(_02125_));
 sky130_fd_sc_hd__clkbuf_1 _12385_ (.A(_02125_),
    .X(_01307_));
 sky130_fd_sc_hd__mux2_1 _12386_ (.A0(_06334_),
    .A1(net620),
    .S(_02113_),
    .X(_02126_));
 sky130_fd_sc_hd__clkbuf_1 _12387_ (.A(_02126_),
    .X(_01308_));
 sky130_fd_sc_hd__mux2_1 _12388_ (.A0(_06336_),
    .A1(net1333),
    .S(_02113_),
    .X(_02127_));
 sky130_fd_sc_hd__clkbuf_1 _12389_ (.A(_02127_),
    .X(_01309_));
 sky130_fd_sc_hd__mux2_1 _12390_ (.A0(_06338_),
    .A1(net951),
    .S(_02113_),
    .X(_02128_));
 sky130_fd_sc_hd__clkbuf_1 _12391_ (.A(_02128_),
    .X(_01310_));
 sky130_fd_sc_hd__mux2_1 _12392_ (.A0(_06340_),
    .A1(net729),
    .S(_02113_),
    .X(_02129_));
 sky130_fd_sc_hd__clkbuf_1 _12393_ (.A(_02129_),
    .X(_01311_));
 sky130_fd_sc_hd__mux2_1 _12394_ (.A0(_06342_),
    .A1(net1592),
    .S(_02113_),
    .X(_02130_));
 sky130_fd_sc_hd__clkbuf_1 _12395_ (.A(_02130_),
    .X(_01312_));
 sky130_fd_sc_hd__nor2_4 _12396_ (.A(_06399_),
    .B(_04569_),
    .Y(_02131_));
 sky130_fd_sc_hd__buf_4 _12397_ (.A(_02131_),
    .X(_02132_));
 sky130_fd_sc_hd__mux2_1 _12398_ (.A0(net321),
    .A1(_04498_),
    .S(_02132_),
    .X(_02133_));
 sky130_fd_sc_hd__clkbuf_1 _12399_ (.A(_02133_),
    .X(_01313_));
 sky130_fd_sc_hd__mux2_1 _12400_ (.A0(net516),
    .A1(_04505_),
    .S(_02132_),
    .X(_02134_));
 sky130_fd_sc_hd__clkbuf_1 _12401_ (.A(_02134_),
    .X(_01314_));
 sky130_fd_sc_hd__mux2_1 _12402_ (.A0(net825),
    .A1(_04508_),
    .S(_02132_),
    .X(_02135_));
 sky130_fd_sc_hd__clkbuf_1 _12403_ (.A(_02135_),
    .X(_01315_));
 sky130_fd_sc_hd__mux2_1 _12404_ (.A0(net509),
    .A1(_04511_),
    .S(_02132_),
    .X(_02136_));
 sky130_fd_sc_hd__clkbuf_1 _12405_ (.A(_02136_),
    .X(_01316_));
 sky130_fd_sc_hd__mux2_1 _12406_ (.A0(net631),
    .A1(_04514_),
    .S(_02132_),
    .X(_02137_));
 sky130_fd_sc_hd__clkbuf_1 _12407_ (.A(_02137_),
    .X(_01317_));
 sky130_fd_sc_hd__mux2_1 _12408_ (.A0(net558),
    .A1(_04517_),
    .S(_02132_),
    .X(_02138_));
 sky130_fd_sc_hd__clkbuf_1 _12409_ (.A(_02138_),
    .X(_01318_));
 sky130_fd_sc_hd__mux2_1 _12410_ (.A0(net95),
    .A1(_04520_),
    .S(_02132_),
    .X(_02139_));
 sky130_fd_sc_hd__clkbuf_1 _12411_ (.A(_02139_),
    .X(_01319_));
 sky130_fd_sc_hd__mux2_1 _12412_ (.A0(net192),
    .A1(_04523_),
    .S(_02132_),
    .X(_02140_));
 sky130_fd_sc_hd__clkbuf_1 _12413_ (.A(_02140_),
    .X(_01320_));
 sky130_fd_sc_hd__mux2_1 _12414_ (.A0(net1158),
    .A1(_04526_),
    .S(_02132_),
    .X(_02141_));
 sky130_fd_sc_hd__clkbuf_1 _12415_ (.A(_02141_),
    .X(_01321_));
 sky130_fd_sc_hd__mux2_1 _12416_ (.A0(net573),
    .A1(_04529_),
    .S(_02132_),
    .X(_02142_));
 sky130_fd_sc_hd__clkbuf_1 _12417_ (.A(_02142_),
    .X(_01322_));
 sky130_fd_sc_hd__mux2_1 _12418_ (.A0(net947),
    .A1(_04532_),
    .S(_02131_),
    .X(_02143_));
 sky130_fd_sc_hd__clkbuf_1 _12419_ (.A(_02143_),
    .X(_01323_));
 sky130_fd_sc_hd__mux2_1 _12420_ (.A0(net716),
    .A1(_04535_),
    .S(_02131_),
    .X(_02144_));
 sky130_fd_sc_hd__clkbuf_1 _12421_ (.A(_02144_),
    .X(_01324_));
 sky130_fd_sc_hd__mux2_1 _12422_ (.A0(net426),
    .A1(_04538_),
    .S(_02131_),
    .X(_02145_));
 sky130_fd_sc_hd__clkbuf_1 _12423_ (.A(_02145_),
    .X(_01325_));
 sky130_fd_sc_hd__mux2_1 _12424_ (.A0(net526),
    .A1(_04541_),
    .S(_02131_),
    .X(_02146_));
 sky130_fd_sc_hd__clkbuf_1 _12425_ (.A(_02146_),
    .X(_01326_));
 sky130_fd_sc_hd__mux2_1 _12426_ (.A0(net159),
    .A1(_04544_),
    .S(_02131_),
    .X(_02147_));
 sky130_fd_sc_hd__clkbuf_1 _12427_ (.A(_02147_),
    .X(_01327_));
 sky130_fd_sc_hd__mux2_1 _12428_ (.A0(net528),
    .A1(_04547_),
    .S(_02131_),
    .X(_02148_));
 sky130_fd_sc_hd__clkbuf_1 _12429_ (.A(_02148_),
    .X(_01328_));
 sky130_fd_sc_hd__or2_1 _12430_ (.A(_04184_),
    .B(_04325_),
    .X(_02149_));
 sky130_fd_sc_hd__clkbuf_4 _12431_ (.A(_02149_),
    .X(_02150_));
 sky130_fd_sc_hd__buf_4 _12432_ (.A(_02150_),
    .X(_02151_));
 sky130_fd_sc_hd__mux2_1 _12433_ (.A0(_06309_),
    .A1(net592),
    .S(_02151_),
    .X(_02152_));
 sky130_fd_sc_hd__clkbuf_1 _12434_ (.A(_02152_),
    .X(_01329_));
 sky130_fd_sc_hd__mux2_1 _12435_ (.A0(_06314_),
    .A1(net1237),
    .S(_02151_),
    .X(_02153_));
 sky130_fd_sc_hd__clkbuf_1 _12436_ (.A(_02153_),
    .X(_01330_));
 sky130_fd_sc_hd__mux2_1 _12437_ (.A0(_06316_),
    .A1(net675),
    .S(_02151_),
    .X(_02154_));
 sky130_fd_sc_hd__clkbuf_1 _12438_ (.A(_02154_),
    .X(_01331_));
 sky130_fd_sc_hd__mux2_1 _12439_ (.A0(_06318_),
    .A1(net506),
    .S(_02151_),
    .X(_02155_));
 sky130_fd_sc_hd__clkbuf_1 _12440_ (.A(_02155_),
    .X(_01332_));
 sky130_fd_sc_hd__mux2_1 _12441_ (.A0(_06320_),
    .A1(net1145),
    .S(_02151_),
    .X(_02156_));
 sky130_fd_sc_hd__clkbuf_1 _12442_ (.A(_02156_),
    .X(_01333_));
 sky130_fd_sc_hd__mux2_1 _12443_ (.A0(_06322_),
    .A1(net1528),
    .S(_02151_),
    .X(_02157_));
 sky130_fd_sc_hd__clkbuf_1 _12444_ (.A(_02157_),
    .X(_01334_));
 sky130_fd_sc_hd__mux2_1 _12445_ (.A0(_06324_),
    .A1(net1118),
    .S(_02151_),
    .X(_02158_));
 sky130_fd_sc_hd__clkbuf_1 _12446_ (.A(_02158_),
    .X(_01335_));
 sky130_fd_sc_hd__mux2_1 _12447_ (.A0(_06326_),
    .A1(net1523),
    .S(_02151_),
    .X(_02159_));
 sky130_fd_sc_hd__clkbuf_1 _12448_ (.A(_02159_),
    .X(_01336_));
 sky130_fd_sc_hd__mux2_1 _12449_ (.A0(_06328_),
    .A1(net1413),
    .S(_02151_),
    .X(_02160_));
 sky130_fd_sc_hd__clkbuf_1 _12450_ (.A(_02160_),
    .X(_01337_));
 sky130_fd_sc_hd__mux2_1 _12451_ (.A0(_06330_),
    .A1(net966),
    .S(_02151_),
    .X(_02161_));
 sky130_fd_sc_hd__clkbuf_1 _12452_ (.A(_02161_),
    .X(_01338_));
 sky130_fd_sc_hd__mux2_1 _12453_ (.A0(_06332_),
    .A1(net1341),
    .S(_02150_),
    .X(_02162_));
 sky130_fd_sc_hd__clkbuf_1 _12454_ (.A(_02162_),
    .X(_01339_));
 sky130_fd_sc_hd__mux2_1 _12455_ (.A0(_06334_),
    .A1(net1018),
    .S(_02150_),
    .X(_02163_));
 sky130_fd_sc_hd__clkbuf_1 _12456_ (.A(_02163_),
    .X(_01340_));
 sky130_fd_sc_hd__mux2_1 _12457_ (.A0(_06336_),
    .A1(net253),
    .S(_02150_),
    .X(_02164_));
 sky130_fd_sc_hd__clkbuf_1 _12458_ (.A(_02164_),
    .X(_01341_));
 sky130_fd_sc_hd__mux2_1 _12459_ (.A0(_06338_),
    .A1(net1426),
    .S(_02150_),
    .X(_02165_));
 sky130_fd_sc_hd__clkbuf_1 _12460_ (.A(_02165_),
    .X(_01342_));
 sky130_fd_sc_hd__mux2_1 _12461_ (.A0(_06340_),
    .A1(net2009),
    .S(_02150_),
    .X(_02166_));
 sky130_fd_sc_hd__clkbuf_1 _12462_ (.A(_02166_),
    .X(_01343_));
 sky130_fd_sc_hd__mux2_1 _12463_ (.A0(_06342_),
    .A1(net683),
    .S(_02150_),
    .X(_02167_));
 sky130_fd_sc_hd__clkbuf_1 _12464_ (.A(_02167_),
    .X(_01344_));
 sky130_fd_sc_hd__or2_1 _12465_ (.A(_06399_),
    .B(_04607_),
    .X(_02168_));
 sky130_fd_sc_hd__buf_4 _12466_ (.A(_02168_),
    .X(_02169_));
 sky130_fd_sc_hd__buf_4 _12467_ (.A(_02169_),
    .X(_02170_));
 sky130_fd_sc_hd__mux2_1 _12468_ (.A0(_06309_),
    .A1(net1132),
    .S(_02170_),
    .X(_02171_));
 sky130_fd_sc_hd__clkbuf_1 _12469_ (.A(_02171_),
    .X(_01345_));
 sky130_fd_sc_hd__mux2_1 _12470_ (.A0(_06314_),
    .A1(net1048),
    .S(_02170_),
    .X(_02172_));
 sky130_fd_sc_hd__clkbuf_1 _12471_ (.A(_02172_),
    .X(_01346_));
 sky130_fd_sc_hd__mux2_1 _12472_ (.A0(_06316_),
    .A1(net1008),
    .S(_02170_),
    .X(_02173_));
 sky130_fd_sc_hd__clkbuf_1 _12473_ (.A(_02173_),
    .X(_01347_));
 sky130_fd_sc_hd__mux2_1 _12474_ (.A0(_06318_),
    .A1(net340),
    .S(_02170_),
    .X(_02174_));
 sky130_fd_sc_hd__clkbuf_1 _12475_ (.A(_02174_),
    .X(_01348_));
 sky130_fd_sc_hd__mux2_1 _12476_ (.A0(_06320_),
    .A1(net1414),
    .S(_02170_),
    .X(_02175_));
 sky130_fd_sc_hd__clkbuf_1 _12477_ (.A(_02175_),
    .X(_01349_));
 sky130_fd_sc_hd__mux2_1 _12478_ (.A0(_06322_),
    .A1(net1865),
    .S(_02170_),
    .X(_02176_));
 sky130_fd_sc_hd__clkbuf_1 _12479_ (.A(_02176_),
    .X(_01350_));
 sky130_fd_sc_hd__mux2_1 _12480_ (.A0(_06324_),
    .A1(net1065),
    .S(_02170_),
    .X(_02177_));
 sky130_fd_sc_hd__clkbuf_1 _12481_ (.A(_02177_),
    .X(_01351_));
 sky130_fd_sc_hd__mux2_1 _12482_ (.A0(_06326_),
    .A1(net818),
    .S(_02170_),
    .X(_02178_));
 sky130_fd_sc_hd__clkbuf_1 _12483_ (.A(_02178_),
    .X(_01352_));
 sky130_fd_sc_hd__mux2_1 _12484_ (.A0(_06328_),
    .A1(net851),
    .S(_02170_),
    .X(_02179_));
 sky130_fd_sc_hd__clkbuf_1 _12485_ (.A(_02179_),
    .X(_01353_));
 sky130_fd_sc_hd__mux2_1 _12486_ (.A0(_06330_),
    .A1(net1204),
    .S(_02170_),
    .X(_02180_));
 sky130_fd_sc_hd__clkbuf_1 _12487_ (.A(_02180_),
    .X(_01354_));
 sky130_fd_sc_hd__mux2_1 _12488_ (.A0(_06332_),
    .A1(net1381),
    .S(_02169_),
    .X(_02181_));
 sky130_fd_sc_hd__clkbuf_1 _12489_ (.A(_02181_),
    .X(_01355_));
 sky130_fd_sc_hd__mux2_1 _12490_ (.A0(_06334_),
    .A1(net1395),
    .S(_02169_),
    .X(_02182_));
 sky130_fd_sc_hd__clkbuf_1 _12491_ (.A(_02182_),
    .X(_01356_));
 sky130_fd_sc_hd__mux2_1 _12492_ (.A0(_06336_),
    .A1(net718),
    .S(_02169_),
    .X(_02183_));
 sky130_fd_sc_hd__clkbuf_1 _12493_ (.A(_02183_),
    .X(_01357_));
 sky130_fd_sc_hd__mux2_1 _12494_ (.A0(_06338_),
    .A1(net728),
    .S(_02169_),
    .X(_02184_));
 sky130_fd_sc_hd__clkbuf_1 _12495_ (.A(_02184_),
    .X(_01358_));
 sky130_fd_sc_hd__mux2_1 _12496_ (.A0(_06340_),
    .A1(net1788),
    .S(_02169_),
    .X(_02185_));
 sky130_fd_sc_hd__clkbuf_1 _12497_ (.A(_02185_),
    .X(_01359_));
 sky130_fd_sc_hd__mux2_1 _12498_ (.A0(_06342_),
    .A1(net1253),
    .S(_02169_),
    .X(_02186_));
 sky130_fd_sc_hd__clkbuf_1 _12499_ (.A(_02186_),
    .X(_01360_));
 sky130_fd_sc_hd__or3_1 _12500_ (.A(_02506_),
    .B(_02644_),
    .C(_04367_),
    .X(_02187_));
 sky130_fd_sc_hd__clkbuf_4 _12501_ (.A(_02187_),
    .X(_02188_));
 sky130_fd_sc_hd__buf_4 _12502_ (.A(_02188_),
    .X(_02189_));
 sky130_fd_sc_hd__mux2_1 _12503_ (.A0(_06309_),
    .A1(net2021),
    .S(_02189_),
    .X(_02190_));
 sky130_fd_sc_hd__clkbuf_1 _12504_ (.A(_02190_),
    .X(_01361_));
 sky130_fd_sc_hd__mux2_1 _12505_ (.A0(_06314_),
    .A1(net766),
    .S(_02189_),
    .X(_02191_));
 sky130_fd_sc_hd__clkbuf_1 _12506_ (.A(_02191_),
    .X(_01362_));
 sky130_fd_sc_hd__mux2_1 _12507_ (.A0(_06316_),
    .A1(net2056),
    .S(_02189_),
    .X(_02192_));
 sky130_fd_sc_hd__clkbuf_1 _12508_ (.A(_02192_),
    .X(_01363_));
 sky130_fd_sc_hd__mux2_1 _12509_ (.A0(_06318_),
    .A1(net2012),
    .S(_02189_),
    .X(_02193_));
 sky130_fd_sc_hd__clkbuf_1 _12510_ (.A(_02193_),
    .X(_01364_));
 sky130_fd_sc_hd__mux2_1 _12511_ (.A0(_06320_),
    .A1(net2027),
    .S(_02189_),
    .X(_02194_));
 sky130_fd_sc_hd__clkbuf_1 _12512_ (.A(_02194_),
    .X(_01365_));
 sky130_fd_sc_hd__mux2_1 _12513_ (.A0(_06322_),
    .A1(net1723),
    .S(_02189_),
    .X(_02195_));
 sky130_fd_sc_hd__clkbuf_1 _12514_ (.A(_02195_),
    .X(_01366_));
 sky130_fd_sc_hd__mux2_1 _12515_ (.A0(_06324_),
    .A1(net1949),
    .S(_02189_),
    .X(_02196_));
 sky130_fd_sc_hd__clkbuf_1 _12516_ (.A(_02196_),
    .X(_01367_));
 sky130_fd_sc_hd__mux2_1 _12517_ (.A0(_06326_),
    .A1(net2024),
    .S(_02189_),
    .X(_02197_));
 sky130_fd_sc_hd__clkbuf_1 _12518_ (.A(_02197_),
    .X(_01368_));
 sky130_fd_sc_hd__mux2_1 _12519_ (.A0(_06328_),
    .A1(net1526),
    .S(_02189_),
    .X(_02198_));
 sky130_fd_sc_hd__clkbuf_1 _12520_ (.A(_02198_),
    .X(_01369_));
 sky130_fd_sc_hd__mux2_1 _12521_ (.A0(_06330_),
    .A1(net1218),
    .S(_02189_),
    .X(_02199_));
 sky130_fd_sc_hd__clkbuf_1 _12522_ (.A(_02199_),
    .X(_01370_));
 sky130_fd_sc_hd__mux2_1 _12523_ (.A0(_06332_),
    .A1(net1751),
    .S(_02188_),
    .X(_02200_));
 sky130_fd_sc_hd__clkbuf_1 _12524_ (.A(_02200_),
    .X(_01371_));
 sky130_fd_sc_hd__mux2_1 _12525_ (.A0(_06334_),
    .A1(net1519),
    .S(_02188_),
    .X(_02201_));
 sky130_fd_sc_hd__clkbuf_1 _12526_ (.A(_02201_),
    .X(_01372_));
 sky130_fd_sc_hd__mux2_1 _12527_ (.A0(_06336_),
    .A1(net1818),
    .S(_02188_),
    .X(_02202_));
 sky130_fd_sc_hd__clkbuf_1 _12528_ (.A(_02202_),
    .X(_01373_));
 sky130_fd_sc_hd__mux2_1 _12529_ (.A0(_06338_),
    .A1(net1967),
    .S(_02188_),
    .X(_02203_));
 sky130_fd_sc_hd__clkbuf_1 _12530_ (.A(_02203_),
    .X(_01374_));
 sky130_fd_sc_hd__mux2_1 _12531_ (.A0(_06340_),
    .A1(net1520),
    .S(_02188_),
    .X(_02204_));
 sky130_fd_sc_hd__clkbuf_1 _12532_ (.A(_02204_),
    .X(_01375_));
 sky130_fd_sc_hd__mux2_1 _12533_ (.A0(_06342_),
    .A1(net1673),
    .S(_02188_),
    .X(_02205_));
 sky130_fd_sc_hd__clkbuf_1 _12534_ (.A(_02205_),
    .X(_01376_));
 sky130_fd_sc_hd__nor2_4 _12535_ (.A(_06399_),
    .B(_04646_),
    .Y(_02206_));
 sky130_fd_sc_hd__buf_4 _12536_ (.A(_02206_),
    .X(_02207_));
 sky130_fd_sc_hd__mux2_1 _12537_ (.A0(net1440),
    .A1(_04498_),
    .S(_02207_),
    .X(_02208_));
 sky130_fd_sc_hd__clkbuf_1 _12538_ (.A(_02208_),
    .X(_01377_));
 sky130_fd_sc_hd__mux2_1 _12539_ (.A0(net1431),
    .A1(_04505_),
    .S(_02207_),
    .X(_02209_));
 sky130_fd_sc_hd__clkbuf_1 _12540_ (.A(_02209_),
    .X(_01378_));
 sky130_fd_sc_hd__mux2_1 _12541_ (.A0(net806),
    .A1(_04508_),
    .S(_02207_),
    .X(_02210_));
 sky130_fd_sc_hd__clkbuf_1 _12542_ (.A(_02210_),
    .X(_01379_));
 sky130_fd_sc_hd__mux2_1 _12543_ (.A0(net1051),
    .A1(_04511_),
    .S(_02207_),
    .X(_02211_));
 sky130_fd_sc_hd__clkbuf_1 _12544_ (.A(_02211_),
    .X(_01380_));
 sky130_fd_sc_hd__mux2_1 _12545_ (.A0(net43),
    .A1(_04514_),
    .S(_02207_),
    .X(_02212_));
 sky130_fd_sc_hd__clkbuf_1 _12546_ (.A(_02212_),
    .X(_01381_));
 sky130_fd_sc_hd__mux2_1 _12547_ (.A0(net367),
    .A1(_04517_),
    .S(_02207_),
    .X(_02213_));
 sky130_fd_sc_hd__clkbuf_1 _12548_ (.A(_02213_),
    .X(_01382_));
 sky130_fd_sc_hd__mux2_1 _12549_ (.A0(net774),
    .A1(_04520_),
    .S(_02207_),
    .X(_02214_));
 sky130_fd_sc_hd__clkbuf_1 _12550_ (.A(_02214_),
    .X(_01383_));
 sky130_fd_sc_hd__mux2_1 _12551_ (.A0(net194),
    .A1(_04523_),
    .S(_02207_),
    .X(_02215_));
 sky130_fd_sc_hd__clkbuf_1 _12552_ (.A(_02215_),
    .X(_01384_));
 sky130_fd_sc_hd__mux2_1 _12553_ (.A0(net364),
    .A1(_04526_),
    .S(_02207_),
    .X(_02216_));
 sky130_fd_sc_hd__clkbuf_1 _12554_ (.A(_02216_),
    .X(_01385_));
 sky130_fd_sc_hd__mux2_1 _12555_ (.A0(net1443),
    .A1(_04529_),
    .S(_02207_),
    .X(_02217_));
 sky130_fd_sc_hd__clkbuf_1 _12556_ (.A(_02217_),
    .X(_01386_));
 sky130_fd_sc_hd__mux2_1 _12557_ (.A0(net303),
    .A1(_04532_),
    .S(_02206_),
    .X(_02218_));
 sky130_fd_sc_hd__clkbuf_1 _12558_ (.A(_02218_),
    .X(_01387_));
 sky130_fd_sc_hd__mux2_1 _12559_ (.A0(net385),
    .A1(_04535_),
    .S(_02206_),
    .X(_02219_));
 sky130_fd_sc_hd__clkbuf_1 _12560_ (.A(_02219_),
    .X(_01388_));
 sky130_fd_sc_hd__mux2_1 _12561_ (.A0(net1169),
    .A1(_04538_),
    .S(_02206_),
    .X(_02220_));
 sky130_fd_sc_hd__clkbuf_1 _12562_ (.A(_02220_),
    .X(_01389_));
 sky130_fd_sc_hd__mux2_1 _12563_ (.A0(net590),
    .A1(_04541_),
    .S(_02206_),
    .X(_02221_));
 sky130_fd_sc_hd__clkbuf_1 _12564_ (.A(_02221_),
    .X(_01390_));
 sky130_fd_sc_hd__mux2_1 _12565_ (.A0(net396),
    .A1(_04544_),
    .S(_02206_),
    .X(_02222_));
 sky130_fd_sc_hd__clkbuf_1 _12566_ (.A(_02222_),
    .X(_01391_));
 sky130_fd_sc_hd__mux2_1 _12567_ (.A0(net1938),
    .A1(_04547_),
    .S(_02206_),
    .X(_02223_));
 sky130_fd_sc_hd__clkbuf_1 _12568_ (.A(_02223_),
    .X(_01392_));
 sky130_fd_sc_hd__or2_1 _12569_ (.A(_04127_),
    .B(_04325_),
    .X(_02224_));
 sky130_fd_sc_hd__clkbuf_4 _12570_ (.A(_02224_),
    .X(_02225_));
 sky130_fd_sc_hd__buf_4 _12571_ (.A(_02225_),
    .X(_02226_));
 sky130_fd_sc_hd__mux2_1 _12572_ (.A0(_06309_),
    .A1(net423),
    .S(_02226_),
    .X(_02227_));
 sky130_fd_sc_hd__clkbuf_1 _12573_ (.A(_02227_),
    .X(_01393_));
 sky130_fd_sc_hd__mux2_1 _12574_ (.A0(_06314_),
    .A1(net1774),
    .S(_02226_),
    .X(_02228_));
 sky130_fd_sc_hd__clkbuf_1 _12575_ (.A(_02228_),
    .X(_01394_));
 sky130_fd_sc_hd__mux2_1 _12576_ (.A0(_06316_),
    .A1(net1106),
    .S(_02226_),
    .X(_02229_));
 sky130_fd_sc_hd__clkbuf_1 _12577_ (.A(_02229_),
    .X(_01395_));
 sky130_fd_sc_hd__mux2_1 _12578_ (.A0(_06318_),
    .A1(net567),
    .S(_02226_),
    .X(_02230_));
 sky130_fd_sc_hd__clkbuf_1 _12579_ (.A(_02230_),
    .X(_01396_));
 sky130_fd_sc_hd__mux2_1 _12580_ (.A0(_06320_),
    .A1(net813),
    .S(_02226_),
    .X(_02231_));
 sky130_fd_sc_hd__clkbuf_1 _12581_ (.A(_02231_),
    .X(_01397_));
 sky130_fd_sc_hd__mux2_1 _12582_ (.A0(_06322_),
    .A1(net640),
    .S(_02226_),
    .X(_02232_));
 sky130_fd_sc_hd__clkbuf_1 _12583_ (.A(_02232_),
    .X(_01398_));
 sky130_fd_sc_hd__mux2_1 _12584_ (.A0(_06324_),
    .A1(net1226),
    .S(_02226_),
    .X(_02233_));
 sky130_fd_sc_hd__clkbuf_1 _12585_ (.A(_02233_),
    .X(_01399_));
 sky130_fd_sc_hd__mux2_1 _12586_ (.A0(_06326_),
    .A1(net757),
    .S(_02226_),
    .X(_02234_));
 sky130_fd_sc_hd__clkbuf_1 _12587_ (.A(_02234_),
    .X(_01400_));
 sky130_fd_sc_hd__mux2_1 _12588_ (.A0(_06328_),
    .A1(net1365),
    .S(_02226_),
    .X(_02235_));
 sky130_fd_sc_hd__clkbuf_1 _12589_ (.A(_02235_),
    .X(_01401_));
 sky130_fd_sc_hd__mux2_1 _12590_ (.A0(_06330_),
    .A1(net1386),
    .S(_02226_),
    .X(_02236_));
 sky130_fd_sc_hd__clkbuf_1 _12591_ (.A(_02236_),
    .X(_01402_));
 sky130_fd_sc_hd__mux2_1 _12592_ (.A0(_06332_),
    .A1(net1725),
    .S(_02225_),
    .X(_02237_));
 sky130_fd_sc_hd__clkbuf_1 _12593_ (.A(_02237_),
    .X(_01403_));
 sky130_fd_sc_hd__mux2_1 _12594_ (.A0(_06334_),
    .A1(net700),
    .S(_02225_),
    .X(_02238_));
 sky130_fd_sc_hd__clkbuf_1 _12595_ (.A(_02238_),
    .X(_01404_));
 sky130_fd_sc_hd__mux2_1 _12596_ (.A0(_06336_),
    .A1(net1879),
    .S(_02225_),
    .X(_02239_));
 sky130_fd_sc_hd__clkbuf_1 _12597_ (.A(_02239_),
    .X(_01405_));
 sky130_fd_sc_hd__mux2_1 _12598_ (.A0(_06338_),
    .A1(net284),
    .S(_02225_),
    .X(_02240_));
 sky130_fd_sc_hd__clkbuf_1 _12599_ (.A(_02240_),
    .X(_01406_));
 sky130_fd_sc_hd__mux2_1 _12600_ (.A0(_06340_),
    .A1(net800),
    .S(_02225_),
    .X(_02241_));
 sky130_fd_sc_hd__clkbuf_1 _12601_ (.A(_02241_),
    .X(_01407_));
 sky130_fd_sc_hd__mux2_1 _12602_ (.A0(_06342_),
    .A1(net863),
    .S(_02225_),
    .X(_02242_));
 sky130_fd_sc_hd__clkbuf_1 _12603_ (.A(_02242_),
    .X(_01408_));
 sky130_fd_sc_hd__or2_1 _12604_ (.A(_06399_),
    .B(_04684_),
    .X(_02243_));
 sky130_fd_sc_hd__buf_4 _12605_ (.A(_02243_),
    .X(_02244_));
 sky130_fd_sc_hd__buf_4 _12606_ (.A(_02244_),
    .X(_02245_));
 sky130_fd_sc_hd__mux2_1 _12607_ (.A0(_06309_),
    .A1(net1131),
    .S(_02245_),
    .X(_02246_));
 sky130_fd_sc_hd__clkbuf_1 _12608_ (.A(_02246_),
    .X(_01409_));
 sky130_fd_sc_hd__mux2_1 _12609_ (.A0(_06314_),
    .A1(net1115),
    .S(_02245_),
    .X(_02247_));
 sky130_fd_sc_hd__clkbuf_1 _12610_ (.A(_02247_),
    .X(_01410_));
 sky130_fd_sc_hd__mux2_1 _12611_ (.A0(_06316_),
    .A1(net1354),
    .S(_02245_),
    .X(_02248_));
 sky130_fd_sc_hd__clkbuf_1 _12612_ (.A(_02248_),
    .X(_01411_));
 sky130_fd_sc_hd__mux2_1 _12613_ (.A0(_06318_),
    .A1(net878),
    .S(_02245_),
    .X(_02249_));
 sky130_fd_sc_hd__clkbuf_1 _12614_ (.A(_02249_),
    .X(_01412_));
 sky130_fd_sc_hd__mux2_1 _12615_ (.A0(_06320_),
    .A1(net1828),
    .S(_02245_),
    .X(_02250_));
 sky130_fd_sc_hd__clkbuf_1 _12616_ (.A(_02250_),
    .X(_01413_));
 sky130_fd_sc_hd__mux2_1 _12617_ (.A0(_06322_),
    .A1(net727),
    .S(_02245_),
    .X(_02251_));
 sky130_fd_sc_hd__clkbuf_1 _12618_ (.A(_02251_),
    .X(_01414_));
 sky130_fd_sc_hd__mux2_1 _12619_ (.A0(_06324_),
    .A1(net1570),
    .S(_02245_),
    .X(_02252_));
 sky130_fd_sc_hd__clkbuf_1 _12620_ (.A(_02252_),
    .X(_01415_));
 sky130_fd_sc_hd__mux2_1 _12621_ (.A0(_06326_),
    .A1(net740),
    .S(_02245_),
    .X(_02253_));
 sky130_fd_sc_hd__clkbuf_1 _12622_ (.A(_02253_),
    .X(_01416_));
 sky130_fd_sc_hd__mux2_1 _12623_ (.A0(_06328_),
    .A1(net1389),
    .S(_02245_),
    .X(_02254_));
 sky130_fd_sc_hd__clkbuf_1 _12624_ (.A(_02254_),
    .X(_01417_));
 sky130_fd_sc_hd__mux2_1 _12625_ (.A0(_06330_),
    .A1(net1664),
    .S(_02245_),
    .X(_02255_));
 sky130_fd_sc_hd__clkbuf_1 _12626_ (.A(_02255_),
    .X(_01418_));
 sky130_fd_sc_hd__mux2_1 _12627_ (.A0(_06332_),
    .A1(net1284),
    .S(_02244_),
    .X(_02256_));
 sky130_fd_sc_hd__clkbuf_1 _12628_ (.A(_02256_),
    .X(_01419_));
 sky130_fd_sc_hd__mux2_1 _12629_ (.A0(_06334_),
    .A1(net888),
    .S(_02244_),
    .X(_02257_));
 sky130_fd_sc_hd__clkbuf_1 _12630_ (.A(_02257_),
    .X(_01420_));
 sky130_fd_sc_hd__mux2_1 _12631_ (.A0(_06336_),
    .A1(net549),
    .S(_02244_),
    .X(_02258_));
 sky130_fd_sc_hd__clkbuf_1 _12632_ (.A(_02258_),
    .X(_01421_));
 sky130_fd_sc_hd__mux2_1 _12633_ (.A0(_06338_),
    .A1(net1359),
    .S(_02244_),
    .X(_02259_));
 sky130_fd_sc_hd__clkbuf_1 _12634_ (.A(_02259_),
    .X(_01422_));
 sky130_fd_sc_hd__mux2_1 _12635_ (.A0(_06340_),
    .A1(net566),
    .S(_02244_),
    .X(_02260_));
 sky130_fd_sc_hd__clkbuf_1 _12636_ (.A(_02260_),
    .X(_01423_));
 sky130_fd_sc_hd__mux2_1 _12637_ (.A0(_06342_),
    .A1(net706),
    .S(_02244_),
    .X(_02261_));
 sky130_fd_sc_hd__clkbuf_1 _12638_ (.A(_02261_),
    .X(_01424_));
 sky130_fd_sc_hd__or3_1 _12639_ (.A(_02506_),
    .B(_02644_),
    .C(_04325_),
    .X(_02262_));
 sky130_fd_sc_hd__buf_4 _12640_ (.A(_02262_),
    .X(_02263_));
 sky130_fd_sc_hd__buf_4 _12641_ (.A(_02263_),
    .X(_02264_));
 sky130_fd_sc_hd__mux2_1 _12642_ (.A0(_06309_),
    .A1(net1357),
    .S(_02264_),
    .X(_02265_));
 sky130_fd_sc_hd__clkbuf_1 _12643_ (.A(_02265_),
    .X(_01425_));
 sky130_fd_sc_hd__mux2_1 _12644_ (.A0(_06314_),
    .A1(net893),
    .S(_02264_),
    .X(_02266_));
 sky130_fd_sc_hd__clkbuf_1 _12645_ (.A(_02266_),
    .X(_01426_));
 sky130_fd_sc_hd__mux2_1 _12646_ (.A0(_06316_),
    .A1(net1425),
    .S(_02264_),
    .X(_02267_));
 sky130_fd_sc_hd__clkbuf_1 _12647_ (.A(_02267_),
    .X(_01427_));
 sky130_fd_sc_hd__mux2_1 _12648_ (.A0(_06318_),
    .A1(net1063),
    .S(_02264_),
    .X(_02268_));
 sky130_fd_sc_hd__clkbuf_1 _12649_ (.A(_02268_),
    .X(_01428_));
 sky130_fd_sc_hd__mux2_1 _12650_ (.A0(_06320_),
    .A1(net1411),
    .S(_02264_),
    .X(_02269_));
 sky130_fd_sc_hd__clkbuf_1 _12651_ (.A(_02269_),
    .X(_01429_));
 sky130_fd_sc_hd__mux2_1 _12652_ (.A0(_06322_),
    .A1(net1202),
    .S(_02264_),
    .X(_02270_));
 sky130_fd_sc_hd__clkbuf_1 _12653_ (.A(_02270_),
    .X(_01430_));
 sky130_fd_sc_hd__mux2_1 _12654_ (.A0(_06324_),
    .A1(net919),
    .S(_02264_),
    .X(_02271_));
 sky130_fd_sc_hd__clkbuf_1 _12655_ (.A(_02271_),
    .X(_01431_));
 sky130_fd_sc_hd__mux2_1 _12656_ (.A0(_06326_),
    .A1(net1677),
    .S(_02264_),
    .X(_02272_));
 sky130_fd_sc_hd__clkbuf_1 _12657_ (.A(_02272_),
    .X(_01432_));
 sky130_fd_sc_hd__mux2_1 _12658_ (.A0(_06328_),
    .A1(net1134),
    .S(_02264_),
    .X(_02273_));
 sky130_fd_sc_hd__clkbuf_1 _12659_ (.A(_02273_),
    .X(_01433_));
 sky130_fd_sc_hd__mux2_1 _12660_ (.A0(_06330_),
    .A1(net1522),
    .S(_02264_),
    .X(_02274_));
 sky130_fd_sc_hd__clkbuf_1 _12661_ (.A(_02274_),
    .X(_01434_));
 sky130_fd_sc_hd__mux2_1 _12662_ (.A0(_06332_),
    .A1(net1630),
    .S(_02263_),
    .X(_02275_));
 sky130_fd_sc_hd__clkbuf_1 _12663_ (.A(_02275_),
    .X(_01435_));
 sky130_fd_sc_hd__mux2_1 _12664_ (.A0(_06334_),
    .A1(net991),
    .S(_02263_),
    .X(_02276_));
 sky130_fd_sc_hd__clkbuf_1 _12665_ (.A(_02276_),
    .X(_01436_));
 sky130_fd_sc_hd__mux2_1 _12666_ (.A0(_06336_),
    .A1(net1028),
    .S(_02263_),
    .X(_02277_));
 sky130_fd_sc_hd__clkbuf_1 _12667_ (.A(_02277_),
    .X(_01437_));
 sky130_fd_sc_hd__mux2_1 _12668_ (.A0(_06338_),
    .A1(net449),
    .S(_02263_),
    .X(_02278_));
 sky130_fd_sc_hd__clkbuf_1 _12669_ (.A(_02278_),
    .X(_01438_));
 sky130_fd_sc_hd__mux2_1 _12670_ (.A0(_06340_),
    .A1(net1340),
    .S(_02263_),
    .X(_02279_));
 sky130_fd_sc_hd__clkbuf_1 _12671_ (.A(_02279_),
    .X(_01439_));
 sky130_fd_sc_hd__mux2_1 _12672_ (.A0(_06342_),
    .A1(net1399),
    .S(_02263_),
    .X(_02280_));
 sky130_fd_sc_hd__clkbuf_1 _12673_ (.A(_02280_),
    .X(_01440_));
 sky130_fd_sc_hd__or2_1 _12674_ (.A(_06399_),
    .B(_04365_),
    .X(_02281_));
 sky130_fd_sc_hd__clkbuf_4 _12675_ (.A(_02281_),
    .X(_02282_));
 sky130_fd_sc_hd__buf_4 _12676_ (.A(_02282_),
    .X(_02283_));
 sky130_fd_sc_hd__mux2_1 _12677_ (.A0(_04070_),
    .A1(net1583),
    .S(_02283_),
    .X(_02284_));
 sky130_fd_sc_hd__clkbuf_1 _12678_ (.A(_02284_),
    .X(_01441_));
 sky130_fd_sc_hd__mux2_1 _12679_ (.A0(_04081_),
    .A1(net661),
    .S(_02283_),
    .X(_02285_));
 sky130_fd_sc_hd__clkbuf_1 _12680_ (.A(_02285_),
    .X(_01442_));
 sky130_fd_sc_hd__mux2_1 _12681_ (.A0(_04084_),
    .A1(net1133),
    .S(_02283_),
    .X(_02286_));
 sky130_fd_sc_hd__clkbuf_1 _12682_ (.A(_02286_),
    .X(_01443_));
 sky130_fd_sc_hd__mux2_1 _12683_ (.A0(_04087_),
    .A1(net221),
    .S(_02283_),
    .X(_02287_));
 sky130_fd_sc_hd__clkbuf_1 _12684_ (.A(_02287_),
    .X(_01444_));
 sky130_fd_sc_hd__mux2_1 _12685_ (.A0(_04090_),
    .A1(net770),
    .S(_02283_),
    .X(_02288_));
 sky130_fd_sc_hd__clkbuf_1 _12686_ (.A(_02288_),
    .X(_01445_));
 sky130_fd_sc_hd__mux2_1 _12687_ (.A0(_04093_),
    .A1(net553),
    .S(_02283_),
    .X(_02289_));
 sky130_fd_sc_hd__clkbuf_1 _12688_ (.A(_02289_),
    .X(_01446_));
 sky130_fd_sc_hd__mux2_1 _12689_ (.A0(_04096_),
    .A1(net1360),
    .S(_02283_),
    .X(_02290_));
 sky130_fd_sc_hd__clkbuf_1 _12690_ (.A(_02290_),
    .X(_01447_));
 sky130_fd_sc_hd__mux2_1 _12691_ (.A0(_04099_),
    .A1(net796),
    .S(_02283_),
    .X(_02291_));
 sky130_fd_sc_hd__clkbuf_1 _12692_ (.A(_02291_),
    .X(_01448_));
 sky130_fd_sc_hd__mux2_1 _12693_ (.A0(_04102_),
    .A1(net637),
    .S(_02283_),
    .X(_02292_));
 sky130_fd_sc_hd__clkbuf_1 _12694_ (.A(_02292_),
    .X(_01449_));
 sky130_fd_sc_hd__mux2_1 _12695_ (.A0(_04105_),
    .A1(net1707),
    .S(_02283_),
    .X(_02293_));
 sky130_fd_sc_hd__clkbuf_1 _12696_ (.A(_02293_),
    .X(_01450_));
 sky130_fd_sc_hd__mux2_1 _12697_ (.A0(_04108_),
    .A1(net1172),
    .S(_02282_),
    .X(_02294_));
 sky130_fd_sc_hd__clkbuf_1 _12698_ (.A(_02294_),
    .X(_01451_));
 sky130_fd_sc_hd__mux2_1 _12699_ (.A0(_04111_),
    .A1(net474),
    .S(_02282_),
    .X(_02295_));
 sky130_fd_sc_hd__clkbuf_1 _12700_ (.A(_02295_),
    .X(_01452_));
 sky130_fd_sc_hd__mux2_1 _12701_ (.A0(_04114_),
    .A1(net868),
    .S(_02282_),
    .X(_02296_));
 sky130_fd_sc_hd__clkbuf_1 _12702_ (.A(_02296_),
    .X(_01453_));
 sky130_fd_sc_hd__mux2_1 _12703_ (.A0(_04117_),
    .A1(net624),
    .S(_02282_),
    .X(_02297_));
 sky130_fd_sc_hd__clkbuf_1 _12704_ (.A(_02297_),
    .X(_01454_));
 sky130_fd_sc_hd__mux2_1 _12705_ (.A0(_04120_),
    .A1(net1201),
    .S(_02282_),
    .X(_02298_));
 sky130_fd_sc_hd__clkbuf_1 _12706_ (.A(_02298_),
    .X(_01455_));
 sky130_fd_sc_hd__mux2_1 _12707_ (.A0(_04123_),
    .A1(net1194),
    .S(_02282_),
    .X(_02299_));
 sky130_fd_sc_hd__clkbuf_1 _12708_ (.A(_02299_),
    .X(_01456_));
 sky130_fd_sc_hd__or3_1 _12709_ (.A(_02484_),
    .B(_02737_),
    .C(_04325_),
    .X(_02300_));
 sky130_fd_sc_hd__clkbuf_4 _12710_ (.A(_02300_),
    .X(_02301_));
 sky130_fd_sc_hd__buf_4 _12711_ (.A(_02301_),
    .X(_02302_));
 sky130_fd_sc_hd__mux2_1 _12712_ (.A0(_04070_),
    .A1(net1298),
    .S(_02302_),
    .X(_02303_));
 sky130_fd_sc_hd__clkbuf_1 _12713_ (.A(_02303_),
    .X(_01457_));
 sky130_fd_sc_hd__mux2_1 _12714_ (.A0(_04081_),
    .A1(net1136),
    .S(_02302_),
    .X(_02304_));
 sky130_fd_sc_hd__clkbuf_1 _12715_ (.A(_02304_),
    .X(_01458_));
 sky130_fd_sc_hd__mux2_1 _12716_ (.A0(_04084_),
    .A1(net791),
    .S(_02302_),
    .X(_02305_));
 sky130_fd_sc_hd__clkbuf_1 _12717_ (.A(_02305_),
    .X(_01459_));
 sky130_fd_sc_hd__mux2_1 _12718_ (.A0(_04087_),
    .A1(net348),
    .S(_02302_),
    .X(_02306_));
 sky130_fd_sc_hd__clkbuf_1 _12719_ (.A(_02306_),
    .X(_01460_));
 sky130_fd_sc_hd__mux2_1 _12720_ (.A0(_04090_),
    .A1(net1575),
    .S(_02302_),
    .X(_02307_));
 sky130_fd_sc_hd__clkbuf_1 _12721_ (.A(_02307_),
    .X(_01461_));
 sky130_fd_sc_hd__mux2_1 _12722_ (.A0(_04093_),
    .A1(net436),
    .S(_02302_),
    .X(_02308_));
 sky130_fd_sc_hd__clkbuf_1 _12723_ (.A(_02308_),
    .X(_01462_));
 sky130_fd_sc_hd__mux2_1 _12724_ (.A0(_04096_),
    .A1(net569),
    .S(_02302_),
    .X(_02309_));
 sky130_fd_sc_hd__clkbuf_1 _12725_ (.A(_02309_),
    .X(_01463_));
 sky130_fd_sc_hd__mux2_1 _12726_ (.A0(_04099_),
    .A1(net1468),
    .S(_02302_),
    .X(_02310_));
 sky130_fd_sc_hd__clkbuf_1 _12727_ (.A(_02310_),
    .X(_01464_));
 sky130_fd_sc_hd__mux2_1 _12728_ (.A0(_04102_),
    .A1(net1250),
    .S(_02302_),
    .X(_02311_));
 sky130_fd_sc_hd__clkbuf_1 _12729_ (.A(_02311_),
    .X(_01465_));
 sky130_fd_sc_hd__mux2_1 _12730_ (.A0(_04105_),
    .A1(net1262),
    .S(_02302_),
    .X(_02312_));
 sky130_fd_sc_hd__clkbuf_1 _12731_ (.A(_02312_),
    .X(_01466_));
 sky130_fd_sc_hd__mux2_1 _12732_ (.A0(_04108_),
    .A1(net667),
    .S(_02301_),
    .X(_02313_));
 sky130_fd_sc_hd__clkbuf_1 _12733_ (.A(_02313_),
    .X(_01467_));
 sky130_fd_sc_hd__mux2_1 _12734_ (.A0(_04111_),
    .A1(net1210),
    .S(_02301_),
    .X(_02314_));
 sky130_fd_sc_hd__clkbuf_1 _12735_ (.A(_02314_),
    .X(_01468_));
 sky130_fd_sc_hd__mux2_1 _12736_ (.A0(_04114_),
    .A1(net1517),
    .S(_02301_),
    .X(_02315_));
 sky130_fd_sc_hd__clkbuf_1 _12737_ (.A(_02315_),
    .X(_01469_));
 sky130_fd_sc_hd__mux2_1 _12738_ (.A0(_04117_),
    .A1(net1035),
    .S(_02301_),
    .X(_02316_));
 sky130_fd_sc_hd__clkbuf_1 _12739_ (.A(_02316_),
    .X(_01470_));
 sky130_fd_sc_hd__mux2_1 _12740_ (.A0(_04120_),
    .A1(net410),
    .S(_02301_),
    .X(_02317_));
 sky130_fd_sc_hd__clkbuf_1 _12741_ (.A(_02317_),
    .X(_01471_));
 sky130_fd_sc_hd__mux2_1 _12742_ (.A0(_04123_),
    .A1(net677),
    .S(_02301_),
    .X(_02318_));
 sky130_fd_sc_hd__clkbuf_1 _12743_ (.A(_02318_),
    .X(_01472_));
 sky130_fd_sc_hd__nand2b_4 _12744_ (.A_N(_06399_),
    .B(_04408_),
    .Y(_02319_));
 sky130_fd_sc_hd__buf_4 _12745_ (.A(_02319_),
    .X(_02320_));
 sky130_fd_sc_hd__mux2_1 _12746_ (.A0(_04070_),
    .A1(net1978),
    .S(_02320_),
    .X(_02321_));
 sky130_fd_sc_hd__clkbuf_1 _12747_ (.A(_02321_),
    .X(_01473_));
 sky130_fd_sc_hd__mux2_1 _12748_ (.A0(_04081_),
    .A1(net1521),
    .S(_02320_),
    .X(_02322_));
 sky130_fd_sc_hd__clkbuf_1 _12749_ (.A(_02322_),
    .X(_01474_));
 sky130_fd_sc_hd__mux2_1 _12750_ (.A0(_04084_),
    .A1(net1602),
    .S(_02320_),
    .X(_02323_));
 sky130_fd_sc_hd__clkbuf_1 _12751_ (.A(_02323_),
    .X(_01475_));
 sky130_fd_sc_hd__mux2_1 _12752_ (.A0(_04087_),
    .A1(net1286),
    .S(_02320_),
    .X(_02324_));
 sky130_fd_sc_hd__clkbuf_1 _12753_ (.A(_02324_),
    .X(_01476_));
 sky130_fd_sc_hd__mux2_1 _12754_ (.A0(_04090_),
    .A1(net930),
    .S(_02320_),
    .X(_02325_));
 sky130_fd_sc_hd__clkbuf_1 _12755_ (.A(_02325_),
    .X(_01477_));
 sky130_fd_sc_hd__mux2_1 _12756_ (.A0(_04093_),
    .A1(net514),
    .S(_02320_),
    .X(_02326_));
 sky130_fd_sc_hd__clkbuf_1 _12757_ (.A(_02326_),
    .X(_01478_));
 sky130_fd_sc_hd__mux2_1 _12758_ (.A0(_04096_),
    .A1(net1214),
    .S(_02320_),
    .X(_02327_));
 sky130_fd_sc_hd__clkbuf_1 _12759_ (.A(_02327_),
    .X(_01479_));
 sky130_fd_sc_hd__mux2_1 _12760_ (.A0(_04099_),
    .A1(net1269),
    .S(_02320_),
    .X(_02328_));
 sky130_fd_sc_hd__clkbuf_1 _12761_ (.A(_02328_),
    .X(_01480_));
 sky130_fd_sc_hd__mux2_1 _12762_ (.A0(_04102_),
    .A1(net955),
    .S(_02320_),
    .X(_02329_));
 sky130_fd_sc_hd__clkbuf_1 _12763_ (.A(_02329_),
    .X(_01481_));
 sky130_fd_sc_hd__mux2_1 _12764_ (.A0(_04105_),
    .A1(net1013),
    .S(_02320_),
    .X(_02330_));
 sky130_fd_sc_hd__clkbuf_1 _12765_ (.A(_02330_),
    .X(_01482_));
 sky130_fd_sc_hd__mux2_1 _12766_ (.A0(_04108_),
    .A1(net641),
    .S(_02319_),
    .X(_02331_));
 sky130_fd_sc_hd__clkbuf_1 _12767_ (.A(_02331_),
    .X(_01483_));
 sky130_fd_sc_hd__mux2_1 _12768_ (.A0(_04111_),
    .A1(net407),
    .S(_02319_),
    .X(_02332_));
 sky130_fd_sc_hd__clkbuf_1 _12769_ (.A(_02332_),
    .X(_01484_));
 sky130_fd_sc_hd__mux2_1 _12770_ (.A0(_04114_),
    .A1(net1670),
    .S(_02319_),
    .X(_02333_));
 sky130_fd_sc_hd__clkbuf_1 _12771_ (.A(_02333_),
    .X(_01485_));
 sky130_fd_sc_hd__mux2_1 _12772_ (.A0(_04117_),
    .A1(net568),
    .S(_02319_),
    .X(_02334_));
 sky130_fd_sc_hd__clkbuf_1 _12773_ (.A(_02334_),
    .X(_01486_));
 sky130_fd_sc_hd__mux2_1 _12774_ (.A0(_04120_),
    .A1(net1339),
    .S(_02319_),
    .X(_02335_));
 sky130_fd_sc_hd__clkbuf_1 _12775_ (.A(_02335_),
    .X(_01487_));
 sky130_fd_sc_hd__mux2_1 _12776_ (.A0(_04123_),
    .A1(net622),
    .S(_02319_),
    .X(_02336_));
 sky130_fd_sc_hd__clkbuf_1 _12777_ (.A(_02336_),
    .X(_01488_));
 sky130_fd_sc_hd__nor2_4 _12778_ (.A(_04127_),
    .B(_04368_),
    .Y(_02337_));
 sky130_fd_sc_hd__buf_4 _12779_ (.A(_02337_),
    .X(_02338_));
 sky130_fd_sc_hd__mux2_1 _12780_ (.A0(net2034),
    .A1(_04498_),
    .S(_02338_),
    .X(_02339_));
 sky130_fd_sc_hd__clkbuf_1 _12781_ (.A(_02339_),
    .X(_01489_));
 sky130_fd_sc_hd__mux2_1 _12782_ (.A0(net815),
    .A1(_04505_),
    .S(_02338_),
    .X(_02340_));
 sky130_fd_sc_hd__clkbuf_1 _12783_ (.A(_02340_),
    .X(_01490_));
 sky130_fd_sc_hd__mux2_1 _12784_ (.A0(net1702),
    .A1(_04508_),
    .S(_02338_),
    .X(_02341_));
 sky130_fd_sc_hd__clkbuf_1 _12785_ (.A(_02341_),
    .X(_01491_));
 sky130_fd_sc_hd__mux2_1 _12786_ (.A0(net1024),
    .A1(_04511_),
    .S(_02338_),
    .X(_02342_));
 sky130_fd_sc_hd__clkbuf_1 _12787_ (.A(_02342_),
    .X(_01492_));
 sky130_fd_sc_hd__mux2_1 _12788_ (.A0(net542),
    .A1(_04514_),
    .S(_02338_),
    .X(_02343_));
 sky130_fd_sc_hd__clkbuf_1 _12789_ (.A(_02343_),
    .X(_01493_));
 sky130_fd_sc_hd__mux2_1 _12790_ (.A0(net45),
    .A1(_04517_),
    .S(_02338_),
    .X(_02344_));
 sky130_fd_sc_hd__clkbuf_1 _12791_ (.A(_02344_),
    .X(_01494_));
 sky130_fd_sc_hd__mux2_1 _12792_ (.A0(net993),
    .A1(_04520_),
    .S(_02338_),
    .X(_02345_));
 sky130_fd_sc_hd__clkbuf_1 _12793_ (.A(_02345_),
    .X(_01495_));
 sky130_fd_sc_hd__mux2_1 _12794_ (.A0(net994),
    .A1(_04523_),
    .S(_02338_),
    .X(_02346_));
 sky130_fd_sc_hd__clkbuf_1 _12795_ (.A(_02346_),
    .X(_01496_));
 sky130_fd_sc_hd__mux2_1 _12796_ (.A0(net1057),
    .A1(_04526_),
    .S(_02338_),
    .X(_02347_));
 sky130_fd_sc_hd__clkbuf_1 _12797_ (.A(_02347_),
    .X(_01497_));
 sky130_fd_sc_hd__mux2_1 _12798_ (.A0(net574),
    .A1(_04529_),
    .S(_02338_),
    .X(_02348_));
 sky130_fd_sc_hd__clkbuf_1 _12799_ (.A(_02348_),
    .X(_01498_));
 sky130_fd_sc_hd__mux2_1 _12800_ (.A0(net1705),
    .A1(_04532_),
    .S(_02337_),
    .X(_02349_));
 sky130_fd_sc_hd__clkbuf_1 _12801_ (.A(_02349_),
    .X(_01499_));
 sky130_fd_sc_hd__mux2_1 _12802_ (.A0(net1397),
    .A1(_04535_),
    .S(_02337_),
    .X(_02350_));
 sky130_fd_sc_hd__clkbuf_1 _12803_ (.A(_02350_),
    .X(_01500_));
 sky130_fd_sc_hd__mux2_1 _12804_ (.A0(net1491),
    .A1(_04538_),
    .S(_02337_),
    .X(_02351_));
 sky130_fd_sc_hd__clkbuf_1 _12805_ (.A(_02351_),
    .X(_01501_));
 sky130_fd_sc_hd__mux2_1 _12806_ (.A0(net808),
    .A1(_04541_),
    .S(_02337_),
    .X(_02352_));
 sky130_fd_sc_hd__clkbuf_1 _12807_ (.A(_02352_),
    .X(_01502_));
 sky130_fd_sc_hd__mux2_1 _12808_ (.A0(net699),
    .A1(_04544_),
    .S(_02337_),
    .X(_02353_));
 sky130_fd_sc_hd__clkbuf_1 _12809_ (.A(_02353_),
    .X(_01503_));
 sky130_fd_sc_hd__mux2_1 _12810_ (.A0(net816),
    .A1(_04547_),
    .S(_02337_),
    .X(_02354_));
 sky130_fd_sc_hd__clkbuf_1 _12811_ (.A(_02354_),
    .X(_01504_));
 sky130_fd_sc_hd__dfxtp_1 _12812_ (.CLK(clknet_leaf_106_i_clk),
    .D(_01505_),
    .Q(\mem[49][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12813_ (.CLK(clknet_leaf_109_i_clk),
    .D(_01506_),
    .Q(\mem[49][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12814_ (.CLK(clknet_leaf_105_i_clk),
    .D(_01507_),
    .Q(\mem[49][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12815_ (.CLK(clknet_leaf_110_i_clk),
    .D(_01508_),
    .Q(\mem[49][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12816_ (.CLK(clknet_leaf_106_i_clk),
    .D(_01509_),
    .Q(\mem[49][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12817_ (.CLK(clknet_leaf_107_i_clk),
    .D(_01510_),
    .Q(\mem[49][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12818_ (.CLK(clknet_leaf_106_i_clk),
    .D(_01511_),
    .Q(\mem[49][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12819_ (.CLK(clknet_leaf_107_i_clk),
    .D(_01512_),
    .Q(\mem[49][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12820_ (.CLK(clknet_leaf_107_i_clk),
    .D(_01513_),
    .Q(\mem[49][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12821_ (.CLK(clknet_leaf_106_i_clk),
    .D(_01514_),
    .Q(\mem[49][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12822_ (.CLK(clknet_leaf_105_i_clk),
    .D(_01515_),
    .Q(\mem[49][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12823_ (.CLK(clknet_leaf_107_i_clk),
    .D(_01516_),
    .Q(\mem[49][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12824_ (.CLK(clknet_leaf_100_i_clk),
    .D(_01517_),
    .Q(\mem[49][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12825_ (.CLK(clknet_leaf_107_i_clk),
    .D(_01518_),
    .Q(\mem[49][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12826_ (.CLK(clknet_leaf_100_i_clk),
    .D(_01519_),
    .Q(\mem[49][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12827_ (.CLK(clknet_leaf_100_i_clk),
    .D(_01520_),
    .Q(\mem[49][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12828_ (.CLK(clknet_leaf_219_i_clk),
    .D(_01521_),
    .Q(\mem[89][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12829_ (.CLK(clknet_leaf_206_i_clk),
    .D(_01522_),
    .Q(\mem[89][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12830_ (.CLK(clknet_leaf_218_i_clk),
    .D(_01523_),
    .Q(\mem[89][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12831_ (.CLK(clknet_leaf_219_i_clk),
    .D(_01524_),
    .Q(\mem[89][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12832_ (.CLK(clknet_leaf_216_i_clk),
    .D(_01525_),
    .Q(\mem[89][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12833_ (.CLK(clknet_leaf_207_i_clk),
    .D(_01526_),
    .Q(\mem[89][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12834_ (.CLK(clknet_leaf_207_i_clk),
    .D(_01527_),
    .Q(\mem[89][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12835_ (.CLK(clknet_leaf_217_i_clk),
    .D(_01528_),
    .Q(\mem[89][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12836_ (.CLK(clknet_leaf_212_i_clk),
    .D(_01529_),
    .Q(\mem[89][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12837_ (.CLK(clknet_leaf_212_i_clk),
    .D(_01530_),
    .Q(\mem[89][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12838_ (.CLK(clknet_leaf_209_i_clk),
    .D(_01531_),
    .Q(\mem[89][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12839_ (.CLK(clknet_leaf_244_i_clk),
    .D(_01532_),
    .Q(\mem[89][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12840_ (.CLK(clknet_leaf_211_i_clk),
    .D(_01533_),
    .Q(\mem[89][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12841_ (.CLK(clknet_leaf_186_i_clk),
    .D(_01534_),
    .Q(\mem[89][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12842_ (.CLK(clknet_leaf_206_i_clk),
    .D(_01535_),
    .Q(\mem[89][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12843_ (.CLK(clknet_leaf_206_i_clk),
    .D(_01536_),
    .Q(\mem[89][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12844_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01537_),
    .Q(\mem[59][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12845_ (.CLK(clknet_leaf_70_i_clk),
    .D(_01538_),
    .Q(\mem[59][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12846_ (.CLK(clknet_leaf_76_i_clk),
    .D(_01539_),
    .Q(\mem[59][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12847_ (.CLK(clknet_leaf_72_i_clk),
    .D(_01540_),
    .Q(\mem[59][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12848_ (.CLK(clknet_leaf_72_i_clk),
    .D(_01541_),
    .Q(\mem[59][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12849_ (.CLK(clknet_leaf_70_i_clk),
    .D(_01542_),
    .Q(\mem[59][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12850_ (.CLK(clknet_leaf_71_i_clk),
    .D(_01543_),
    .Q(\mem[59][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12851_ (.CLK(clknet_leaf_83_i_clk),
    .D(_01544_),
    .Q(\mem[59][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12852_ (.CLK(clknet_leaf_78_i_clk),
    .D(_01545_),
    .Q(\mem[59][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12853_ (.CLK(clknet_leaf_78_i_clk),
    .D(_01546_),
    .Q(\mem[59][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12854_ (.CLK(clknet_leaf_81_i_clk),
    .D(_01547_),
    .Q(\mem[59][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12855_ (.CLK(clknet_leaf_81_i_clk),
    .D(_01548_),
    .Q(\mem[59][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12856_ (.CLK(clknet_leaf_82_i_clk),
    .D(_01549_),
    .Q(\mem[59][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12857_ (.CLK(clknet_leaf_85_i_clk),
    .D(_01550_),
    .Q(\mem[59][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12858_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01551_),
    .Q(\mem[59][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12859_ (.CLK(clknet_leaf_82_i_clk),
    .D(_01552_),
    .Q(\mem[59][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12860_ (.CLK(clknet_leaf_123_i_clk),
    .D(_01553_),
    .Q(\mem[69][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12861_ (.CLK(clknet_leaf_175_i_clk),
    .D(_01554_),
    .Q(\mem[69][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12862_ (.CLK(clknet_leaf_123_i_clk),
    .D(_01555_),
    .Q(\mem[69][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12863_ (.CLK(clknet_leaf_123_i_clk),
    .D(_01556_),
    .Q(\mem[69][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12864_ (.CLK(clknet_leaf_123_i_clk),
    .D(_01557_),
    .Q(\mem[69][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12865_ (.CLK(clknet_leaf_179_i_clk),
    .D(_01558_),
    .Q(\mem[69][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12866_ (.CLK(clknet_leaf_174_i_clk),
    .D(_01559_),
    .Q(\mem[69][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12867_ (.CLK(clknet_leaf_123_i_clk),
    .D(_01560_),
    .Q(\mem[69][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12868_ (.CLK(clknet_leaf_122_i_clk),
    .D(_01561_),
    .Q(\mem[69][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12869_ (.CLK(clknet_leaf_120_i_clk),
    .D(_01562_),
    .Q(\mem[69][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12870_ (.CLK(clknet_leaf_158_i_clk),
    .D(_01563_),
    .Q(\mem[69][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12871_ (.CLK(clknet_leaf_174_i_clk),
    .D(_01564_),
    .Q(\mem[69][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12872_ (.CLK(clknet_leaf_158_i_clk),
    .D(_01565_),
    .Q(\mem[69][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12873_ (.CLK(clknet_leaf_174_i_clk),
    .D(_01566_),
    .Q(\mem[69][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12874_ (.CLK(clknet_leaf_172_i_clk),
    .D(_01567_),
    .Q(\mem[69][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12875_ (.CLK(clknet_leaf_121_i_clk),
    .D(_01568_),
    .Q(\mem[69][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12876_ (.CLK(clknet_leaf_202_i_clk),
    .D(_01569_),
    .Q(\mem[79][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12877_ (.CLK(clknet_leaf_196_i_clk),
    .D(_01570_),
    .Q(\mem[79][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12878_ (.CLK(clknet_leaf_202_i_clk),
    .D(_01571_),
    .Q(\mem[79][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12879_ (.CLK(clknet_leaf_202_i_clk),
    .D(_01572_),
    .Q(\mem[79][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12880_ (.CLK(clknet_leaf_199_i_clk),
    .D(_01573_),
    .Q(\mem[79][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12881_ (.CLK(clknet_leaf_195_i_clk),
    .D(_01574_),
    .Q(\mem[79][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12882_ (.CLK(clknet_leaf_192_i_clk),
    .D(_01575_),
    .Q(\mem[79][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12883_ (.CLK(clknet_leaf_202_i_clk),
    .D(_01576_),
    .Q(\mem[79][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12884_ (.CLK(clknet_leaf_202_i_clk),
    .D(_01577_),
    .Q(\mem[79][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12885_ (.CLK(clknet_leaf_197_i_clk),
    .D(_01578_),
    .Q(\mem[79][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12886_ (.CLK(clknet_leaf_194_i_clk),
    .D(_01579_),
    .Q(\mem[79][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12887_ (.CLK(clknet_leaf_184_i_clk),
    .D(_01580_),
    .Q(\mem[79][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12888_ (.CLK(clknet_leaf_194_i_clk),
    .D(_01581_),
    .Q(\mem[79][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12889_ (.CLK(clknet_leaf_185_i_clk),
    .D(_01582_),
    .Q(\mem[79][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12890_ (.CLK(clknet_leaf_194_i_clk),
    .D(_01583_),
    .Q(\mem[79][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12891_ (.CLK(clknet_leaf_185_i_clk),
    .D(_01584_),
    .Q(\mem[79][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12892_ (.CLK(clknet_leaf_240_i_clk),
    .D(_01585_),
    .Q(\mem[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12893_ (.CLK(clknet_leaf_257_i_clk),
    .D(_01586_),
    .Q(\mem[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12894_ (.CLK(clknet_leaf_239_i_clk),
    .D(_01587_),
    .Q(\mem[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12895_ (.CLK(clknet_leaf_267_i_clk),
    .D(_01588_),
    .Q(\mem[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12896_ (.CLK(clknet_leaf_267_i_clk),
    .D(_01589_),
    .Q(\mem[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12897_ (.CLK(clknet_leaf_258_i_clk),
    .D(_01590_),
    .Q(\mem[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12898_ (.CLK(clknet_leaf_267_i_clk),
    .D(_01591_),
    .Q(\mem[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12899_ (.CLK(clknet_leaf_270_i_clk),
    .D(_01592_),
    .Q(\mem[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12900_ (.CLK(clknet_leaf_270_i_clk),
    .D(_01593_),
    .Q(\mem[19][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12901_ (.CLK(clknet_leaf_237_i_clk),
    .D(_01594_),
    .Q(\mem[19][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12902_ (.CLK(clknet_leaf_240_i_clk),
    .D(_01595_),
    .Q(\mem[19][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12903_ (.CLK(clknet_leaf_237_i_clk),
    .D(_01596_),
    .Q(\mem[19][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12904_ (.CLK(clknet_leaf_228_i_clk),
    .D(_01597_),
    .Q(\mem[19][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12905_ (.CLK(clknet_leaf_246_i_clk),
    .D(_01598_),
    .Q(\mem[19][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12906_ (.CLK(clknet_leaf_228_i_clk),
    .D(_01599_),
    .Q(\mem[19][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12907_ (.CLK(clknet_leaf_229_i_clk),
    .D(_01600_),
    .Q(\mem[19][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12908_ (.CLK(clknet_leaf_6_i_clk),
    .D(_01601_),
    .Q(\mem[39][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12909_ (.CLK(clknet_leaf_26_i_clk),
    .D(_01602_),
    .Q(\mem[39][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12910_ (.CLK(clknet_leaf_286_i_clk),
    .D(_01603_),
    .Q(\mem[39][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12911_ (.CLK(clknet_leaf_288_i_clk),
    .D(_01604_),
    .Q(\mem[39][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12912_ (.CLK(clknet_leaf_288_i_clk),
    .D(_01605_),
    .Q(\mem[39][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12913_ (.CLK(clknet_leaf_26_i_clk),
    .D(_01606_),
    .Q(\mem[39][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12914_ (.CLK(clknet_leaf_1_i_clk),
    .D(_01607_),
    .Q(\mem[39][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12915_ (.CLK(clknet_leaf_286_i_clk),
    .D(_01608_),
    .Q(\mem[39][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12916_ (.CLK(clknet_leaf_6_i_clk),
    .D(_01609_),
    .Q(\mem[39][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12917_ (.CLK(clknet_leaf_12_i_clk),
    .D(_01610_),
    .Q(\mem[39][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12918_ (.CLK(clknet_leaf_26_i_clk),
    .D(_01611_),
    .Q(\mem[39][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12919_ (.CLK(clknet_leaf_27_i_clk),
    .D(_01612_),
    .Q(\mem[39][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12920_ (.CLK(clknet_leaf_26_i_clk),
    .D(_01613_),
    .Q(\mem[39][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12921_ (.CLK(clknet_leaf_25_i_clk),
    .D(_01614_),
    .Q(\mem[39][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12922_ (.CLK(clknet_leaf_9_i_clk),
    .D(_01615_),
    .Q(\mem[39][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12923_ (.CLK(clknet_leaf_8_i_clk),
    .D(_01616_),
    .Q(\mem[39][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12924_ (.CLK(clknet_leaf_240_i_clk),
    .D(_01617_),
    .Q(\mem[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12925_ (.CLK(clknet_leaf_247_i_clk),
    .D(_01618_),
    .Q(\mem[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12926_ (.CLK(clknet_leaf_237_i_clk),
    .D(_01619_),
    .Q(\mem[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12927_ (.CLK(clknet_leaf_240_i_clk),
    .D(_01620_),
    .Q(\mem[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12928_ (.CLK(clknet_leaf_238_i_clk),
    .D(_01621_),
    .Q(\mem[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12929_ (.CLK(clknet_leaf_248_i_clk),
    .D(_01622_),
    .Q(\mem[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12930_ (.CLK(clknet_leaf_238_i_clk),
    .D(_01623_),
    .Q(\mem[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12931_ (.CLK(clknet_leaf_236_i_clk),
    .D(_01624_),
    .Q(\mem[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12932_ (.CLK(clknet_leaf_236_i_clk),
    .D(_01625_),
    .Q(\mem[29][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12933_ (.CLK(clknet_leaf_237_i_clk),
    .D(_01626_),
    .Q(\mem[29][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12934_ (.CLK(clknet_leaf_242_i_clk),
    .D(_01627_),
    .Q(\mem[29][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12935_ (.CLK(clknet_leaf_242_i_clk),
    .D(_01628_),
    .Q(\mem[29][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12936_ (.CLK(clknet_leaf_242_i_clk),
    .D(_01629_),
    .Q(\mem[29][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12937_ (.CLK(clknet_leaf_250_i_clk),
    .D(_01630_),
    .Q(\mem[29][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12938_ (.CLK(clknet_leaf_242_i_clk),
    .D(_01631_),
    .Q(\mem[29][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12939_ (.CLK(clknet_leaf_228_i_clk),
    .D(_01632_),
    .Q(\mem[29][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12940_ (.CLK(clknet_leaf_286_i_clk),
    .D(_01633_),
    .Q(\mem[99][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12941_ (.CLK(clknet_leaf_261_i_clk),
    .D(_01634_),
    .Q(\mem[99][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12942_ (.CLK(clknet_leaf_286_i_clk),
    .D(_01635_),
    .Q(\mem[99][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12943_ (.CLK(clknet_leaf_284_i_clk),
    .D(_01636_),
    .Q(\mem[99][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12944_ (.CLK(clknet_leaf_277_i_clk),
    .D(_01637_),
    .Q(\mem[99][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12945_ (.CLK(clknet_leaf_259_i_clk),
    .D(_01638_),
    .Q(\mem[99][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12946_ (.CLK(clknet_leaf_261_i_clk),
    .D(_01639_),
    .Q(\mem[99][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12947_ (.CLK(clknet_leaf_284_i_clk),
    .D(_01640_),
    .Q(\mem[99][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12948_ (.CLK(clknet_leaf_275_i_clk),
    .D(_01641_),
    .Q(\mem[99][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12949_ (.CLK(clknet_leaf_276_i_clk),
    .D(_01642_),
    .Q(\mem[99][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12950_ (.CLK(clknet_leaf_7_i_clk),
    .D(_01643_),
    .Q(\mem[99][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12951_ (.CLK(clknet_leaf_27_i_clk),
    .D(_01644_),
    .Q(\mem[99][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12952_ (.CLK(clknet_leaf_280_i_clk),
    .D(_01645_),
    .Q(\mem[99][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12953_ (.CLK(clknet_leaf_30_i_clk),
    .D(_01646_),
    .Q(\mem[99][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12954_ (.CLK(clknet_leaf_7_i_clk),
    .D(_01647_),
    .Q(\mem[99][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12955_ (.CLK(clknet_leaf_28_i_clk),
    .D(_01648_),
    .Q(\mem[99][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12956_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01649_),
    .Q(\mem[109][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12957_ (.CLK(clknet_leaf_110_i_clk),
    .D(_01650_),
    .Q(\mem[109][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12958_ (.CLK(clknet_leaf_51_i_clk),
    .D(_01651_),
    .Q(\mem[109][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12959_ (.CLK(clknet_leaf_51_i_clk),
    .D(_01652_),
    .Q(\mem[109][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12960_ (.CLK(clknet_leaf_52_i_clk),
    .D(_01653_),
    .Q(\mem[109][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12961_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01654_),
    .Q(\mem[109][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12962_ (.CLK(clknet_leaf_52_i_clk),
    .D(_01655_),
    .Q(\mem[109][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12963_ (.CLK(clknet_leaf_44_i_clk),
    .D(_01656_),
    .Q(\mem[109][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12964_ (.CLK(clknet_leaf_45_i_clk),
    .D(_01657_),
    .Q(\mem[109][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12965_ (.CLK(clknet_leaf_51_i_clk),
    .D(_01658_),
    .Q(\mem[109][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12966_ (.CLK(clknet_leaf_47_i_clk),
    .D(_01659_),
    .Q(\mem[109][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12967_ (.CLK(clknet_leaf_45_i_clk),
    .D(_01660_),
    .Q(\mem[109][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12968_ (.CLK(clknet_leaf_47_i_clk),
    .D(_01661_),
    .Q(\mem[109][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12969_ (.CLK(clknet_leaf_106_i_clk),
    .D(_01662_),
    .Q(\mem[109][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12970_ (.CLK(clknet_leaf_106_i_clk),
    .D(_01663_),
    .Q(\mem[109][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12971_ (.CLK(clknet_leaf_47_i_clk),
    .D(_01664_),
    .Q(\mem[109][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12972_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01665_),
    .Q(\mem[119][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12973_ (.CLK(clknet_leaf_102_i_clk),
    .D(_01666_),
    .Q(\mem[119][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12974_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01667_),
    .Q(\mem[119][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12975_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01668_),
    .Q(\mem[119][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12976_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01669_),
    .Q(\mem[119][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12977_ (.CLK(clknet_leaf_102_i_clk),
    .D(_01670_),
    .Q(\mem[119][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12978_ (.CLK(clknet_leaf_100_i_clk),
    .D(_01671_),
    .Q(\mem[119][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12979_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01672_),
    .Q(\mem[119][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12980_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01673_),
    .Q(\mem[119][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12981_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01674_),
    .Q(\mem[119][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12982_ (.CLK(clknet_leaf_145_i_clk),
    .D(_01675_),
    .Q(\mem[119][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12983_ (.CLK(clknet_leaf_137_i_clk),
    .D(_01676_),
    .Q(\mem[119][11] ));
 sky130_fd_sc_hd__dfxtp_1 _12984_ (.CLK(clknet_leaf_146_i_clk),
    .D(_01677_),
    .Q(\mem[119][12] ));
 sky130_fd_sc_hd__dfxtp_1 _12985_ (.CLK(clknet_leaf_123_i_clk),
    .D(_01678_),
    .Q(\mem[119][13] ));
 sky130_fd_sc_hd__dfxtp_1 _12986_ (.CLK(clknet_leaf_147_i_clk),
    .D(_01679_),
    .Q(\mem[119][14] ));
 sky130_fd_sc_hd__dfxtp_1 _12987_ (.CLK(clknet_leaf_146_i_clk),
    .D(_01680_),
    .Q(\mem[119][15] ));
 sky130_fd_sc_hd__dfxtp_1 _12988_ (.CLK(clknet_leaf_100_i_clk),
    .D(_01681_),
    .Q(\mem[127][0] ));
 sky130_fd_sc_hd__dfxtp_1 _12989_ (.CLK(clknet_leaf_100_i_clk),
    .D(_01682_),
    .Q(\mem[127][1] ));
 sky130_fd_sc_hd__dfxtp_1 _12990_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01683_),
    .Q(\mem[127][2] ));
 sky130_fd_sc_hd__dfxtp_1 _12991_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01684_),
    .Q(\mem[127][3] ));
 sky130_fd_sc_hd__dfxtp_1 _12992_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01685_),
    .Q(\mem[127][4] ));
 sky130_fd_sc_hd__dfxtp_1 _12993_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01686_),
    .Q(\mem[127][5] ));
 sky130_fd_sc_hd__dfxtp_1 _12994_ (.CLK(clknet_leaf_127_i_clk),
    .D(_01687_),
    .Q(\mem[127][6] ));
 sky130_fd_sc_hd__dfxtp_1 _12995_ (.CLK(clknet_leaf_127_i_clk),
    .D(_01688_),
    .Q(\mem[127][7] ));
 sky130_fd_sc_hd__dfxtp_1 _12996_ (.CLK(clknet_leaf_128_i_clk),
    .D(_01689_),
    .Q(\mem[127][8] ));
 sky130_fd_sc_hd__dfxtp_1 _12997_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01690_),
    .Q(\mem[127][9] ));
 sky130_fd_sc_hd__dfxtp_1 _12998_ (.CLK(clknet_leaf_144_i_clk),
    .D(_01691_),
    .Q(\mem[127][10] ));
 sky130_fd_sc_hd__dfxtp_1 _12999_ (.CLK(clknet_leaf_136_i_clk),
    .D(_01692_),
    .Q(\mem[127][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13000_ (.CLK(clknet_leaf_143_i_clk),
    .D(_01693_),
    .Q(\mem[127][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13001_ (.CLK(clknet_leaf_124_i_clk),
    .D(_01694_),
    .Q(\mem[127][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13002_ (.CLK(clknet_leaf_144_i_clk),
    .D(_01695_),
    .Q(\mem[127][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13003_ (.CLK(clknet_leaf_136_i_clk),
    .D(_01696_),
    .Q(\mem[127][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13004_ (.CLK(clknet_leaf_112_i_clk),
    .D(_01697_),
    .Q(\mem[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13005_ (.CLK(clknet_leaf_110_i_clk),
    .D(_01698_),
    .Q(\mem[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13006_ (.CLK(clknet_leaf_108_i_clk),
    .D(_01699_),
    .Q(\mem[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13007_ (.CLK(clknet_leaf_108_i_clk),
    .D(_01700_),
    .Q(\mem[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13008_ (.CLK(clknet_leaf_107_i_clk),
    .D(_01701_),
    .Q(\mem[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13009_ (.CLK(clknet_leaf_111_i_clk),
    .D(_01702_),
    .Q(\mem[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13010_ (.CLK(clknet_leaf_107_i_clk),
    .D(_01703_),
    .Q(\mem[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13011_ (.CLK(clknet_leaf_108_i_clk),
    .D(_01704_),
    .Q(\mem[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13012_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01705_),
    .Q(\mem[12][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13013_ (.CLK(clknet_leaf_110_i_clk),
    .D(_01706_),
    .Q(\mem[12][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13014_ (.CLK(clknet_leaf_113_i_clk),
    .D(_01707_),
    .Q(\mem[12][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13015_ (.CLK(clknet_leaf_179_i_clk),
    .D(_01708_),
    .Q(\mem[12][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13016_ (.CLK(clknet_leaf_179_i_clk),
    .D(_01709_),
    .Q(\mem[12][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13017_ (.CLK(clknet_leaf_111_i_clk),
    .D(_01710_),
    .Q(\mem[12][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13018_ (.CLK(clknet_leaf_179_i_clk),
    .D(_01711_),
    .Q(\mem[12][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13019_ (.CLK(clknet_leaf_179_i_clk),
    .D(_01712_),
    .Q(\mem[12][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13020_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01713_),
    .Q(\mem[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13021_ (.CLK(clknet_leaf_110_i_clk),
    .D(_01714_),
    .Q(\mem[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13022_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01715_),
    .Q(\mem[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13023_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01716_),
    .Q(\mem[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13024_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01717_),
    .Q(\mem[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13025_ (.CLK(clknet_leaf_111_i_clk),
    .D(_01718_),
    .Q(\mem[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13026_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01719_),
    .Q(\mem[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13027_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01720_),
    .Q(\mem[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13028_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01721_),
    .Q(\mem[13][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13029_ (.CLK(clknet_leaf_112_i_clk),
    .D(_01722_),
    .Q(\mem[13][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13030_ (.CLK(clknet_leaf_180_i_clk),
    .D(_01723_),
    .Q(\mem[13][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13031_ (.CLK(clknet_leaf_180_i_clk),
    .D(_01724_),
    .Q(\mem[13][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13032_ (.CLK(clknet_leaf_180_i_clk),
    .D(_01725_),
    .Q(\mem[13][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13033_ (.CLK(clknet_leaf_112_i_clk),
    .D(_01726_),
    .Q(\mem[13][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13034_ (.CLK(clknet_leaf_178_i_clk),
    .D(_01727_),
    .Q(\mem[13][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13035_ (.CLK(clknet_leaf_178_i_clk),
    .D(_01728_),
    .Q(\mem[13][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13036_ (.CLK(clknet_leaf_180_i_clk),
    .D(_01729_),
    .Q(\mem[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13037_ (.CLK(clknet_leaf_109_i_clk),
    .D(_01730_),
    .Q(\mem[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13038_ (.CLK(clknet_leaf_109_i_clk),
    .D(_01731_),
    .Q(\mem[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13039_ (.CLK(clknet_leaf_108_i_clk),
    .D(_01732_),
    .Q(\mem[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13040_ (.CLK(clknet_leaf_108_i_clk),
    .D(_01733_),
    .Q(\mem[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13041_ (.CLK(clknet_leaf_109_i_clk),
    .D(_01734_),
    .Q(\mem[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13042_ (.CLK(clknet_leaf_109_i_clk),
    .D(_01735_),
    .Q(\mem[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13043_ (.CLK(clknet_leaf_108_i_clk),
    .D(_01736_),
    .Q(\mem[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13044_ (.CLK(clknet_leaf_39_i_clk),
    .D(_01737_),
    .Q(\mem[14][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13045_ (.CLK(clknet_leaf_112_i_clk),
    .D(_01738_),
    .Q(\mem[14][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13046_ (.CLK(clknet_leaf_113_i_clk),
    .D(_01739_),
    .Q(\mem[14][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13047_ (.CLK(clknet_leaf_180_i_clk),
    .D(_01740_),
    .Q(\mem[14][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13048_ (.CLK(clknet_leaf_178_i_clk),
    .D(_01741_),
    .Q(\mem[14][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13049_ (.CLK(clknet_leaf_113_i_clk),
    .D(_01742_),
    .Q(\mem[14][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13050_ (.CLK(clknet_leaf_178_i_clk),
    .D(_01743_),
    .Q(\mem[14][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13051_ (.CLK(clknet_leaf_178_i_clk),
    .D(_01744_),
    .Q(\mem[14][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13052_ (.CLK(clknet_leaf_113_i_clk),
    .D(_01745_),
    .Q(\mem[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13053_ (.CLK(clknet_leaf_111_i_clk),
    .D(_01746_),
    .Q(\mem[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13054_ (.CLK(clknet_leaf_108_i_clk),
    .D(_01747_),
    .Q(\mem[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13055_ (.CLK(clknet_leaf_108_i_clk),
    .D(_01748_),
    .Q(\mem[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13056_ (.CLK(clknet_leaf_109_i_clk),
    .D(_01749_),
    .Q(\mem[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13057_ (.CLK(clknet_leaf_109_i_clk),
    .D(_01750_),
    .Q(\mem[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13058_ (.CLK(clknet_leaf_110_i_clk),
    .D(_01751_),
    .Q(\mem[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13059_ (.CLK(clknet_leaf_108_i_clk),
    .D(_01752_),
    .Q(\mem[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13060_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01753_),
    .Q(\mem[15][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13061_ (.CLK(clknet_leaf_111_i_clk),
    .D(_01754_),
    .Q(\mem[15][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13062_ (.CLK(clknet_leaf_113_i_clk),
    .D(_01755_),
    .Q(\mem[15][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13063_ (.CLK(clknet_leaf_180_i_clk),
    .D(_01756_),
    .Q(\mem[15][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13064_ (.CLK(clknet_leaf_179_i_clk),
    .D(_01757_),
    .Q(\mem[15][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13065_ (.CLK(clknet_leaf_114_i_clk),
    .D(_01758_),
    .Q(\mem[15][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13066_ (.CLK(clknet_leaf_178_i_clk),
    .D(_01759_),
    .Q(\mem[15][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13067_ (.CLK(clknet_leaf_178_i_clk),
    .D(_01760_),
    .Q(\mem[15][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13068_ (.CLK(clknet_leaf_242_i_clk),
    .D(_01761_),
    .Q(\mem[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13069_ (.CLK(clknet_leaf_249_i_clk),
    .D(_01762_),
    .Q(\mem[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13070_ (.CLK(clknet_leaf_239_i_clk),
    .D(_01763_),
    .Q(\mem[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13071_ (.CLK(clknet_leaf_239_i_clk),
    .D(_01764_),
    .Q(\mem[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13072_ (.CLK(clknet_leaf_238_i_clk),
    .D(_01765_),
    .Q(\mem[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13073_ (.CLK(clknet_leaf_248_i_clk),
    .D(_01766_),
    .Q(\mem[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13074_ (.CLK(clknet_leaf_238_i_clk),
    .D(_01767_),
    .Q(\mem[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13075_ (.CLK(clknet_leaf_236_i_clk),
    .D(_01768_),
    .Q(\mem[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13076_ (.CLK(clknet_leaf_236_i_clk),
    .D(_01769_),
    .Q(\mem[16][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13077_ (.CLK(clknet_leaf_237_i_clk),
    .D(_01770_),
    .Q(\mem[16][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13078_ (.CLK(clknet_leaf_241_i_clk),
    .D(_01771_),
    .Q(\mem[16][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13079_ (.CLK(clknet_leaf_229_i_clk),
    .D(_01772_),
    .Q(\mem[16][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13080_ (.CLK(clknet_leaf_229_i_clk),
    .D(_01773_),
    .Q(\mem[16][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13081_ (.CLK(clknet_leaf_244_i_clk),
    .D(_01774_),
    .Q(\mem[16][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13082_ (.CLK(clknet_leaf_228_i_clk),
    .D(_01775_),
    .Q(\mem[16][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13083_ (.CLK(clknet_leaf_228_i_clk),
    .D(_01776_),
    .Q(\mem[16][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13084_ (.CLK(clknet_leaf_242_i_clk),
    .D(_01777_),
    .Q(\mem[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13085_ (.CLK(clknet_leaf_257_i_clk),
    .D(_01778_),
    .Q(\mem[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13086_ (.CLK(clknet_leaf_239_i_clk),
    .D(_01779_),
    .Q(\mem[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13087_ (.CLK(clknet_leaf_266_i_clk),
    .D(_01780_),
    .Q(\mem[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13088_ (.CLK(clknet_leaf_267_i_clk),
    .D(_01781_),
    .Q(\mem[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13089_ (.CLK(clknet_leaf_256_i_clk),
    .D(_01782_),
    .Q(\mem[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13090_ (.CLK(clknet_leaf_267_i_clk),
    .D(_01783_),
    .Q(\mem[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13091_ (.CLK(clknet_leaf_267_i_clk),
    .D(_01784_),
    .Q(\mem[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13092_ (.CLK(clknet_leaf_267_i_clk),
    .D(_01785_),
    .Q(\mem[17][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13093_ (.CLK(clknet_leaf_237_i_clk),
    .D(_01786_),
    .Q(\mem[17][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13094_ (.CLK(clknet_leaf_241_i_clk),
    .D(_01787_),
    .Q(\mem[17][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13095_ (.CLK(clknet_leaf_241_i_clk),
    .D(_01788_),
    .Q(\mem[17][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13096_ (.CLK(clknet_leaf_229_i_clk),
    .D(_01789_),
    .Q(\mem[17][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13097_ (.CLK(clknet_leaf_246_i_clk),
    .D(_01790_),
    .Q(\mem[17][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13098_ (.CLK(clknet_leaf_228_i_clk),
    .D(_01791_),
    .Q(\mem[17][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13099_ (.CLK(clknet_leaf_230_i_clk),
    .D(_01792_),
    .Q(\mem[17][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13100_ (.CLK(clknet_leaf_240_i_clk),
    .D(_01793_),
    .Q(\mem[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13101_ (.CLK(clknet_leaf_249_i_clk),
    .D(_01794_),
    .Q(\mem[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13102_ (.CLK(clknet_leaf_239_i_clk),
    .D(_01795_),
    .Q(\mem[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13103_ (.CLK(clknet_leaf_265_i_clk),
    .D(_01796_),
    .Q(\mem[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13104_ (.CLK(clknet_leaf_268_i_clk),
    .D(_01797_),
    .Q(\mem[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13105_ (.CLK(clknet_leaf_257_i_clk),
    .D(_01798_),
    .Q(\mem[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13106_ (.CLK(clknet_leaf_268_i_clk),
    .D(_01799_),
    .Q(\mem[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13107_ (.CLK(clknet_leaf_268_i_clk),
    .D(_01800_),
    .Q(\mem[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13108_ (.CLK(clknet_leaf_268_i_clk),
    .D(_01801_),
    .Q(\mem[18][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13109_ (.CLK(clknet_leaf_237_i_clk),
    .D(_01802_),
    .Q(\mem[18][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13110_ (.CLK(clknet_leaf_240_i_clk),
    .D(_01803_),
    .Q(\mem[18][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13111_ (.CLK(clknet_leaf_241_i_clk),
    .D(_01804_),
    .Q(\mem[18][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13112_ (.CLK(clknet_leaf_228_i_clk),
    .D(_01805_),
    .Q(\mem[18][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13113_ (.CLK(clknet_leaf_245_i_clk),
    .D(_01806_),
    .Q(\mem[18][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13114_ (.CLK(clknet_leaf_228_i_clk),
    .D(_01807_),
    .Q(\mem[18][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13115_ (.CLK(clknet_leaf_228_i_clk),
    .D(_01808_),
    .Q(\mem[18][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13116_ (.CLK(clknet_leaf_251_i_clk),
    .D(_01809_),
    .Q(\mem[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13117_ (.CLK(clknet_leaf_252_i_clk),
    .D(_01810_),
    .Q(\mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13118_ (.CLK(clknet_leaf_249_i_clk),
    .D(_01811_),
    .Q(\mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13119_ (.CLK(clknet_leaf_259_i_clk),
    .D(_01812_),
    .Q(\mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13120_ (.CLK(clknet_leaf_255_i_clk),
    .D(_01813_),
    .Q(\mem[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13121_ (.CLK(clknet_leaf_254_i_clk),
    .D(_01814_),
    .Q(\mem[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13122_ (.CLK(clknet_leaf_259_i_clk),
    .D(_01815_),
    .Q(\mem[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13123_ (.CLK(clknet_leaf_255_i_clk),
    .D(_01816_),
    .Q(\mem[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13124_ (.CLK(clknet_leaf_254_i_clk),
    .D(_01817_),
    .Q(\mem[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13125_ (.CLK(clknet_leaf_254_i_clk),
    .D(_01818_),
    .Q(\mem[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13126_ (.CLK(clknet_leaf_251_i_clk),
    .D(_01819_),
    .Q(\mem[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13127_ (.CLK(clknet_leaf_250_i_clk),
    .D(_01820_),
    .Q(\mem[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13128_ (.CLK(clknet_leaf_250_i_clk),
    .D(_01821_),
    .Q(\mem[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13129_ (.CLK(clknet_leaf_251_i_clk),
    .D(_01822_),
    .Q(\mem[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13130_ (.CLK(clknet_leaf_183_i_clk),
    .D(_01823_),
    .Q(\mem[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13131_ (.CLK(clknet_leaf_183_i_clk),
    .D(_01824_),
    .Q(\mem[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13132_ (.CLK(clknet_leaf_266_i_clk),
    .D(_01825_),
    .Q(\mem[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13133_ (.CLK(clknet_leaf_266_i_clk),
    .D(_01826_),
    .Q(\mem[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13134_ (.CLK(clknet_leaf_263_i_clk),
    .D(_01827_),
    .Q(\mem[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13135_ (.CLK(clknet_leaf_263_i_clk),
    .D(_01828_),
    .Q(\mem[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13136_ (.CLK(clknet_leaf_273_i_clk),
    .D(_01829_),
    .Q(\mem[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13137_ (.CLK(clknet_leaf_265_i_clk),
    .D(_01830_),
    .Q(\mem[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13138_ (.CLK(clknet_leaf_273_i_clk),
    .D(_01831_),
    .Q(\mem[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13139_ (.CLK(clknet_leaf_274_i_clk),
    .D(_01832_),
    .Q(\mem[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13140_ (.CLK(clknet_leaf_274_i_clk),
    .D(_01833_),
    .Q(\mem[20][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13141_ (.CLK(clknet_leaf_271_i_clk),
    .D(_01834_),
    .Q(\mem[20][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13142_ (.CLK(clknet_leaf_235_i_clk),
    .D(_01835_),
    .Q(\mem[20][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13143_ (.CLK(clknet_leaf_235_i_clk),
    .D(_01836_),
    .Q(\mem[20][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13144_ (.CLK(clknet_leaf_234_i_clk),
    .D(_01837_),
    .Q(\mem[20][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13145_ (.CLK(clknet_leaf_249_i_clk),
    .D(_01838_),
    .Q(\mem[20][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13146_ (.CLK(clknet_leaf_234_i_clk),
    .D(_01839_),
    .Q(\mem[20][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13147_ (.CLK(clknet_leaf_232_i_clk),
    .D(_01840_),
    .Q(\mem[20][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13148_ (.CLK(clknet_leaf_266_i_clk),
    .D(_01841_),
    .Q(\mem[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13149_ (.CLK(clknet_leaf_248_i_clk),
    .D(_01842_),
    .Q(\mem[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13150_ (.CLK(clknet_leaf_264_i_clk),
    .D(_01843_),
    .Q(\mem[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13151_ (.CLK(clknet_leaf_265_i_clk),
    .D(_01844_),
    .Q(\mem[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13152_ (.CLK(clknet_leaf_269_i_clk),
    .D(_01845_),
    .Q(\mem[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13153_ (.CLK(clknet_leaf_257_i_clk),
    .D(_01846_),
    .Q(\mem[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13154_ (.CLK(clknet_leaf_270_i_clk),
    .D(_01847_),
    .Q(\mem[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13155_ (.CLK(clknet_leaf_272_i_clk),
    .D(_01848_),
    .Q(\mem[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13156_ (.CLK(clknet_leaf_271_i_clk),
    .D(_01849_),
    .Q(\mem[21][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13157_ (.CLK(clknet_leaf_271_i_clk),
    .D(_01850_),
    .Q(\mem[21][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13158_ (.CLK(clknet_leaf_235_i_clk),
    .D(_01851_),
    .Q(\mem[21][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13159_ (.CLK(clknet_leaf_235_i_clk),
    .D(_01852_),
    .Q(\mem[21][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13160_ (.CLK(clknet_leaf_234_i_clk),
    .D(_01853_),
    .Q(\mem[21][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13161_ (.CLK(clknet_leaf_249_i_clk),
    .D(_01854_),
    .Q(\mem[21][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13162_ (.CLK(clknet_leaf_234_i_clk),
    .D(_01855_),
    .Q(\mem[21][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13163_ (.CLK(clknet_leaf_232_i_clk),
    .D(_01856_),
    .Q(\mem[21][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13164_ (.CLK(clknet_leaf_266_i_clk),
    .D(_01857_),
    .Q(\mem[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13165_ (.CLK(clknet_leaf_266_i_clk),
    .D(_01858_),
    .Q(\mem[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13166_ (.CLK(clknet_leaf_264_i_clk),
    .D(_01859_),
    .Q(\mem[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13167_ (.CLK(clknet_leaf_265_i_clk),
    .D(_01860_),
    .Q(\mem[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13168_ (.CLK(clknet_leaf_273_i_clk),
    .D(_01861_),
    .Q(\mem[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13169_ (.CLK(clknet_leaf_265_i_clk),
    .D(_01862_),
    .Q(\mem[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13170_ (.CLK(clknet_leaf_273_i_clk),
    .D(_01863_),
    .Q(\mem[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13171_ (.CLK(clknet_leaf_272_i_clk),
    .D(_01864_),
    .Q(\mem[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13172_ (.CLK(clknet_leaf_272_i_clk),
    .D(_01865_),
    .Q(\mem[22][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13173_ (.CLK(clknet_leaf_271_i_clk),
    .D(_01866_),
    .Q(\mem[22][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13174_ (.CLK(clknet_leaf_235_i_clk),
    .D(_01867_),
    .Q(\mem[22][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13175_ (.CLK(clknet_leaf_235_i_clk),
    .D(_01868_),
    .Q(\mem[22][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13176_ (.CLK(clknet_leaf_234_i_clk),
    .D(_01869_),
    .Q(\mem[22][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13177_ (.CLK(clknet_leaf_249_i_clk),
    .D(_01870_),
    .Q(\mem[22][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13178_ (.CLK(clknet_leaf_234_i_clk),
    .D(_01871_),
    .Q(\mem[22][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13179_ (.CLK(clknet_leaf_232_i_clk),
    .D(_01872_),
    .Q(\mem[22][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13180_ (.CLK(clknet_leaf_265_i_clk),
    .D(_01873_),
    .Q(\mem[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13181_ (.CLK(clknet_leaf_258_i_clk),
    .D(_01874_),
    .Q(\mem[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13182_ (.CLK(clknet_leaf_263_i_clk),
    .D(_01875_),
    .Q(\mem[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13183_ (.CLK(clknet_leaf_265_i_clk),
    .D(_01876_),
    .Q(\mem[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13184_ (.CLK(clknet_leaf_278_i_clk),
    .D(_01877_),
    .Q(\mem[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13185_ (.CLK(clknet_leaf_258_i_clk),
    .D(_01878_),
    .Q(\mem[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13186_ (.CLK(clknet_leaf_273_i_clk),
    .D(_01879_),
    .Q(\mem[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13187_ (.CLK(clknet_leaf_273_i_clk),
    .D(_01880_),
    .Q(\mem[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13188_ (.CLK(clknet_leaf_272_i_clk),
    .D(_01881_),
    .Q(\mem[23][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13189_ (.CLK(clknet_leaf_271_i_clk),
    .D(_01882_),
    .Q(\mem[23][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13190_ (.CLK(clknet_leaf_235_i_clk),
    .D(_01883_),
    .Q(\mem[23][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13191_ (.CLK(clknet_leaf_235_i_clk),
    .D(_01884_),
    .Q(\mem[23][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13192_ (.CLK(clknet_leaf_234_i_clk),
    .D(_01885_),
    .Q(\mem[23][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13193_ (.CLK(clknet_leaf_249_i_clk),
    .D(_01886_),
    .Q(\mem[23][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13194_ (.CLK(clknet_leaf_234_i_clk),
    .D(_01887_),
    .Q(\mem[23][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13195_ (.CLK(clknet_leaf_232_i_clk),
    .D(_01888_),
    .Q(\mem[23][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13196_ (.CLK(clknet_leaf_247_i_clk),
    .D(_01889_),
    .Q(\mem[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13197_ (.CLK(clknet_leaf_248_i_clk),
    .D(_01890_),
    .Q(\mem[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13198_ (.CLK(clknet_leaf_268_i_clk),
    .D(_01891_),
    .Q(\mem[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13199_ (.CLK(clknet_leaf_268_i_clk),
    .D(_01892_),
    .Q(\mem[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13200_ (.CLK(clknet_leaf_273_i_clk),
    .D(_01893_),
    .Q(\mem[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13201_ (.CLK(clknet_leaf_248_i_clk),
    .D(_01894_),
    .Q(\mem[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13202_ (.CLK(clknet_leaf_272_i_clk),
    .D(_01895_),
    .Q(\mem[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13203_ (.CLK(clknet_leaf_272_i_clk),
    .D(_01896_),
    .Q(\mem[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13204_ (.CLK(clknet_leaf_272_i_clk),
    .D(_01897_),
    .Q(\mem[24][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13205_ (.CLK(clknet_leaf_271_i_clk),
    .D(_01898_),
    .Q(\mem[24][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13206_ (.CLK(clknet_leaf_231_i_clk),
    .D(_01899_),
    .Q(\mem[24][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13207_ (.CLK(clknet_leaf_232_i_clk),
    .D(_01900_),
    .Q(\mem[24][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13208_ (.CLK(clknet_leaf_231_i_clk),
    .D(_01901_),
    .Q(\mem[24][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13209_ (.CLK(clknet_leaf_246_i_clk),
    .D(_01902_),
    .Q(\mem[24][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13210_ (.CLK(clknet_leaf_223_i_clk),
    .D(_01903_),
    .Q(\mem[24][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13211_ (.CLK(clknet_leaf_223_i_clk),
    .D(_01904_),
    .Q(\mem[24][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13212_ (.CLK(clknet_leaf_247_i_clk),
    .D(_01905_),
    .Q(\mem[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13213_ (.CLK(clknet_leaf_258_i_clk),
    .D(_01906_),
    .Q(\mem[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13214_ (.CLK(clknet_leaf_278_i_clk),
    .D(_01907_),
    .Q(\mem[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13215_ (.CLK(clknet_leaf_264_i_clk),
    .D(_01908_),
    .Q(\mem[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13216_ (.CLK(clknet_leaf_278_i_clk),
    .D(_01909_),
    .Q(\mem[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13217_ (.CLK(clknet_leaf_258_i_clk),
    .D(_01910_),
    .Q(\mem[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13218_ (.CLK(clknet_leaf_273_i_clk),
    .D(_01911_),
    .Q(\mem[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13219_ (.CLK(clknet_leaf_274_i_clk),
    .D(_01912_),
    .Q(\mem[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13220_ (.CLK(clknet_leaf_274_i_clk),
    .D(_01913_),
    .Q(\mem[25][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13221_ (.CLK(clknet_leaf_271_i_clk),
    .D(_01914_),
    .Q(\mem[25][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13222_ (.CLK(clknet_leaf_231_i_clk),
    .D(_01915_),
    .Q(\mem[25][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13223_ (.CLK(clknet_leaf_232_i_clk),
    .D(_01916_),
    .Q(\mem[25][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13224_ (.CLK(clknet_leaf_231_i_clk),
    .D(_01917_),
    .Q(\mem[25][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13225_ (.CLK(clknet_leaf_250_i_clk),
    .D(_01918_),
    .Q(\mem[25][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13226_ (.CLK(clknet_leaf_223_i_clk),
    .D(_01919_),
    .Q(\mem[25][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13227_ (.CLK(clknet_leaf_223_i_clk),
    .D(_01920_),
    .Q(\mem[25][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13228_ (.CLK(clknet_leaf_247_i_clk),
    .D(_01921_),
    .Q(\mem[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13229_ (.CLK(clknet_leaf_258_i_clk),
    .D(_01922_),
    .Q(\mem[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13230_ (.CLK(clknet_leaf_264_i_clk),
    .D(_01923_),
    .Q(\mem[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13231_ (.CLK(clknet_leaf_269_i_clk),
    .D(_01924_),
    .Q(\mem[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13232_ (.CLK(clknet_leaf_273_i_clk),
    .D(_01925_),
    .Q(\mem[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13233_ (.CLK(clknet_leaf_258_i_clk),
    .D(_01926_),
    .Q(\mem[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13234_ (.CLK(clknet_leaf_272_i_clk),
    .D(_01927_),
    .Q(\mem[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13235_ (.CLK(clknet_leaf_272_i_clk),
    .D(_01928_),
    .Q(\mem[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13236_ (.CLK(clknet_leaf_274_i_clk),
    .D(_01929_),
    .Q(\mem[26][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13237_ (.CLK(clknet_leaf_271_i_clk),
    .D(_01930_),
    .Q(\mem[26][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13238_ (.CLK(clknet_leaf_231_i_clk),
    .D(_01931_),
    .Q(\mem[26][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13239_ (.CLK(clknet_leaf_232_i_clk),
    .D(_01932_),
    .Q(\mem[26][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13240_ (.CLK(clknet_leaf_231_i_clk),
    .D(_01933_),
    .Q(\mem[26][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13241_ (.CLK(clknet_leaf_245_i_clk),
    .D(_01934_),
    .Q(\mem[26][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13242_ (.CLK(clknet_leaf_223_i_clk),
    .D(_01935_),
    .Q(\mem[26][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13243_ (.CLK(clknet_leaf_223_i_clk),
    .D(_01936_),
    .Q(\mem[26][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13244_ (.CLK(clknet_leaf_247_i_clk),
    .D(_01937_),
    .Q(\mem[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13245_ (.CLK(clknet_leaf_258_i_clk),
    .D(_01938_),
    .Q(\mem[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13246_ (.CLK(clknet_leaf_278_i_clk),
    .D(_01939_),
    .Q(\mem[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13247_ (.CLK(clknet_leaf_278_i_clk),
    .D(_01940_),
    .Q(\mem[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13248_ (.CLK(clknet_leaf_278_i_clk),
    .D(_01941_),
    .Q(\mem[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13249_ (.CLK(clknet_leaf_258_i_clk),
    .D(_01942_),
    .Q(\mem[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13250_ (.CLK(clknet_leaf_273_i_clk),
    .D(_01943_),
    .Q(\mem[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13251_ (.CLK(clknet_leaf_274_i_clk),
    .D(_01944_),
    .Q(\mem[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13252_ (.CLK(clknet_leaf_274_i_clk),
    .D(_01945_),
    .Q(\mem[27][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13253_ (.CLK(clknet_leaf_272_i_clk),
    .D(_01946_),
    .Q(\mem[27][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13254_ (.CLK(clknet_leaf_231_i_clk),
    .D(_01947_),
    .Q(\mem[27][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13255_ (.CLK(clknet_leaf_232_i_clk),
    .D(_01948_),
    .Q(\mem[27][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13256_ (.CLK(clknet_leaf_231_i_clk),
    .D(_01949_),
    .Q(\mem[27][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13257_ (.CLK(clknet_leaf_250_i_clk),
    .D(_01950_),
    .Q(\mem[27][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13258_ (.CLK(clknet_leaf_231_i_clk),
    .D(_01951_),
    .Q(\mem[27][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13259_ (.CLK(clknet_leaf_231_i_clk),
    .D(_01952_),
    .Q(\mem[27][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13260_ (.CLK(clknet_leaf_239_i_clk),
    .D(_01953_),
    .Q(\mem[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13261_ (.CLK(clknet_leaf_248_i_clk),
    .D(_01954_),
    .Q(\mem[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13262_ (.CLK(clknet_leaf_238_i_clk),
    .D(_01955_),
    .Q(\mem[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13263_ (.CLK(clknet_leaf_268_i_clk),
    .D(_01956_),
    .Q(\mem[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13264_ (.CLK(clknet_leaf_270_i_clk),
    .D(_01957_),
    .Q(\mem[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13265_ (.CLK(clknet_leaf_239_i_clk),
    .D(_01958_),
    .Q(\mem[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13266_ (.CLK(clknet_leaf_270_i_clk),
    .D(_01959_),
    .Q(\mem[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13267_ (.CLK(clknet_leaf_270_i_clk),
    .D(_01960_),
    .Q(\mem[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13268_ (.CLK(clknet_leaf_270_i_clk),
    .D(_01961_),
    .Q(\mem[28][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13269_ (.CLK(clknet_leaf_235_i_clk),
    .D(_01962_),
    .Q(\mem[28][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13270_ (.CLK(clknet_leaf_233_i_clk),
    .D(_01963_),
    .Q(\mem[28][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13271_ (.CLK(clknet_leaf_233_i_clk),
    .D(_01964_),
    .Q(\mem[28][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13272_ (.CLK(clknet_leaf_233_i_clk),
    .D(_01965_),
    .Q(\mem[28][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13273_ (.CLK(clknet_leaf_251_i_clk),
    .D(_01966_),
    .Q(\mem[28][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13274_ (.CLK(clknet_leaf_230_i_clk),
    .D(_01967_),
    .Q(\mem[28][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13275_ (.CLK(clknet_leaf_230_i_clk),
    .D(_01968_),
    .Q(\mem[28][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13276_ (.CLK(clknet_leaf_251_i_clk),
    .D(_01969_),
    .Q(\mem[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13277_ (.CLK(clknet_leaf_252_i_clk),
    .D(_01970_),
    .Q(\mem[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13278_ (.CLK(clknet_leaf_257_i_clk),
    .D(_01971_),
    .Q(\mem[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13279_ (.CLK(clknet_leaf_256_i_clk),
    .D(_01972_),
    .Q(\mem[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13280_ (.CLK(clknet_leaf_255_i_clk),
    .D(_01973_),
    .Q(\mem[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13281_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01974_),
    .Q(\mem[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13282_ (.CLK(clknet_leaf_256_i_clk),
    .D(_01975_),
    .Q(\mem[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13283_ (.CLK(clknet_leaf_253_i_clk),
    .D(_01976_),
    .Q(\mem[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13284_ (.CLK(clknet_leaf_253_i_clk),
    .D(_01977_),
    .Q(\mem[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13285_ (.CLK(clknet_leaf_253_i_clk),
    .D(_01978_),
    .Q(\mem[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13286_ (.CLK(clknet_leaf_251_i_clk),
    .D(_01979_),
    .Q(\mem[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13287_ (.CLK(clknet_leaf_181_i_clk),
    .D(_01980_),
    .Q(\mem[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13288_ (.CLK(clknet_leaf_182_i_clk),
    .D(_01981_),
    .Q(\mem[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13289_ (.CLK(clknet_leaf_252_i_clk),
    .D(_01982_),
    .Q(\mem[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13290_ (.CLK(clknet_leaf_183_i_clk),
    .D(_01983_),
    .Q(\mem[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13291_ (.CLK(clknet_leaf_183_i_clk),
    .D(_01984_),
    .Q(\mem[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13292_ (.CLK(clknet_leaf_240_i_clk),
    .D(_01985_),
    .Q(\mem[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13293_ (.CLK(clknet_leaf_239_i_clk),
    .D(_01986_),
    .Q(\mem[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13294_ (.CLK(clknet_leaf_238_i_clk),
    .D(_01987_),
    .Q(\mem[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13295_ (.CLK(clknet_leaf_266_i_clk),
    .D(_01988_),
    .Q(\mem[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13296_ (.CLK(clknet_leaf_270_i_clk),
    .D(_01989_),
    .Q(\mem[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13297_ (.CLK(clknet_leaf_247_i_clk),
    .D(_01990_),
    .Q(\mem[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13298_ (.CLK(clknet_leaf_236_i_clk),
    .D(_01991_),
    .Q(\mem[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13299_ (.CLK(clknet_leaf_271_i_clk),
    .D(_01992_),
    .Q(\mem[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13300_ (.CLK(clknet_leaf_235_i_clk),
    .D(_01993_),
    .Q(\mem[30][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13301_ (.CLK(clknet_leaf_236_i_clk),
    .D(_01994_),
    .Q(\mem[30][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13302_ (.CLK(clknet_leaf_233_i_clk),
    .D(_01995_),
    .Q(\mem[30][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13303_ (.CLK(clknet_leaf_233_i_clk),
    .D(_01996_),
    .Q(\mem[30][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13304_ (.CLK(clknet_leaf_233_i_clk),
    .D(_01997_),
    .Q(\mem[30][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13305_ (.CLK(clknet_leaf_250_i_clk),
    .D(_01998_),
    .Q(\mem[30][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13306_ (.CLK(clknet_leaf_229_i_clk),
    .D(_01999_),
    .Q(\mem[30][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13307_ (.CLK(clknet_leaf_230_i_clk),
    .D(_02000_),
    .Q(\mem[30][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13308_ (.CLK(clknet_leaf_239_i_clk),
    .D(_02001_),
    .Q(\mem[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13309_ (.CLK(clknet_leaf_247_i_clk),
    .D(_02002_),
    .Q(\mem[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13310_ (.CLK(clknet_leaf_238_i_clk),
    .D(_02003_),
    .Q(\mem[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13311_ (.CLK(clknet_leaf_266_i_clk),
    .D(_02004_),
    .Q(\mem[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13312_ (.CLK(clknet_leaf_270_i_clk),
    .D(_02005_),
    .Q(\mem[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13313_ (.CLK(clknet_leaf_248_i_clk),
    .D(_02006_),
    .Q(\mem[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13314_ (.CLK(clknet_leaf_236_i_clk),
    .D(_02007_),
    .Q(\mem[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13315_ (.CLK(clknet_leaf_270_i_clk),
    .D(_02008_),
    .Q(\mem[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13316_ (.CLK(clknet_leaf_236_i_clk),
    .D(_02009_),
    .Q(\mem[31][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13317_ (.CLK(clknet_leaf_236_i_clk),
    .D(_02010_),
    .Q(\mem[31][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13318_ (.CLK(clknet_leaf_233_i_clk),
    .D(_02011_),
    .Q(\mem[31][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13319_ (.CLK(clknet_leaf_233_i_clk),
    .D(_02012_),
    .Q(\mem[31][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13320_ (.CLK(clknet_leaf_233_i_clk),
    .D(_02013_),
    .Q(\mem[31][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13321_ (.CLK(clknet_leaf_250_i_clk),
    .D(_02014_),
    .Q(\mem[31][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13322_ (.CLK(clknet_leaf_229_i_clk),
    .D(_02015_),
    .Q(\mem[31][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13323_ (.CLK(clknet_leaf_231_i_clk),
    .D(_02016_),
    .Q(\mem[31][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13324_ (.CLK(clknet_leaf_7_i_clk),
    .D(_02017_),
    .Q(\mem[32][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13325_ (.CLK(clknet_leaf_25_i_clk),
    .D(_02018_),
    .Q(\mem[32][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13326_ (.CLK(clknet_leaf_282_i_clk),
    .D(_02019_),
    .Q(\mem[32][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13327_ (.CLK(clknet_leaf_287_i_clk),
    .D(_02020_),
    .Q(\mem[32][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13328_ (.CLK(clknet_leaf_0_i_clk),
    .D(_02021_),
    .Q(\mem[32][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13329_ (.CLK(clknet_leaf_21_i_clk),
    .D(_02022_),
    .Q(\mem[32][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13330_ (.CLK(clknet_leaf_0_i_clk),
    .D(_02023_),
    .Q(\mem[32][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13331_ (.CLK(clknet_leaf_0_i_clk),
    .D(_02024_),
    .Q(\mem[32][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13332_ (.CLK(clknet_leaf_1_i_clk),
    .D(_02025_),
    .Q(\mem[32][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13333_ (.CLK(clknet_leaf_12_i_clk),
    .D(_02026_),
    .Q(\mem[32][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13334_ (.CLK(clknet_leaf_15_i_clk),
    .D(_02027_),
    .Q(\mem[32][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13335_ (.CLK(clknet_leaf_13_i_clk),
    .D(_02028_),
    .Q(\mem[32][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13336_ (.CLK(clknet_leaf_14_i_clk),
    .D(_02029_),
    .Q(\mem[32][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13337_ (.CLK(clknet_leaf_28_i_clk),
    .D(_02030_),
    .Q(\mem[32][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13338_ (.CLK(clknet_leaf_11_i_clk),
    .D(_02031_),
    .Q(\mem[32][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13339_ (.CLK(clknet_leaf_28_i_clk),
    .D(_02032_),
    .Q(\mem[32][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13340_ (.CLK(clknet_leaf_7_i_clk),
    .D(_02033_),
    .Q(\mem[33][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13341_ (.CLK(clknet_leaf_22_i_clk),
    .D(_02034_),
    .Q(\mem[33][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13342_ (.CLK(clknet_leaf_282_i_clk),
    .D(_02035_),
    .Q(\mem[33][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13343_ (.CLK(clknet_leaf_288_i_clk),
    .D(_02036_),
    .Q(\mem[33][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13344_ (.CLK(clknet_leaf_288_i_clk),
    .D(_02037_),
    .Q(\mem[33][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13345_ (.CLK(clknet_leaf_21_i_clk),
    .D(_02038_),
    .Q(\mem[33][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13346_ (.CLK(clknet_leaf_0_i_clk),
    .D(_02039_),
    .Q(\mem[33][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13347_ (.CLK(clknet_leaf_0_i_clk),
    .D(_02040_),
    .Q(\mem[33][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13348_ (.CLK(clknet_leaf_2_i_clk),
    .D(_02041_),
    .Q(\mem[33][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13349_ (.CLK(clknet_leaf_13_i_clk),
    .D(_02042_),
    .Q(\mem[33][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13350_ (.CLK(clknet_leaf_15_i_clk),
    .D(_02043_),
    .Q(\mem[33][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13351_ (.CLK(clknet_leaf_13_i_clk),
    .D(_02044_),
    .Q(\mem[33][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13352_ (.CLK(clknet_leaf_14_i_clk),
    .D(_02045_),
    .Q(\mem[33][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13353_ (.CLK(clknet_leaf_28_i_clk),
    .D(_02046_),
    .Q(\mem[33][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13354_ (.CLK(clknet_leaf_11_i_clk),
    .D(_02047_),
    .Q(\mem[33][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13355_ (.CLK(clknet_leaf_28_i_clk),
    .D(_02048_),
    .Q(\mem[33][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13356_ (.CLK(clknet_leaf_9_i_clk),
    .D(_02049_),
    .Q(\mem[34][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13357_ (.CLK(clknet_leaf_21_i_clk),
    .D(_02050_),
    .Q(\mem[34][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13358_ (.CLK(clknet_leaf_282_i_clk),
    .D(_02051_),
    .Q(\mem[34][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13359_ (.CLK(clknet_leaf_287_i_clk),
    .D(_02052_),
    .Q(\mem[34][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13360_ (.CLK(clknet_leaf_0_i_clk),
    .D(_02053_),
    .Q(\mem[34][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13361_ (.CLK(clknet_leaf_21_i_clk),
    .D(_02054_),
    .Q(\mem[34][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13362_ (.CLK(clknet_leaf_0_i_clk),
    .D(_02055_),
    .Q(\mem[34][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13363_ (.CLK(clknet_leaf_0_i_clk),
    .D(_02056_),
    .Q(\mem[34][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13364_ (.CLK(clknet_leaf_2_i_clk),
    .D(_02057_),
    .Q(\mem[34][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13365_ (.CLK(clknet_leaf_13_i_clk),
    .D(_02058_),
    .Q(\mem[34][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13366_ (.CLK(clknet_leaf_15_i_clk),
    .D(_02059_),
    .Q(\mem[34][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13367_ (.CLK(clknet_leaf_13_i_clk),
    .D(_02060_),
    .Q(\mem[34][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13368_ (.CLK(clknet_leaf_14_i_clk),
    .D(_02061_),
    .Q(\mem[34][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13369_ (.CLK(clknet_leaf_27_i_clk),
    .D(_02062_),
    .Q(\mem[34][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13370_ (.CLK(clknet_leaf_11_i_clk),
    .D(_02063_),
    .Q(\mem[34][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13371_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00016_),
    .Q(\mem[34][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13372_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00017_),
    .Q(\mem[35][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13373_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00018_),
    .Q(\mem[35][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13374_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00019_),
    .Q(\mem[35][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13375_ (.CLK(clknet_leaf_287_i_clk),
    .D(_00020_),
    .Q(\mem[35][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13376_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00021_),
    .Q(\mem[35][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13377_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00022_),
    .Q(\mem[35][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13378_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00023_),
    .Q(\mem[35][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13379_ (.CLK(clknet_leaf_0_i_clk),
    .D(_00024_),
    .Q(\mem[35][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13380_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00025_),
    .Q(\mem[35][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13381_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00026_),
    .Q(\mem[35][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13382_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00027_),
    .Q(\mem[35][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13383_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00028_),
    .Q(\mem[35][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13384_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00029_),
    .Q(\mem[35][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13385_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00030_),
    .Q(\mem[35][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13386_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00031_),
    .Q(\mem[35][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13387_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00032_),
    .Q(\mem[35][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13388_ (.CLK(clknet_leaf_280_i_clk),
    .D(_00033_),
    .Q(\mem[36][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13389_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00034_),
    .Q(\mem[36][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13390_ (.CLK(clknet_leaf_283_i_clk),
    .D(_00035_),
    .Q(\mem[36][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13391_ (.CLK(clknet_leaf_286_i_clk),
    .D(_00036_),
    .Q(\mem[36][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13392_ (.CLK(clknet_leaf_288_i_clk),
    .D(_00037_),
    .Q(\mem[36][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13393_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00038_),
    .Q(\mem[36][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13394_ (.CLK(clknet_leaf_283_i_clk),
    .D(_00039_),
    .Q(\mem[36][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13395_ (.CLK(clknet_leaf_286_i_clk),
    .D(_00040_),
    .Q(\mem[36][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13396_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00041_),
    .Q(\mem[36][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13397_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00042_),
    .Q(\mem[36][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13398_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00043_),
    .Q(\mem[36][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13399_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00044_),
    .Q(\mem[36][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13400_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00045_),
    .Q(\mem[36][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13401_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00046_),
    .Q(\mem[36][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13402_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00047_),
    .Q(\mem[36][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13403_ (.CLK(clknet_leaf_8_i_clk),
    .D(_00048_),
    .Q(\mem[36][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13404_ (.CLK(clknet_leaf_7_i_clk),
    .D(_00049_),
    .Q(\mem[37][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13405_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00050_),
    .Q(\mem[37][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13406_ (.CLK(clknet_leaf_283_i_clk),
    .D(_00051_),
    .Q(\mem[37][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13407_ (.CLK(clknet_leaf_286_i_clk),
    .D(_00052_),
    .Q(\mem[37][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13408_ (.CLK(clknet_leaf_288_i_clk),
    .D(_00053_),
    .Q(\mem[37][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13409_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00054_),
    .Q(\mem[37][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13410_ (.CLK(clknet_leaf_287_i_clk),
    .D(_00055_),
    .Q(\mem[37][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13411_ (.CLK(clknet_leaf_283_i_clk),
    .D(_00056_),
    .Q(\mem[37][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13412_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00057_),
    .Q(\mem[37][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13413_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00058_),
    .Q(\mem[37][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13414_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00059_),
    .Q(\mem[37][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13415_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00060_),
    .Q(\mem[37][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13416_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00061_),
    .Q(\mem[37][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13417_ (.CLK(clknet_leaf_27_i_clk),
    .D(_00062_),
    .Q(\mem[37][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13418_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00063_),
    .Q(\mem[37][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13419_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00064_),
    .Q(\mem[37][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13420_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00065_),
    .Q(\mem[38][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13421_ (.CLK(clknet_leaf_26_i_clk),
    .D(_00066_),
    .Q(\mem[38][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13422_ (.CLK(clknet_leaf_282_i_clk),
    .D(_00067_),
    .Q(\mem[38][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13423_ (.CLK(clknet_leaf_288_i_clk),
    .D(_00068_),
    .Q(\mem[38][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13424_ (.CLK(clknet_leaf_288_i_clk),
    .D(_00069_),
    .Q(\mem[38][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13425_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00070_),
    .Q(\mem[38][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13426_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00071_),
    .Q(\mem[38][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13427_ (.CLK(clknet_leaf_286_i_clk),
    .D(_00072_),
    .Q(\mem[38][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13428_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00073_),
    .Q(\mem[38][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13429_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00074_),
    .Q(\mem[38][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13430_ (.CLK(clknet_leaf_15_i_clk),
    .D(_00075_),
    .Q(\mem[38][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13431_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00076_),
    .Q(\mem[38][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13432_ (.CLK(clknet_leaf_10_i_clk),
    .D(_00077_),
    .Q(\mem[38][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13433_ (.CLK(clknet_leaf_25_i_clk),
    .D(_00078_),
    .Q(\mem[38][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13434_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00079_),
    .Q(\mem[38][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13435_ (.CLK(clknet_leaf_9_i_clk),
    .D(_00080_),
    .Q(\mem[38][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13436_ (.CLK(clknet_leaf_32_i_clk),
    .D(_00081_),
    .Q(\mem[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13437_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00082_),
    .Q(\mem[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13438_ (.CLK(clknet_leaf_259_i_clk),
    .D(_00083_),
    .Q(\mem[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13439_ (.CLK(clknet_leaf_260_i_clk),
    .D(_00084_),
    .Q(\mem[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13440_ (.CLK(clknet_leaf_260_i_clk),
    .D(_00085_),
    .Q(\mem[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13441_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00086_),
    .Q(\mem[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13442_ (.CLK(clknet_leaf_259_i_clk),
    .D(_00087_),
    .Q(\mem[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13443_ (.CLK(clknet_leaf_255_i_clk),
    .D(_00088_),
    .Q(\mem[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13444_ (.CLK(clknet_leaf_254_i_clk),
    .D(_00089_),
    .Q(\mem[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13445_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00090_),
    .Q(\mem[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13446_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00091_),
    .Q(\mem[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13447_ (.CLK(clknet_leaf_254_i_clk),
    .D(_00092_),
    .Q(\mem[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13448_ (.CLK(clknet_leaf_36_i_clk),
    .D(_00093_),
    .Q(\mem[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13449_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00094_),
    .Q(\mem[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13450_ (.CLK(clknet_leaf_35_i_clk),
    .D(_00095_),
    .Q(\mem[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13451_ (.CLK(clknet_leaf_37_i_clk),
    .D(_00096_),
    .Q(\mem[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13452_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00097_),
    .Q(\mem[40][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13453_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00098_),
    .Q(\mem[40][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13454_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00099_),
    .Q(\mem[40][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13455_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00100_),
    .Q(\mem[40][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13456_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00101_),
    .Q(\mem[40][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13457_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00102_),
    .Q(\mem[40][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13458_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00103_),
    .Q(\mem[40][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13459_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00104_),
    .Q(\mem[40][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13460_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00105_),
    .Q(\mem[40][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13461_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00106_),
    .Q(\mem[40][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13462_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00107_),
    .Q(\mem[40][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13463_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00108_),
    .Q(\mem[40][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13464_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00109_),
    .Q(\mem[40][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13465_ (.CLK(clknet_leaf_23_i_clk),
    .D(_00110_),
    .Q(\mem[40][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13466_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00111_),
    .Q(\mem[40][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13467_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00112_),
    .Q(\mem[40][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13468_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00113_),
    .Q(\mem[41][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13469_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00114_),
    .Q(\mem[41][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13470_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00115_),
    .Q(\mem[41][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13471_ (.CLK(clknet_leaf_1_i_clk),
    .D(_00116_),
    .Q(\mem[41][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13472_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00117_),
    .Q(\mem[41][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13473_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00118_),
    .Q(\mem[41][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13474_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00119_),
    .Q(\mem[41][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13475_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00120_),
    .Q(\mem[41][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13476_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00121_),
    .Q(\mem[41][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13477_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00122_),
    .Q(\mem[41][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13478_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00123_),
    .Q(\mem[41][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13479_ (.CLK(clknet_leaf_19_i_clk),
    .D(_00124_),
    .Q(\mem[41][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13480_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00125_),
    .Q(\mem[41][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13481_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00126_),
    .Q(\mem[41][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13482_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00127_),
    .Q(\mem[41][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13483_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00128_),
    .Q(\mem[41][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13484_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00129_),
    .Q(\mem[42][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13485_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00130_),
    .Q(\mem[42][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13486_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00131_),
    .Q(\mem[42][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13487_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00132_),
    .Q(\mem[42][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13488_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00133_),
    .Q(\mem[42][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13489_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00134_),
    .Q(\mem[42][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13490_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00135_),
    .Q(\mem[42][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13491_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00136_),
    .Q(\mem[42][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13492_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00137_),
    .Q(\mem[42][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13493_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00138_),
    .Q(\mem[42][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13494_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00139_),
    .Q(\mem[42][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13495_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00140_),
    .Q(\mem[42][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13496_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00141_),
    .Q(\mem[42][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13497_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00142_),
    .Q(\mem[42][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13498_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00143_),
    .Q(\mem[42][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13499_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00144_),
    .Q(\mem[42][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13500_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00145_),
    .Q(\mem[43][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13501_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00146_),
    .Q(\mem[43][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13502_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00147_),
    .Q(\mem[43][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13503_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00148_),
    .Q(\mem[43][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13504_ (.CLK(clknet_leaf_2_i_clk),
    .D(_00149_),
    .Q(\mem[43][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13505_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00150_),
    .Q(\mem[43][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13506_ (.CLK(clknet_leaf_13_i_clk),
    .D(_00151_),
    .Q(\mem[43][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13507_ (.CLK(clknet_leaf_14_i_clk),
    .D(_00152_),
    .Q(\mem[43][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13508_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00153_),
    .Q(\mem[43][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13509_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00154_),
    .Q(\mem[43][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13510_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00155_),
    .Q(\mem[43][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13511_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00156_),
    .Q(\mem[43][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13512_ (.CLK(clknet_leaf_18_i_clk),
    .D(_00157_),
    .Q(\mem[43][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13513_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00158_),
    .Q(\mem[43][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13514_ (.CLK(clknet_leaf_20_i_clk),
    .D(_00159_),
    .Q(\mem[43][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13515_ (.CLK(clknet_leaf_22_i_clk),
    .D(_00160_),
    .Q(\mem[43][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13516_ (.CLK(clknet_leaf_11_i_clk),
    .D(_00161_),
    .Q(\mem[44][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13517_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00162_),
    .Q(\mem[44][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13518_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00163_),
    .Q(\mem[44][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13519_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00164_),
    .Q(\mem[44][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13520_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00165_),
    .Q(\mem[44][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13521_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00166_),
    .Q(\mem[44][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13522_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00167_),
    .Q(\mem[44][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13523_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00168_),
    .Q(\mem[44][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13524_ (.CLK(clknet_leaf_21_i_clk),
    .D(_00169_),
    .Q(\mem[44][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13525_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00170_),
    .Q(\mem[44][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13526_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00171_),
    .Q(\mem[44][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13527_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00172_),
    .Q(\mem[44][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13528_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00173_),
    .Q(\mem[44][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13529_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00174_),
    .Q(\mem[44][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13530_ (.CLK(clknet_leaf_55_i_clk),
    .D(_00175_),
    .Q(\mem[44][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13531_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00176_),
    .Q(\mem[44][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13532_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00177_),
    .Q(\mem[45][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13533_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00178_),
    .Q(\mem[45][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13534_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00179_),
    .Q(\mem[45][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13535_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00180_),
    .Q(\mem[45][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13536_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00181_),
    .Q(\mem[45][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13537_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00182_),
    .Q(\mem[45][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13538_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00183_),
    .Q(\mem[45][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13539_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00184_),
    .Q(\mem[45][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13540_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00185_),
    .Q(\mem[45][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13541_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00186_),
    .Q(\mem[45][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13542_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00187_),
    .Q(\mem[45][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13543_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00188_),
    .Q(\mem[45][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13544_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00189_),
    .Q(\mem[45][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13545_ (.CLK(clknet_leaf_52_i_clk),
    .D(_00190_),
    .Q(\mem[45][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13546_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00191_),
    .Q(\mem[45][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13547_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00192_),
    .Q(\mem[45][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13548_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00193_),
    .Q(\mem[46][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13549_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00194_),
    .Q(\mem[46][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13550_ (.CLK(clknet_leaf_6_i_clk),
    .D(_00195_),
    .Q(\mem[46][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13551_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00196_),
    .Q(\mem[46][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13552_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00197_),
    .Q(\mem[46][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13553_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00198_),
    .Q(\mem[46][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13554_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00199_),
    .Q(\mem[46][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13555_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00200_),
    .Q(\mem[46][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13556_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00201_),
    .Q(\mem[46][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13557_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00202_),
    .Q(\mem[46][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13558_ (.CLK(clknet_leaf_57_i_clk),
    .D(_00203_),
    .Q(\mem[46][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13559_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00204_),
    .Q(\mem[46][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13560_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00205_),
    .Q(\mem[46][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13561_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00206_),
    .Q(\mem[46][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13562_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00207_),
    .Q(\mem[46][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13563_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00208_),
    .Q(\mem[46][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13564_ (.CLK(clknet_leaf_12_i_clk),
    .D(_00209_),
    .Q(\mem[47][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13565_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00210_),
    .Q(\mem[47][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13566_ (.CLK(clknet_leaf_5_i_clk),
    .D(_00211_),
    .Q(\mem[47][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13567_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00212_),
    .Q(\mem[47][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13568_ (.CLK(clknet_leaf_3_i_clk),
    .D(_00213_),
    .Q(\mem[47][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13569_ (.CLK(clknet_leaf_56_i_clk),
    .D(_00214_),
    .Q(\mem[47][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13570_ (.CLK(clknet_leaf_4_i_clk),
    .D(_00215_),
    .Q(\mem[47][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13571_ (.CLK(clknet_leaf_17_i_clk),
    .D(_00216_),
    .Q(\mem[47][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13572_ (.CLK(clknet_leaf_16_i_clk),
    .D(_00217_),
    .Q(\mem[47][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13573_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00218_),
    .Q(\mem[47][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13574_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00219_),
    .Q(\mem[47][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13575_ (.CLK(clknet_leaf_58_i_clk),
    .D(_00220_),
    .Q(\mem[47][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13576_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00221_),
    .Q(\mem[47][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13577_ (.CLK(clknet_leaf_53_i_clk),
    .D(_00222_),
    .Q(\mem[47][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13578_ (.CLK(clknet_leaf_59_i_clk),
    .D(_00223_),
    .Q(\mem[47][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13579_ (.CLK(clknet_leaf_54_i_clk),
    .D(_00224_),
    .Q(\mem[47][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13580_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00225_),
    .Q(\mem[48][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13581_ (.CLK(clknet_leaf_47_i_clk),
    .D(_00226_),
    .Q(\mem[48][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13582_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00227_),
    .Q(\mem[48][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13583_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00228_),
    .Q(\mem[48][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13584_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00229_),
    .Q(\mem[48][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13585_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00230_),
    .Q(\mem[48][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13586_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00231_),
    .Q(\mem[48][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13587_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00232_),
    .Q(\mem[48][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13588_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00233_),
    .Q(\mem[48][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13589_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00234_),
    .Q(\mem[48][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13590_ (.CLK(clknet_leaf_105_i_clk),
    .D(_00235_),
    .Q(\mem[48][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13591_ (.CLK(clknet_leaf_102_i_clk),
    .D(_00236_),
    .Q(\mem[48][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13592_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00237_),
    .Q(\mem[48][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13593_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00238_),
    .Q(\mem[48][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13594_ (.CLK(clknet_leaf_103_i_clk),
    .D(_00239_),
    .Q(\mem[48][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13595_ (.CLK(clknet_leaf_102_i_clk),
    .D(_00240_),
    .Q(\mem[48][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13596_ (.CLK(clknet_leaf_160_i_clk),
    .D(_00241_),
    .Q(\mem[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13597_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00242_),
    .Q(\mem[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13598_ (.CLK(clknet_leaf_164_i_clk),
    .D(_00243_),
    .Q(\mem[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13599_ (.CLK(clknet_leaf_163_i_clk),
    .D(_00244_),
    .Q(\mem[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13600_ (.CLK(clknet_leaf_162_i_clk),
    .D(_00245_),
    .Q(\mem[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13601_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00246_),
    .Q(\mem[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13602_ (.CLK(clknet_leaf_159_i_clk),
    .D(_00247_),
    .Q(\mem[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13603_ (.CLK(clknet_leaf_161_i_clk),
    .D(_00248_),
    .Q(\mem[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13604_ (.CLK(clknet_leaf_161_i_clk),
    .D(_00249_),
    .Q(\mem[4][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13605_ (.CLK(clknet_leaf_160_i_clk),
    .D(_00250_),
    .Q(\mem[4][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13606_ (.CLK(clknet_leaf_156_i_clk),
    .D(_00251_),
    .Q(\mem[4][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13607_ (.CLK(clknet_leaf_139_i_clk),
    .D(_00252_),
    .Q(\mem[4][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13608_ (.CLK(clknet_leaf_156_i_clk),
    .D(_00253_),
    .Q(\mem[4][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13609_ (.CLK(clknet_leaf_117_i_clk),
    .D(_00254_),
    .Q(\mem[4][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13610_ (.CLK(clknet_leaf_140_i_clk),
    .D(_00255_),
    .Q(\mem[4][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13611_ (.CLK(clknet_leaf_139_i_clk),
    .D(_00256_),
    .Q(\mem[4][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13612_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00257_),
    .Q(\mem[50][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13613_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00258_),
    .Q(\mem[50][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13614_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00259_),
    .Q(\mem[50][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13615_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00260_),
    .Q(\mem[50][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13616_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00261_),
    .Q(\mem[50][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13617_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00262_),
    .Q(\mem[50][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13618_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00263_),
    .Q(\mem[50][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13619_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00264_),
    .Q(\mem[50][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13620_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00265_),
    .Q(\mem[50][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13621_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00266_),
    .Q(\mem[50][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13622_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00267_),
    .Q(\mem[50][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13623_ (.CLK(clknet_leaf_105_i_clk),
    .D(_00268_),
    .Q(\mem[50][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13624_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00269_),
    .Q(\mem[50][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13625_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00270_),
    .Q(\mem[50][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13626_ (.CLK(clknet_leaf_103_i_clk),
    .D(_00271_),
    .Q(\mem[50][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13627_ (.CLK(clknet_leaf_102_i_clk),
    .D(_00272_),
    .Q(\mem[50][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13628_ (.CLK(clknet_leaf_60_i_clk),
    .D(_00273_),
    .Q(\mem[51][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13629_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00274_),
    .Q(\mem[51][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13630_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00275_),
    .Q(\mem[51][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13631_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00276_),
    .Q(\mem[51][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13632_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00277_),
    .Q(\mem[51][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13633_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00278_),
    .Q(\mem[51][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13634_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00279_),
    .Q(\mem[51][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13635_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00280_),
    .Q(\mem[51][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13636_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00281_),
    .Q(\mem[51][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13637_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00282_),
    .Q(\mem[51][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13638_ (.CLK(clknet_leaf_105_i_clk),
    .D(_00283_),
    .Q(\mem[51][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13639_ (.CLK(clknet_leaf_105_i_clk),
    .D(_00284_),
    .Q(\mem[51][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13640_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00285_),
    .Q(\mem[51][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13641_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00286_),
    .Q(\mem[51][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13642_ (.CLK(clknet_leaf_104_i_clk),
    .D(_00287_),
    .Q(\mem[51][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13643_ (.CLK(clknet_leaf_102_i_clk),
    .D(_00288_),
    .Q(\mem[51][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13644_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00289_),
    .Q(\mem[52][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13645_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00290_),
    .Q(\mem[52][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13646_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00291_),
    .Q(\mem[52][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13647_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00292_),
    .Q(\mem[52][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13648_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00293_),
    .Q(\mem[52][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13649_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00294_),
    .Q(\mem[52][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13650_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00295_),
    .Q(\mem[52][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13651_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00296_),
    .Q(\mem[52][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13652_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00297_),
    .Q(\mem[52][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13653_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00298_),
    .Q(\mem[52][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13654_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00299_),
    .Q(\mem[52][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13655_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00300_),
    .Q(\mem[52][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13656_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00301_),
    .Q(\mem[52][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13657_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00302_),
    .Q(\mem[52][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13658_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00303_),
    .Q(\mem[52][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13659_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00304_),
    .Q(\mem[52][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13660_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00305_),
    .Q(\mem[53][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13661_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00306_),
    .Q(\mem[53][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13662_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00307_),
    .Q(\mem[53][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13663_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00308_),
    .Q(\mem[53][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13664_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00309_),
    .Q(\mem[53][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13665_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00310_),
    .Q(\mem[53][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13666_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00311_),
    .Q(\mem[53][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13667_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00312_),
    .Q(\mem[53][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13668_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00313_),
    .Q(\mem[53][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13669_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00314_),
    .Q(\mem[53][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13670_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00315_),
    .Q(\mem[53][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13671_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00316_),
    .Q(\mem[53][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13672_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00317_),
    .Q(\mem[53][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13673_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00318_),
    .Q(\mem[53][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13674_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00319_),
    .Q(\mem[53][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13675_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00320_),
    .Q(\mem[53][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13676_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00321_),
    .Q(\mem[54][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13677_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00322_),
    .Q(\mem[54][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13678_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00323_),
    .Q(\mem[54][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13679_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00324_),
    .Q(\mem[54][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13680_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00325_),
    .Q(\mem[54][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13681_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00326_),
    .Q(\mem[54][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13682_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00327_),
    .Q(\mem[54][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13683_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00328_),
    .Q(\mem[54][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13684_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00329_),
    .Q(\mem[54][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13685_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00330_),
    .Q(\mem[54][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13686_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00331_),
    .Q(\mem[54][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13687_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00332_),
    .Q(\mem[54][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13688_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00333_),
    .Q(\mem[54][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13689_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00334_),
    .Q(\mem[54][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13690_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00335_),
    .Q(\mem[54][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13691_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00336_),
    .Q(\mem[54][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13692_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00337_),
    .Q(\mem[55][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13693_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00338_),
    .Q(\mem[55][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13694_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00339_),
    .Q(\mem[55][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13695_ (.CLK(clknet_leaf_74_i_clk),
    .D(_00340_),
    .Q(\mem[55][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13696_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00341_),
    .Q(\mem[55][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13697_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00342_),
    .Q(\mem[55][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13698_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00343_),
    .Q(\mem[55][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13699_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00344_),
    .Q(\mem[55][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13700_ (.CLK(clknet_leaf_77_i_clk),
    .D(_00345_),
    .Q(\mem[55][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13701_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00346_),
    .Q(\mem[55][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13702_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00347_),
    .Q(\mem[55][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13703_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00348_),
    .Q(\mem[55][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13704_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00349_),
    .Q(\mem[55][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13705_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00350_),
    .Q(\mem[55][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13706_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00351_),
    .Q(\mem[55][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13707_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00352_),
    .Q(\mem[55][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13708_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00353_),
    .Q(\mem[56][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13709_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00354_),
    .Q(\mem[56][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13710_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00355_),
    .Q(\mem[56][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13711_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00356_),
    .Q(\mem[56][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13712_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00357_),
    .Q(\mem[56][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13713_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00358_),
    .Q(\mem[56][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13714_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00359_),
    .Q(\mem[56][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13715_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00360_),
    .Q(\mem[56][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13716_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00361_),
    .Q(\mem[56][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13717_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00362_),
    .Q(\mem[56][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13718_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00363_),
    .Q(\mem[56][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13719_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00364_),
    .Q(\mem[56][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13720_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00365_),
    .Q(\mem[56][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13721_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00366_),
    .Q(\mem[56][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13722_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00367_),
    .Q(\mem[56][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13723_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00368_),
    .Q(\mem[56][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13724_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00369_),
    .Q(\mem[57][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13725_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00370_),
    .Q(\mem[57][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13726_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00371_),
    .Q(\mem[57][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13727_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00372_),
    .Q(\mem[57][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13728_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00373_),
    .Q(\mem[57][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13729_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00374_),
    .Q(\mem[57][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13730_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00375_),
    .Q(\mem[57][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13731_ (.CLK(clknet_leaf_83_i_clk),
    .D(_00376_),
    .Q(\mem[57][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13732_ (.CLK(clknet_leaf_79_i_clk),
    .D(_00377_),
    .Q(\mem[57][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13733_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00378_),
    .Q(\mem[57][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13734_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00379_),
    .Q(\mem[57][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13735_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00380_),
    .Q(\mem[57][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13736_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00381_),
    .Q(\mem[57][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13737_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00382_),
    .Q(\mem[57][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13738_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00383_),
    .Q(\mem[57][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13739_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00384_),
    .Q(\mem[57][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13740_ (.CLK(clknet_leaf_71_i_clk),
    .D(_00385_),
    .Q(\mem[58][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13741_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00386_),
    .Q(\mem[58][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13742_ (.CLK(clknet_leaf_75_i_clk),
    .D(_00387_),
    .Q(\mem[58][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13743_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00388_),
    .Q(\mem[58][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13744_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00389_),
    .Q(\mem[58][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13745_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00390_),
    .Q(\mem[58][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13746_ (.CLK(clknet_leaf_76_i_clk),
    .D(_00391_),
    .Q(\mem[58][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13747_ (.CLK(clknet_leaf_84_i_clk),
    .D(_00392_),
    .Q(\mem[58][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13748_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00393_),
    .Q(\mem[58][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13749_ (.CLK(clknet_leaf_78_i_clk),
    .D(_00394_),
    .Q(\mem[58][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13750_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00395_),
    .Q(\mem[58][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13751_ (.CLK(clknet_leaf_80_i_clk),
    .D(_00396_),
    .Q(\mem[58][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13752_ (.CLK(clknet_leaf_81_i_clk),
    .D(_00397_),
    .Q(\mem[58][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13753_ (.CLK(clknet_leaf_82_i_clk),
    .D(_00398_),
    .Q(\mem[58][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13754_ (.CLK(clknet_leaf_90_i_clk),
    .D(_00399_),
    .Q(\mem[58][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13755_ (.CLK(clknet_leaf_89_i_clk),
    .D(_00400_),
    .Q(\mem[58][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13756_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00401_),
    .Q(\mem[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13757_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00402_),
    .Q(\mem[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13758_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00403_),
    .Q(\mem[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13759_ (.CLK(clknet_leaf_115_i_clk),
    .D(_00404_),
    .Q(\mem[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13760_ (.CLK(clknet_leaf_118_i_clk),
    .D(_00405_),
    .Q(\mem[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13761_ (.CLK(clknet_leaf_116_i_clk),
    .D(_00406_),
    .Q(\mem[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13762_ (.CLK(clknet_leaf_118_i_clk),
    .D(_00407_),
    .Q(\mem[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13763_ (.CLK(clknet_leaf_118_i_clk),
    .D(_00408_),
    .Q(\mem[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13764_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00409_),
    .Q(\mem[5][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13765_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00410_),
    .Q(\mem[5][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13766_ (.CLK(clknet_leaf_120_i_clk),
    .D(_00411_),
    .Q(\mem[5][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13767_ (.CLK(clknet_leaf_120_i_clk),
    .D(_00412_),
    .Q(\mem[5][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13768_ (.CLK(clknet_leaf_121_i_clk),
    .D(_00413_),
    .Q(\mem[5][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13769_ (.CLK(clknet_leaf_117_i_clk),
    .D(_00414_),
    .Q(\mem[5][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13770_ (.CLK(clknet_leaf_121_i_clk),
    .D(_00415_),
    .Q(\mem[5][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13771_ (.CLK(clknet_leaf_121_i_clk),
    .D(_00416_),
    .Q(\mem[5][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13772_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00417_),
    .Q(\mem[60][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13773_ (.CLK(clknet_leaf_50_i_clk),
    .D(_00418_),
    .Q(\mem[60][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13774_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00419_),
    .Q(\mem[60][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13775_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00420_),
    .Q(\mem[60][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13776_ (.CLK(clknet_leaf_65_i_clk),
    .D(_00421_),
    .Q(\mem[60][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13777_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00422_),
    .Q(\mem[60][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13778_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00423_),
    .Q(\mem[60][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13779_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00424_),
    .Q(\mem[60][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13780_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00425_),
    .Q(\mem[60][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13781_ (.CLK(clknet_leaf_48_i_clk),
    .D(_00426_),
    .Q(\mem[60][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13782_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00427_),
    .Q(\mem[60][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13783_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00428_),
    .Q(\mem[60][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13784_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00429_),
    .Q(\mem[60][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13785_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00430_),
    .Q(\mem[60][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13786_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00431_),
    .Q(\mem[60][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13787_ (.CLK(clknet_leaf_102_i_clk),
    .D(_00432_),
    .Q(\mem[60][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13788_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00433_),
    .Q(\mem[61][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13789_ (.CLK(clknet_leaf_67_i_clk),
    .D(_00434_),
    .Q(\mem[61][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13790_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00435_),
    .Q(\mem[61][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13791_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00436_),
    .Q(\mem[61][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13792_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00437_),
    .Q(\mem[61][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13793_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00438_),
    .Q(\mem[61][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13794_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00439_),
    .Q(\mem[61][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13795_ (.CLK(clknet_leaf_73_i_clk),
    .D(_00440_),
    .Q(\mem[61][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13796_ (.CLK(clknet_leaf_72_i_clk),
    .D(_00441_),
    .Q(\mem[61][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13797_ (.CLK(clknet_leaf_49_i_clk),
    .D(_00442_),
    .Q(\mem[61][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13798_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00443_),
    .Q(\mem[61][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13799_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00444_),
    .Q(\mem[61][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13800_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00445_),
    .Q(\mem[61][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13801_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00446_),
    .Q(\mem[61][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13802_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00447_),
    .Q(\mem[61][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13803_ (.CLK(clknet_leaf_103_i_clk),
    .D(_00448_),
    .Q(\mem[61][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13804_ (.CLK(clknet_leaf_61_i_clk),
    .D(_00449_),
    .Q(\mem[62][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13805_ (.CLK(clknet_leaf_51_i_clk),
    .D(_00450_),
    .Q(\mem[62][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13806_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00451_),
    .Q(\mem[62][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13807_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00452_),
    .Q(\mem[62][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13808_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00453_),
    .Q(\mem[62][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13809_ (.CLK(clknet_leaf_70_i_clk),
    .D(_00454_),
    .Q(\mem[62][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13810_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00455_),
    .Q(\mem[62][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13811_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00456_),
    .Q(\mem[62][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13812_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00457_),
    .Q(\mem[62][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13813_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00458_),
    .Q(\mem[62][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13814_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00459_),
    .Q(\mem[62][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13815_ (.CLK(clknet_leaf_86_i_clk),
    .D(_00460_),
    .Q(\mem[62][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13816_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00461_),
    .Q(\mem[62][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13817_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00462_),
    .Q(\mem[62][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13818_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00463_),
    .Q(\mem[62][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13819_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00464_),
    .Q(\mem[62][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13820_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00465_),
    .Q(\mem[63][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13821_ (.CLK(clknet_leaf_66_i_clk),
    .D(_00466_),
    .Q(\mem[63][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13822_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00467_),
    .Q(\mem[63][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13823_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00468_),
    .Q(\mem[63][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13824_ (.CLK(clknet_leaf_62_i_clk),
    .D(_00469_),
    .Q(\mem[63][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13825_ (.CLK(clknet_leaf_68_i_clk),
    .D(_00470_),
    .Q(\mem[63][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13826_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00471_),
    .Q(\mem[63][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13827_ (.CLK(clknet_leaf_63_i_clk),
    .D(_00472_),
    .Q(\mem[63][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13828_ (.CLK(clknet_leaf_64_i_clk),
    .D(_00473_),
    .Q(\mem[63][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13829_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00474_),
    .Q(\mem[63][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13830_ (.CLK(clknet_leaf_69_i_clk),
    .D(_00475_),
    .Q(\mem[63][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13831_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00476_),
    .Q(\mem[63][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13832_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00477_),
    .Q(\mem[63][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13833_ (.CLK(clknet_leaf_85_i_clk),
    .D(_00478_),
    .Q(\mem[63][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13834_ (.CLK(clknet_leaf_87_i_clk),
    .D(_00479_),
    .Q(\mem[63][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13835_ (.CLK(clknet_leaf_103_i_clk),
    .D(_00480_),
    .Q(\mem[63][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13836_ (.CLK(clknet_leaf_198_i_clk),
    .D(_00481_),
    .Q(\mem[64][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13837_ (.CLK(clknet_leaf_168_i_clk),
    .D(_00482_),
    .Q(\mem[64][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13838_ (.CLK(clknet_leaf_198_i_clk),
    .D(_00483_),
    .Q(\mem[64][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13839_ (.CLK(clknet_leaf_199_i_clk),
    .D(_00484_),
    .Q(\mem[64][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13840_ (.CLK(clknet_leaf_165_i_clk),
    .D(_00485_),
    .Q(\mem[64][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13841_ (.CLK(clknet_leaf_168_i_clk),
    .D(_00486_),
    .Q(\mem[64][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13842_ (.CLK(clknet_leaf_169_i_clk),
    .D(_00487_),
    .Q(\mem[64][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13843_ (.CLK(clknet_leaf_167_i_clk),
    .D(_00488_),
    .Q(\mem[64][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13844_ (.CLK(clknet_leaf_166_i_clk),
    .D(_00489_),
    .Q(\mem[64][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13845_ (.CLK(clknet_leaf_167_i_clk),
    .D(_00490_),
    .Q(\mem[64][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13846_ (.CLK(clknet_leaf_168_i_clk),
    .D(_00491_),
    .Q(\mem[64][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13847_ (.CLK(clknet_leaf_177_i_clk),
    .D(_00492_),
    .Q(\mem[64][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13848_ (.CLK(clknet_leaf_168_i_clk),
    .D(_00493_),
    .Q(\mem[64][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13849_ (.CLK(clknet_leaf_177_i_clk),
    .D(_00494_),
    .Q(\mem[64][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13850_ (.CLK(clknet_leaf_169_i_clk),
    .D(_00495_),
    .Q(\mem[64][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13851_ (.CLK(clknet_leaf_177_i_clk),
    .D(_00496_),
    .Q(\mem[64][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13852_ (.CLK(clknet_leaf_167_i_clk),
    .D(_00497_),
    .Q(\mem[65][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13853_ (.CLK(clknet_leaf_167_i_clk),
    .D(_00498_),
    .Q(\mem[65][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13854_ (.CLK(clknet_leaf_167_i_clk),
    .D(_00499_),
    .Q(\mem[65][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13855_ (.CLK(clknet_leaf_166_i_clk),
    .D(_00500_),
    .Q(\mem[65][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13856_ (.CLK(clknet_leaf_165_i_clk),
    .D(_00501_),
    .Q(\mem[65][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13857_ (.CLK(clknet_leaf_167_i_clk),
    .D(_00502_),
    .Q(\mem[65][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13858_ (.CLK(clknet_leaf_168_i_clk),
    .D(_00503_),
    .Q(\mem[65][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13859_ (.CLK(clknet_leaf_165_i_clk),
    .D(_00504_),
    .Q(\mem[65][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13860_ (.CLK(clknet_leaf_165_i_clk),
    .D(_00505_),
    .Q(\mem[65][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13861_ (.CLK(clknet_leaf_167_i_clk),
    .D(_00506_),
    .Q(\mem[65][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13862_ (.CLK(clknet_leaf_170_i_clk),
    .D(_00507_),
    .Q(\mem[65][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13863_ (.CLK(clknet_leaf_178_i_clk),
    .D(_00508_),
    .Q(\mem[65][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13864_ (.CLK(clknet_leaf_170_i_clk),
    .D(_00509_),
    .Q(\mem[65][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13865_ (.CLK(clknet_leaf_176_i_clk),
    .D(_00510_),
    .Q(\mem[65][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13866_ (.CLK(clknet_leaf_170_i_clk),
    .D(_00511_),
    .Q(\mem[65][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13867_ (.CLK(clknet_leaf_176_i_clk),
    .D(_00512_),
    .Q(\mem[65][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13868_ (.CLK(clknet_leaf_195_i_clk),
    .D(_00513_),
    .Q(\mem[66][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13869_ (.CLK(clknet_leaf_168_i_clk),
    .D(_00514_),
    .Q(\mem[66][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13870_ (.CLK(clknet_leaf_198_i_clk),
    .D(_00515_),
    .Q(\mem[66][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13871_ (.CLK(clknet_leaf_166_i_clk),
    .D(_00516_),
    .Q(\mem[66][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13872_ (.CLK(clknet_leaf_166_i_clk),
    .D(_00517_),
    .Q(\mem[66][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13873_ (.CLK(clknet_leaf_168_i_clk),
    .D(_00518_),
    .Q(\mem[66][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13874_ (.CLK(clknet_leaf_168_i_clk),
    .D(_00519_),
    .Q(\mem[66][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13875_ (.CLK(clknet_leaf_166_i_clk),
    .D(_00520_),
    .Q(\mem[66][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13876_ (.CLK(clknet_leaf_166_i_clk),
    .D(_00521_),
    .Q(\mem[66][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13877_ (.CLK(clknet_leaf_167_i_clk),
    .D(_00522_),
    .Q(\mem[66][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13878_ (.CLK(clknet_leaf_168_i_clk),
    .D(_00523_),
    .Q(\mem[66][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13879_ (.CLK(clknet_leaf_177_i_clk),
    .D(_00524_),
    .Q(\mem[66][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13880_ (.CLK(clknet_leaf_169_i_clk),
    .D(_00525_),
    .Q(\mem[66][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13881_ (.CLK(clknet_leaf_177_i_clk),
    .D(_00526_),
    .Q(\mem[66][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13882_ (.CLK(clknet_leaf_169_i_clk),
    .D(_00527_),
    .Q(\mem[66][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13883_ (.CLK(clknet_leaf_177_i_clk),
    .D(_00528_),
    .Q(\mem[66][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13884_ (.CLK(clknet_leaf_167_i_clk),
    .D(_00529_),
    .Q(\mem[67][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13885_ (.CLK(clknet_leaf_167_i_clk),
    .D(_00530_),
    .Q(\mem[67][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13886_ (.CLK(clknet_leaf_166_i_clk),
    .D(_00531_),
    .Q(\mem[67][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13887_ (.CLK(clknet_leaf_166_i_clk),
    .D(_00532_),
    .Q(\mem[67][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13888_ (.CLK(clknet_leaf_165_i_clk),
    .D(_00533_),
    .Q(\mem[67][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13889_ (.CLK(clknet_leaf_168_i_clk),
    .D(_00534_),
    .Q(\mem[67][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13890_ (.CLK(clknet_leaf_169_i_clk),
    .D(_00535_),
    .Q(\mem[67][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13891_ (.CLK(clknet_leaf_165_i_clk),
    .D(_00536_),
    .Q(\mem[67][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13892_ (.CLK(clknet_leaf_165_i_clk),
    .D(_00537_),
    .Q(\mem[67][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13893_ (.CLK(clknet_leaf_164_i_clk),
    .D(_00538_),
    .Q(\mem[67][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13894_ (.CLK(clknet_leaf_170_i_clk),
    .D(_00539_),
    .Q(\mem[67][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13895_ (.CLK(clknet_leaf_178_i_clk),
    .D(_00540_),
    .Q(\mem[67][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13896_ (.CLK(clknet_leaf_170_i_clk),
    .D(_00541_),
    .Q(\mem[67][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13897_ (.CLK(clknet_leaf_176_i_clk),
    .D(_00542_),
    .Q(\mem[67][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13898_ (.CLK(clknet_leaf_170_i_clk),
    .D(_00543_),
    .Q(\mem[67][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13899_ (.CLK(clknet_leaf_176_i_clk),
    .D(_00544_),
    .Q(\mem[67][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13900_ (.CLK(clknet_leaf_142_i_clk),
    .D(_00545_),
    .Q(\mem[68][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13901_ (.CLK(clknet_leaf_160_i_clk),
    .D(_00546_),
    .Q(\mem[68][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13902_ (.CLK(clknet_leaf_151_i_clk),
    .D(_00547_),
    .Q(\mem[68][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13903_ (.CLK(clknet_leaf_151_i_clk),
    .D(_00548_),
    .Q(\mem[68][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13904_ (.CLK(clknet_leaf_154_i_clk),
    .D(_00549_),
    .Q(\mem[68][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13905_ (.CLK(clknet_leaf_171_i_clk),
    .D(_00550_),
    .Q(\mem[68][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13906_ (.CLK(clknet_leaf_172_i_clk),
    .D(_00551_),
    .Q(\mem[68][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13907_ (.CLK(clknet_leaf_155_i_clk),
    .D(_00552_),
    .Q(\mem[68][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13908_ (.CLK(clknet_leaf_154_i_clk),
    .D(_00553_),
    .Q(\mem[68][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13909_ (.CLK(clknet_leaf_154_i_clk),
    .D(_00554_),
    .Q(\mem[68][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13910_ (.CLK(clknet_leaf_157_i_clk),
    .D(_00555_),
    .Q(\mem[68][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13911_ (.CLK(clknet_leaf_174_i_clk),
    .D(_00556_),
    .Q(\mem[68][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13912_ (.CLK(clknet_leaf_140_i_clk),
    .D(_00557_),
    .Q(\mem[68][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13913_ (.CLK(clknet_leaf_173_i_clk),
    .D(_00558_),
    .Q(\mem[68][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13914_ (.CLK(clknet_leaf_140_i_clk),
    .D(_00559_),
    .Q(\mem[68][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13915_ (.CLK(clknet_leaf_140_i_clk),
    .D(_00560_),
    .Q(\mem[68][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13916_ (.CLK(clknet_leaf_160_i_clk),
    .D(_00561_),
    .Q(\mem[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13917_ (.CLK(clknet_leaf_164_i_clk),
    .D(_00562_),
    .Q(\mem[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13918_ (.CLK(clknet_leaf_162_i_clk),
    .D(_00563_),
    .Q(\mem[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13919_ (.CLK(clknet_leaf_162_i_clk),
    .D(_00564_),
    .Q(\mem[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13920_ (.CLK(clknet_leaf_162_i_clk),
    .D(_00565_),
    .Q(\mem[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13921_ (.CLK(clknet_leaf_164_i_clk),
    .D(_00566_),
    .Q(\mem[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13922_ (.CLK(clknet_leaf_160_i_clk),
    .D(_00567_),
    .Q(\mem[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13923_ (.CLK(clknet_leaf_162_i_clk),
    .D(_00568_),
    .Q(\mem[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13924_ (.CLK(clknet_leaf_162_i_clk),
    .D(_00569_),
    .Q(\mem[6][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13925_ (.CLK(clknet_leaf_161_i_clk),
    .D(_00570_),
    .Q(\mem[6][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13926_ (.CLK(clknet_leaf_159_i_clk),
    .D(_00571_),
    .Q(\mem[6][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13927_ (.CLK(clknet_leaf_173_i_clk),
    .D(_00572_),
    .Q(\mem[6][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13928_ (.CLK(clknet_leaf_157_i_clk),
    .D(_00573_),
    .Q(\mem[6][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13929_ (.CLK(clknet_leaf_173_i_clk),
    .D(_00574_),
    .Q(\mem[6][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13930_ (.CLK(clknet_leaf_140_i_clk),
    .D(_00575_),
    .Q(\mem[6][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13931_ (.CLK(clknet_leaf_139_i_clk),
    .D(_00576_),
    .Q(\mem[6][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13932_ (.CLK(clknet_leaf_156_i_clk),
    .D(_00577_),
    .Q(\mem[70][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13933_ (.CLK(clknet_leaf_160_i_clk),
    .D(_00578_),
    .Q(\mem[70][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13934_ (.CLK(clknet_leaf_155_i_clk),
    .D(_00579_),
    .Q(\mem[70][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13935_ (.CLK(clknet_leaf_155_i_clk),
    .D(_00580_),
    .Q(\mem[70][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13936_ (.CLK(clknet_leaf_154_i_clk),
    .D(_00581_),
    .Q(\mem[70][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13937_ (.CLK(clknet_leaf_171_i_clk),
    .D(_00582_),
    .Q(\mem[70][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13938_ (.CLK(clknet_leaf_171_i_clk),
    .D(_00583_),
    .Q(\mem[70][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13939_ (.CLK(clknet_leaf_151_i_clk),
    .D(_00584_),
    .Q(\mem[70][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13940_ (.CLK(clknet_leaf_153_i_clk),
    .D(_00585_),
    .Q(\mem[70][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13941_ (.CLK(clknet_leaf_154_i_clk),
    .D(_00586_),
    .Q(\mem[70][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13942_ (.CLK(clknet_leaf_157_i_clk),
    .D(_00587_),
    .Q(\mem[70][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13943_ (.CLK(clknet_leaf_174_i_clk),
    .D(_00588_),
    .Q(\mem[70][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13944_ (.CLK(clknet_leaf_157_i_clk),
    .D(_00589_),
    .Q(\mem[70][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13945_ (.CLK(clknet_leaf_172_i_clk),
    .D(_00590_),
    .Q(\mem[70][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13946_ (.CLK(clknet_leaf_140_i_clk),
    .D(_00591_),
    .Q(\mem[70][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13947_ (.CLK(clknet_leaf_139_i_clk),
    .D(_00592_),
    .Q(\mem[70][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13948_ (.CLK(clknet_leaf_156_i_clk),
    .D(_00593_),
    .Q(\mem[71][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13949_ (.CLK(clknet_leaf_171_i_clk),
    .D(_00594_),
    .Q(\mem[71][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13950_ (.CLK(clknet_leaf_155_i_clk),
    .D(_00595_),
    .Q(\mem[71][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13951_ (.CLK(clknet_leaf_156_i_clk),
    .D(_00596_),
    .Q(\mem[71][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13952_ (.CLK(clknet_leaf_156_i_clk),
    .D(_00597_),
    .Q(\mem[71][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13953_ (.CLK(clknet_leaf_171_i_clk),
    .D(_00598_),
    .Q(\mem[71][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13954_ (.CLK(clknet_leaf_172_i_clk),
    .D(_00599_),
    .Q(\mem[71][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13955_ (.CLK(clknet_leaf_156_i_clk),
    .D(_00600_),
    .Q(\mem[71][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13956_ (.CLK(clknet_leaf_156_i_clk),
    .D(_00601_),
    .Q(\mem[71][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13957_ (.CLK(clknet_leaf_156_i_clk),
    .D(_00602_),
    .Q(\mem[71][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13958_ (.CLK(clknet_leaf_140_i_clk),
    .D(_00603_),
    .Q(\mem[71][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13959_ (.CLK(clknet_leaf_122_i_clk),
    .D(_00604_),
    .Q(\mem[71][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13960_ (.CLK(clknet_leaf_141_i_clk),
    .D(_00605_),
    .Q(\mem[71][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13961_ (.CLK(clknet_leaf_139_i_clk),
    .D(_00606_),
    .Q(\mem[71][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13962_ (.CLK(clknet_leaf_140_i_clk),
    .D(_00607_),
    .Q(\mem[71][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13963_ (.CLK(clknet_leaf_139_i_clk),
    .D(_00608_),
    .Q(\mem[71][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13964_ (.CLK(clknet_leaf_151_i_clk),
    .D(_00609_),
    .Q(\mem[72][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13965_ (.CLK(clknet_leaf_164_i_clk),
    .D(_00610_),
    .Q(\mem[72][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13966_ (.CLK(clknet_leaf_151_i_clk),
    .D(_00611_),
    .Q(\mem[72][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13967_ (.CLK(clknet_leaf_150_i_clk),
    .D(_00612_),
    .Q(\mem[72][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13968_ (.CLK(clknet_leaf_153_i_clk),
    .D(_00613_),
    .Q(\mem[72][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13969_ (.CLK(clknet_leaf_171_i_clk),
    .D(_00614_),
    .Q(\mem[72][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13970_ (.CLK(clknet_leaf_171_i_clk),
    .D(_00615_),
    .Q(\mem[72][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13971_ (.CLK(clknet_leaf_152_i_clk),
    .D(_00616_),
    .Q(\mem[72][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13972_ (.CLK(clknet_leaf_153_i_clk),
    .D(_00617_),
    .Q(\mem[72][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13973_ (.CLK(clknet_leaf_153_i_clk),
    .D(_00618_),
    .Q(\mem[72][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13974_ (.CLK(clknet_leaf_159_i_clk),
    .D(_00619_),
    .Q(\mem[72][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13975_ (.CLK(clknet_leaf_175_i_clk),
    .D(_00620_),
    .Q(\mem[72][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13976_ (.CLK(clknet_leaf_159_i_clk),
    .D(_00621_),
    .Q(\mem[72][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13977_ (.CLK(clknet_leaf_170_i_clk),
    .D(_00622_),
    .Q(\mem[72][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13978_ (.CLK(clknet_leaf_172_i_clk),
    .D(_00623_),
    .Q(\mem[72][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13979_ (.CLK(clknet_leaf_173_i_clk),
    .D(_00624_),
    .Q(\mem[72][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13980_ (.CLK(clknet_leaf_151_i_clk),
    .D(_00625_),
    .Q(\mem[73][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13981_ (.CLK(clknet_leaf_165_i_clk),
    .D(_00626_),
    .Q(\mem[73][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13982_ (.CLK(clknet_leaf_152_i_clk),
    .D(_00627_),
    .Q(\mem[73][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13983_ (.CLK(clknet_leaf_152_i_clk),
    .D(_00628_),
    .Q(\mem[73][3] ));
 sky130_fd_sc_hd__dfxtp_1 _13984_ (.CLK(clknet_leaf_153_i_clk),
    .D(_00629_),
    .Q(\mem[73][4] ));
 sky130_fd_sc_hd__dfxtp_1 _13985_ (.CLK(clknet_leaf_164_i_clk),
    .D(_00630_),
    .Q(\mem[73][5] ));
 sky130_fd_sc_hd__dfxtp_1 _13986_ (.CLK(clknet_leaf_171_i_clk),
    .D(_00631_),
    .Q(\mem[73][6] ));
 sky130_fd_sc_hd__dfxtp_1 _13987_ (.CLK(clknet_leaf_152_i_clk),
    .D(_00632_),
    .Q(\mem[73][7] ));
 sky130_fd_sc_hd__dfxtp_1 _13988_ (.CLK(clknet_leaf_153_i_clk),
    .D(_00633_),
    .Q(\mem[73][8] ));
 sky130_fd_sc_hd__dfxtp_1 _13989_ (.CLK(clknet_leaf_161_i_clk),
    .D(_00634_),
    .Q(\mem[73][9] ));
 sky130_fd_sc_hd__dfxtp_1 _13990_ (.CLK(clknet_leaf_159_i_clk),
    .D(_00635_),
    .Q(\mem[73][10] ));
 sky130_fd_sc_hd__dfxtp_1 _13991_ (.CLK(clknet_leaf_176_i_clk),
    .D(_00636_),
    .Q(\mem[73][11] ));
 sky130_fd_sc_hd__dfxtp_1 _13992_ (.CLK(clknet_leaf_159_i_clk),
    .D(_00637_),
    .Q(\mem[73][12] ));
 sky130_fd_sc_hd__dfxtp_1 _13993_ (.CLK(clknet_leaf_170_i_clk),
    .D(_00638_),
    .Q(\mem[73][13] ));
 sky130_fd_sc_hd__dfxtp_1 _13994_ (.CLK(clknet_leaf_172_i_clk),
    .D(_00639_),
    .Q(\mem[73][14] ));
 sky130_fd_sc_hd__dfxtp_1 _13995_ (.CLK(clknet_leaf_172_i_clk),
    .D(_00640_),
    .Q(\mem[73][15] ));
 sky130_fd_sc_hd__dfxtp_1 _13996_ (.CLK(clknet_leaf_151_i_clk),
    .D(_00641_),
    .Q(\mem[74][0] ));
 sky130_fd_sc_hd__dfxtp_1 _13997_ (.CLK(clknet_leaf_165_i_clk),
    .D(_00642_),
    .Q(\mem[74][1] ));
 sky130_fd_sc_hd__dfxtp_1 _13998_ (.CLK(clknet_leaf_150_i_clk),
    .D(_00643_),
    .Q(\mem[74][2] ));
 sky130_fd_sc_hd__dfxtp_1 _13999_ (.CLK(clknet_leaf_150_i_clk),
    .D(_00644_),
    .Q(\mem[74][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14000_ (.CLK(clknet_leaf_153_i_clk),
    .D(_00645_),
    .Q(\mem[74][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14001_ (.CLK(clknet_leaf_164_i_clk),
    .D(_00646_),
    .Q(\mem[74][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14002_ (.CLK(clknet_leaf_171_i_clk),
    .D(_00647_),
    .Q(\mem[74][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14003_ (.CLK(clknet_leaf_152_i_clk),
    .D(_00648_),
    .Q(\mem[74][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14004_ (.CLK(clknet_leaf_153_i_clk),
    .D(_00649_),
    .Q(\mem[74][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14005_ (.CLK(clknet_leaf_161_i_clk),
    .D(_00650_),
    .Q(\mem[74][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14006_ (.CLK(clknet_leaf_157_i_clk),
    .D(_00651_),
    .Q(\mem[74][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14007_ (.CLK(clknet_leaf_173_i_clk),
    .D(_00652_),
    .Q(\mem[74][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14008_ (.CLK(clknet_leaf_157_i_clk),
    .D(_00653_),
    .Q(\mem[74][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14009_ (.CLK(clknet_leaf_172_i_clk),
    .D(_00654_),
    .Q(\mem[74][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14010_ (.CLK(clknet_leaf_158_i_clk),
    .D(_00655_),
    .Q(\mem[74][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14011_ (.CLK(clknet_leaf_158_i_clk),
    .D(_00656_),
    .Q(\mem[74][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14012_ (.CLK(clknet_leaf_151_i_clk),
    .D(_00657_),
    .Q(\mem[75][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14013_ (.CLK(clknet_leaf_165_i_clk),
    .D(_00658_),
    .Q(\mem[75][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14014_ (.CLK(clknet_leaf_152_i_clk),
    .D(_00659_),
    .Q(\mem[75][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14015_ (.CLK(clknet_leaf_152_i_clk),
    .D(_00660_),
    .Q(\mem[75][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14016_ (.CLK(clknet_leaf_153_i_clk),
    .D(_00661_),
    .Q(\mem[75][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14017_ (.CLK(clknet_leaf_165_i_clk),
    .D(_00662_),
    .Q(\mem[75][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14018_ (.CLK(clknet_leaf_164_i_clk),
    .D(_00663_),
    .Q(\mem[75][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14019_ (.CLK(clknet_leaf_152_i_clk),
    .D(_00664_),
    .Q(\mem[75][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14020_ (.CLK(clknet_leaf_161_i_clk),
    .D(_00665_),
    .Q(\mem[75][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14021_ (.CLK(clknet_leaf_161_i_clk),
    .D(_00666_),
    .Q(\mem[75][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14022_ (.CLK(clknet_leaf_161_i_clk),
    .D(_00667_),
    .Q(\mem[75][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14023_ (.CLK(clknet_leaf_174_i_clk),
    .D(_00668_),
    .Q(\mem[75][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14024_ (.CLK(clknet_leaf_159_i_clk),
    .D(_00669_),
    .Q(\mem[75][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14025_ (.CLK(clknet_leaf_171_i_clk),
    .D(_00670_),
    .Q(\mem[75][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14026_ (.CLK(clknet_leaf_159_i_clk),
    .D(_00671_),
    .Q(\mem[75][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14027_ (.CLK(clknet_leaf_173_i_clk),
    .D(_00672_),
    .Q(\mem[75][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14028_ (.CLK(clknet_leaf_203_i_clk),
    .D(_00673_),
    .Q(\mem[76][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14029_ (.CLK(clknet_leaf_196_i_clk),
    .D(_00674_),
    .Q(\mem[76][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14030_ (.CLK(clknet_leaf_203_i_clk),
    .D(_00675_),
    .Q(\mem[76][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14031_ (.CLK(clknet_leaf_204_i_clk),
    .D(_00676_),
    .Q(\mem[76][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14032_ (.CLK(clknet_leaf_200_i_clk),
    .D(_00677_),
    .Q(\mem[76][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14033_ (.CLK(clknet_leaf_196_i_clk),
    .D(_00678_),
    .Q(\mem[76][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14034_ (.CLK(clknet_leaf_192_i_clk),
    .D(_00679_),
    .Q(\mem[76][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14035_ (.CLK(clknet_leaf_202_i_clk),
    .D(_00680_),
    .Q(\mem[76][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14036_ (.CLK(clknet_leaf_201_i_clk),
    .D(_00681_),
    .Q(\mem[76][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14037_ (.CLK(clknet_leaf_197_i_clk),
    .D(_00682_),
    .Q(\mem[76][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14038_ (.CLK(clknet_leaf_196_i_clk),
    .D(_00683_),
    .Q(\mem[76][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14039_ (.CLK(clknet_leaf_184_i_clk),
    .D(_00684_),
    .Q(\mem[76][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14040_ (.CLK(clknet_leaf_193_i_clk),
    .D(_00685_),
    .Q(\mem[76][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14041_ (.CLK(clknet_leaf_185_i_clk),
    .D(_00686_),
    .Q(\mem[76][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14042_ (.CLK(clknet_leaf_193_i_clk),
    .D(_00687_),
    .Q(\mem[76][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14043_ (.CLK(clknet_leaf_186_i_clk),
    .D(_00688_),
    .Q(\mem[76][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14044_ (.CLK(clknet_leaf_200_i_clk),
    .D(_00689_),
    .Q(\mem[77][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14045_ (.CLK(clknet_leaf_197_i_clk),
    .D(_00690_),
    .Q(\mem[77][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14046_ (.CLK(clknet_leaf_198_i_clk),
    .D(_00691_),
    .Q(\mem[77][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14047_ (.CLK(clknet_leaf_199_i_clk),
    .D(_00692_),
    .Q(\mem[77][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14048_ (.CLK(clknet_leaf_200_i_clk),
    .D(_00693_),
    .Q(\mem[77][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14049_ (.CLK(clknet_leaf_195_i_clk),
    .D(_00694_),
    .Q(\mem[77][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14050_ (.CLK(clknet_leaf_192_i_clk),
    .D(_00695_),
    .Q(\mem[77][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14051_ (.CLK(clknet_leaf_200_i_clk),
    .D(_00696_),
    .Q(\mem[77][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14052_ (.CLK(clknet_leaf_199_i_clk),
    .D(_00697_),
    .Q(\mem[77][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14053_ (.CLK(clknet_leaf_197_i_clk),
    .D(_00698_),
    .Q(\mem[77][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14054_ (.CLK(clknet_leaf_194_i_clk),
    .D(_00699_),
    .Q(\mem[77][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14055_ (.CLK(clknet_leaf_184_i_clk),
    .D(_00700_),
    .Q(\mem[77][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14056_ (.CLK(clknet_leaf_194_i_clk),
    .D(_00701_),
    .Q(\mem[77][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14057_ (.CLK(clknet_leaf_185_i_clk),
    .D(_00702_),
    .Q(\mem[77][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14058_ (.CLK(clknet_leaf_194_i_clk),
    .D(_00703_),
    .Q(\mem[77][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14059_ (.CLK(clknet_leaf_184_i_clk),
    .D(_00704_),
    .Q(\mem[77][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14060_ (.CLK(clknet_leaf_201_i_clk),
    .D(_00705_),
    .Q(\mem[78][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14061_ (.CLK(clknet_leaf_197_i_clk),
    .D(_00706_),
    .Q(\mem[78][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14062_ (.CLK(clknet_leaf_201_i_clk),
    .D(_00707_),
    .Q(\mem[78][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14063_ (.CLK(clknet_leaf_201_i_clk),
    .D(_00708_),
    .Q(\mem[78][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14064_ (.CLK(clknet_leaf_200_i_clk),
    .D(_00709_),
    .Q(\mem[78][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14065_ (.CLK(clknet_leaf_195_i_clk),
    .D(_00710_),
    .Q(\mem[78][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14066_ (.CLK(clknet_leaf_196_i_clk),
    .D(_00711_),
    .Q(\mem[78][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14067_ (.CLK(clknet_leaf_200_i_clk),
    .D(_00712_),
    .Q(\mem[78][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14068_ (.CLK(clknet_leaf_201_i_clk),
    .D(_00713_),
    .Q(\mem[78][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14069_ (.CLK(clknet_leaf_197_i_clk),
    .D(_00714_),
    .Q(\mem[78][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14070_ (.CLK(clknet_leaf_195_i_clk),
    .D(_00715_),
    .Q(\mem[78][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14071_ (.CLK(clknet_leaf_184_i_clk),
    .D(_00716_),
    .Q(\mem[78][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14072_ (.CLK(clknet_leaf_194_i_clk),
    .D(_00717_),
    .Q(\mem[78][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14073_ (.CLK(clknet_leaf_185_i_clk),
    .D(_00718_),
    .Q(\mem[78][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14074_ (.CLK(clknet_leaf_194_i_clk),
    .D(_00719_),
    .Q(\mem[78][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14075_ (.CLK(clknet_leaf_185_i_clk),
    .D(_00720_),
    .Q(\mem[78][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14076_ (.CLK(clknet_leaf_160_i_clk),
    .D(_00721_),
    .Q(\mem[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14077_ (.CLK(clknet_leaf_163_i_clk),
    .D(_00722_),
    .Q(\mem[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14078_ (.CLK(clknet_leaf_162_i_clk),
    .D(_00723_),
    .Q(\mem[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14079_ (.CLK(clknet_leaf_163_i_clk),
    .D(_00724_),
    .Q(\mem[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14080_ (.CLK(clknet_leaf_162_i_clk),
    .D(_00725_),
    .Q(\mem[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14081_ (.CLK(clknet_leaf_163_i_clk),
    .D(_00726_),
    .Q(\mem[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14082_ (.CLK(clknet_leaf_159_i_clk),
    .D(_00727_),
    .Q(\mem[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14083_ (.CLK(clknet_leaf_161_i_clk),
    .D(_00728_),
    .Q(\mem[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14084_ (.CLK(clknet_leaf_162_i_clk),
    .D(_00729_),
    .Q(\mem[7][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14085_ (.CLK(clknet_leaf_161_i_clk),
    .D(_00730_),
    .Q(\mem[7][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14086_ (.CLK(clknet_leaf_159_i_clk),
    .D(_00731_),
    .Q(\mem[7][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14087_ (.CLK(clknet_leaf_173_i_clk),
    .D(_00732_),
    .Q(\mem[7][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14088_ (.CLK(clknet_leaf_157_i_clk),
    .D(_00733_),
    .Q(\mem[7][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14089_ (.CLK(clknet_leaf_173_i_clk),
    .D(_00734_),
    .Q(\mem[7][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14090_ (.CLK(clknet_leaf_157_i_clk),
    .D(_00735_),
    .Q(\mem[7][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14091_ (.CLK(clknet_leaf_121_i_clk),
    .D(_00736_),
    .Q(\mem[7][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14092_ (.CLK(clknet_leaf_221_i_clk),
    .D(_00737_),
    .Q(\mem[80][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14093_ (.CLK(clknet_leaf_203_i_clk),
    .D(_00738_),
    .Q(\mem[80][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14094_ (.CLK(clknet_leaf_216_i_clk),
    .D(_00739_),
    .Q(\mem[80][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14095_ (.CLK(clknet_leaf_220_i_clk),
    .D(_00740_),
    .Q(\mem[80][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14096_ (.CLK(clknet_leaf_216_i_clk),
    .D(_00741_),
    .Q(\mem[80][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14097_ (.CLK(clknet_leaf_192_i_clk),
    .D(_00742_),
    .Q(\mem[80][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14098_ (.CLK(clknet_leaf_191_i_clk),
    .D(_00743_),
    .Q(\mem[80][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14099_ (.CLK(clknet_leaf_210_i_clk),
    .D(_00744_),
    .Q(\mem[80][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14100_ (.CLK(clknet_leaf_211_i_clk),
    .D(_00745_),
    .Q(\mem[80][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14101_ (.CLK(clknet_leaf_211_i_clk),
    .D(_00746_),
    .Q(\mem[80][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14102_ (.CLK(clknet_leaf_193_i_clk),
    .D(_00747_),
    .Q(\mem[80][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14103_ (.CLK(clknet_leaf_183_i_clk),
    .D(_00748_),
    .Q(\mem[80][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14104_ (.CLK(clknet_leaf_193_i_clk),
    .D(_00749_),
    .Q(\mem[80][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14105_ (.CLK(clknet_leaf_186_i_clk),
    .D(_00750_),
    .Q(\mem[80][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14106_ (.CLK(clknet_leaf_193_i_clk),
    .D(_00751_),
    .Q(\mem[80][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14107_ (.CLK(clknet_leaf_186_i_clk),
    .D(_00752_),
    .Q(\mem[80][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14108_ (.CLK(clknet_leaf_222_i_clk),
    .D(_00753_),
    .Q(\mem[81][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14109_ (.CLK(clknet_leaf_207_i_clk),
    .D(_00754_),
    .Q(\mem[81][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14110_ (.CLK(clknet_leaf_223_i_clk),
    .D(_00755_),
    .Q(\mem[81][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14111_ (.CLK(clknet_leaf_221_i_clk),
    .D(_00756_),
    .Q(\mem[81][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14112_ (.CLK(clknet_leaf_221_i_clk),
    .D(_00757_),
    .Q(\mem[81][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14113_ (.CLK(clknet_leaf_191_i_clk),
    .D(_00758_),
    .Q(\mem[81][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14114_ (.CLK(clknet_leaf_191_i_clk),
    .D(_00759_),
    .Q(\mem[81][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14115_ (.CLK(clknet_leaf_225_i_clk),
    .D(_00760_),
    .Q(\mem[81][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14116_ (.CLK(clknet_leaf_210_i_clk),
    .D(_00761_),
    .Q(\mem[81][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14117_ (.CLK(clknet_leaf_210_i_clk),
    .D(_00762_),
    .Q(\mem[81][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14118_ (.CLK(clknet_leaf_227_i_clk),
    .D(_00763_),
    .Q(\mem[81][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14119_ (.CLK(clknet_leaf_187_i_clk),
    .D(_00764_),
    .Q(\mem[81][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14120_ (.CLK(clknet_leaf_227_i_clk),
    .D(_00765_),
    .Q(\mem[81][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14121_ (.CLK(clknet_leaf_188_i_clk),
    .D(_00766_),
    .Q(\mem[81][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14122_ (.CLK(clknet_leaf_190_i_clk),
    .D(_00767_),
    .Q(\mem[81][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14123_ (.CLK(clknet_leaf_189_i_clk),
    .D(_00768_),
    .Q(\mem[81][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14124_ (.CLK(clknet_leaf_222_i_clk),
    .D(_00769_),
    .Q(\mem[82][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14125_ (.CLK(clknet_leaf_191_i_clk),
    .D(_00770_),
    .Q(\mem[82][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14126_ (.CLK(clknet_leaf_222_i_clk),
    .D(_00771_),
    .Q(\mem[82][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14127_ (.CLK(clknet_leaf_221_i_clk),
    .D(_00772_),
    .Q(\mem[82][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14128_ (.CLK(clknet_leaf_221_i_clk),
    .D(_00773_),
    .Q(\mem[82][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14129_ (.CLK(clknet_leaf_191_i_clk),
    .D(_00774_),
    .Q(\mem[82][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14130_ (.CLK(clknet_leaf_191_i_clk),
    .D(_00775_),
    .Q(\mem[82][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14131_ (.CLK(clknet_leaf_225_i_clk),
    .D(_00776_),
    .Q(\mem[82][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14132_ (.CLK(clknet_leaf_210_i_clk),
    .D(_00777_),
    .Q(\mem[82][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14133_ (.CLK(clknet_leaf_210_i_clk),
    .D(_00778_),
    .Q(\mem[82][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14134_ (.CLK(clknet_leaf_227_i_clk),
    .D(_00779_),
    .Q(\mem[82][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14135_ (.CLK(clknet_leaf_187_i_clk),
    .D(_00780_),
    .Q(\mem[82][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14136_ (.CLK(clknet_leaf_227_i_clk),
    .D(_00781_),
    .Q(\mem[82][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14137_ (.CLK(clknet_leaf_188_i_clk),
    .D(_00782_),
    .Q(\mem[82][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14138_ (.CLK(clknet_leaf_227_i_clk),
    .D(_00783_),
    .Q(\mem[82][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14139_ (.CLK(clknet_leaf_243_i_clk),
    .D(_00784_),
    .Q(\mem[82][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14140_ (.CLK(clknet_leaf_222_i_clk),
    .D(_00785_),
    .Q(\mem[83][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14141_ (.CLK(clknet_leaf_203_i_clk),
    .D(_00786_),
    .Q(\mem[83][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14142_ (.CLK(clknet_leaf_222_i_clk),
    .D(_00787_),
    .Q(\mem[83][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14143_ (.CLK(clknet_leaf_221_i_clk),
    .D(_00788_),
    .Q(\mem[83][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14144_ (.CLK(clknet_leaf_220_i_clk),
    .D(_00789_),
    .Q(\mem[83][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14145_ (.CLK(clknet_leaf_191_i_clk),
    .D(_00790_),
    .Q(\mem[83][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14146_ (.CLK(clknet_leaf_191_i_clk),
    .D(_00791_),
    .Q(\mem[83][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14147_ (.CLK(clknet_leaf_216_i_clk),
    .D(_00792_),
    .Q(\mem[83][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14148_ (.CLK(clknet_leaf_211_i_clk),
    .D(_00793_),
    .Q(\mem[83][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14149_ (.CLK(clknet_leaf_210_i_clk),
    .D(_00794_),
    .Q(\mem[83][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14150_ (.CLK(clknet_leaf_209_i_clk),
    .D(_00795_),
    .Q(\mem[83][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14151_ (.CLK(clknet_leaf_245_i_clk),
    .D(_00796_),
    .Q(\mem[83][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14152_ (.CLK(clknet_leaf_209_i_clk),
    .D(_00797_),
    .Q(\mem[83][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14153_ (.CLK(clknet_leaf_188_i_clk),
    .D(_00798_),
    .Q(\mem[83][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14154_ (.CLK(clknet_leaf_208_i_clk),
    .D(_00799_),
    .Q(\mem[83][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14155_ (.CLK(clknet_leaf_189_i_clk),
    .D(_00800_),
    .Q(\mem[83][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14156_ (.CLK(clknet_leaf_218_i_clk),
    .D(_00801_),
    .Q(\mem[84][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14157_ (.CLK(clknet_leaf_203_i_clk),
    .D(_00802_),
    .Q(\mem[84][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14158_ (.CLK(clknet_leaf_218_i_clk),
    .D(_00803_),
    .Q(\mem[84][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14159_ (.CLK(clknet_leaf_217_i_clk),
    .D(_00804_),
    .Q(\mem[84][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14160_ (.CLK(clknet_leaf_217_i_clk),
    .D(_00805_),
    .Q(\mem[84][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14161_ (.CLK(clknet_leaf_203_i_clk),
    .D(_00806_),
    .Q(\mem[84][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14162_ (.CLK(clknet_leaf_192_i_clk),
    .D(_00807_),
    .Q(\mem[84][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14163_ (.CLK(clknet_leaf_215_i_clk),
    .D(_00808_),
    .Q(\mem[84][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14164_ (.CLK(clknet_leaf_215_i_clk),
    .D(_00809_),
    .Q(\mem[84][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14165_ (.CLK(clknet_leaf_214_i_clk),
    .D(_00810_),
    .Q(\mem[84][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14166_ (.CLK(clknet_leaf_207_i_clk),
    .D(_00811_),
    .Q(\mem[84][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14167_ (.CLK(clknet_leaf_186_i_clk),
    .D(_00812_),
    .Q(\mem[84][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14168_ (.CLK(clknet_leaf_192_i_clk),
    .D(_00813_),
    .Q(\mem[84][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14169_ (.CLK(clknet_leaf_186_i_clk),
    .D(_00814_),
    .Q(\mem[84][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14170_ (.CLK(clknet_leaf_207_i_clk),
    .D(_00815_),
    .Q(\mem[84][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14171_ (.CLK(clknet_leaf_207_i_clk),
    .D(_00816_),
    .Q(\mem[84][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14172_ (.CLK(clknet_leaf_218_i_clk),
    .D(_00817_),
    .Q(\mem[85][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14173_ (.CLK(clknet_leaf_204_i_clk),
    .D(_00818_),
    .Q(\mem[85][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14174_ (.CLK(clknet_leaf_218_i_clk),
    .D(_00819_),
    .Q(\mem[85][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14175_ (.CLK(clknet_leaf_217_i_clk),
    .D(_00820_),
    .Q(\mem[85][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14176_ (.CLK(clknet_leaf_217_i_clk),
    .D(_00821_),
    .Q(\mem[85][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14177_ (.CLK(clknet_leaf_203_i_clk),
    .D(_00822_),
    .Q(\mem[85][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14178_ (.CLK(clknet_leaf_205_i_clk),
    .D(_00823_),
    .Q(\mem[85][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14179_ (.CLK(clknet_leaf_215_i_clk),
    .D(_00824_),
    .Q(\mem[85][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14180_ (.CLK(clknet_leaf_214_i_clk),
    .D(_00825_),
    .Q(\mem[85][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14181_ (.CLK(clknet_leaf_213_i_clk),
    .D(_00826_),
    .Q(\mem[85][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14182_ (.CLK(clknet_leaf_213_i_clk),
    .D(_00827_),
    .Q(\mem[85][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14183_ (.CLK(clknet_leaf_187_i_clk),
    .D(_00828_),
    .Q(\mem[85][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14184_ (.CLK(clknet_leaf_212_i_clk),
    .D(_00829_),
    .Q(\mem[85][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14185_ (.CLK(clknet_leaf_193_i_clk),
    .D(_00830_),
    .Q(\mem[85][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14186_ (.CLK(clknet_leaf_205_i_clk),
    .D(_00831_),
    .Q(\mem[85][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14187_ (.CLK(clknet_leaf_205_i_clk),
    .D(_00832_),
    .Q(\mem[85][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14188_ (.CLK(clknet_leaf_218_i_clk),
    .D(_00833_),
    .Q(\mem[86][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14189_ (.CLK(clknet_leaf_204_i_clk),
    .D(_00834_),
    .Q(\mem[86][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14190_ (.CLK(clknet_leaf_218_i_clk),
    .D(_00835_),
    .Q(\mem[86][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14191_ (.CLK(clknet_leaf_218_i_clk),
    .D(_00836_),
    .Q(\mem[86][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14192_ (.CLK(clknet_leaf_217_i_clk),
    .D(_00837_),
    .Q(\mem[86][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14193_ (.CLK(clknet_leaf_204_i_clk),
    .D(_00838_),
    .Q(\mem[86][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14194_ (.CLK(clknet_leaf_205_i_clk),
    .D(_00839_),
    .Q(\mem[86][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14195_ (.CLK(clknet_leaf_215_i_clk),
    .D(_00840_),
    .Q(\mem[86][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14196_ (.CLK(clknet_leaf_214_i_clk),
    .D(_00841_),
    .Q(\mem[86][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14197_ (.CLK(clknet_leaf_213_i_clk),
    .D(_00842_),
    .Q(\mem[86][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14198_ (.CLK(clknet_leaf_213_i_clk),
    .D(_00843_),
    .Q(\mem[86][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14199_ (.CLK(clknet_leaf_186_i_clk),
    .D(_00844_),
    .Q(\mem[86][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14200_ (.CLK(clknet_leaf_204_i_clk),
    .D(_00845_),
    .Q(\mem[86][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14201_ (.CLK(clknet_leaf_193_i_clk),
    .D(_00846_),
    .Q(\mem[86][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14202_ (.CLK(clknet_leaf_205_i_clk),
    .D(_00847_),
    .Q(\mem[86][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14203_ (.CLK(clknet_leaf_205_i_clk),
    .D(_00848_),
    .Q(\mem[86][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14204_ (.CLK(clknet_leaf_218_i_clk),
    .D(_00849_),
    .Q(\mem[87][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14205_ (.CLK(clknet_leaf_204_i_clk),
    .D(_00850_),
    .Q(\mem[87][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14206_ (.CLK(clknet_leaf_218_i_clk),
    .D(_00851_),
    .Q(\mem[87][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14207_ (.CLK(clknet_leaf_217_i_clk),
    .D(_00852_),
    .Q(\mem[87][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14208_ (.CLK(clknet_leaf_217_i_clk),
    .D(_00853_),
    .Q(\mem[87][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14209_ (.CLK(clknet_leaf_204_i_clk),
    .D(_00854_),
    .Q(\mem[87][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14210_ (.CLK(clknet_leaf_205_i_clk),
    .D(_00855_),
    .Q(\mem[87][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14211_ (.CLK(clknet_leaf_215_i_clk),
    .D(_00856_),
    .Q(\mem[87][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14212_ (.CLK(clknet_leaf_214_i_clk),
    .D(_00857_),
    .Q(\mem[87][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14213_ (.CLK(clknet_leaf_213_i_clk),
    .D(_00858_),
    .Q(\mem[87][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14214_ (.CLK(clknet_leaf_205_i_clk),
    .D(_00859_),
    .Q(\mem[87][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14215_ (.CLK(clknet_leaf_186_i_clk),
    .D(_00860_),
    .Q(\mem[87][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14216_ (.CLK(clknet_leaf_203_i_clk),
    .D(_00861_),
    .Q(\mem[87][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14217_ (.CLK(clknet_leaf_193_i_clk),
    .D(_00862_),
    .Q(\mem[87][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14218_ (.CLK(clknet_leaf_205_i_clk),
    .D(_00863_),
    .Q(\mem[87][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14219_ (.CLK(clknet_leaf_205_i_clk),
    .D(_00864_),
    .Q(\mem[87][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14220_ (.CLK(clknet_leaf_219_i_clk),
    .D(_00865_),
    .Q(\mem[88][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14221_ (.CLK(clknet_leaf_206_i_clk),
    .D(_00866_),
    .Q(\mem[88][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14222_ (.CLK(clknet_leaf_219_i_clk),
    .D(_00867_),
    .Q(\mem[88][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14223_ (.CLK(clknet_leaf_222_i_clk),
    .D(_00868_),
    .Q(\mem[88][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14224_ (.CLK(clknet_leaf_220_i_clk),
    .D(_00869_),
    .Q(\mem[88][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14225_ (.CLK(clknet_leaf_206_i_clk),
    .D(_00870_),
    .Q(\mem[88][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14226_ (.CLK(clknet_leaf_208_i_clk),
    .D(_00871_),
    .Q(\mem[88][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14227_ (.CLK(clknet_leaf_216_i_clk),
    .D(_00872_),
    .Q(\mem[88][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14228_ (.CLK(clknet_leaf_215_i_clk),
    .D(_00873_),
    .Q(\mem[88][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14229_ (.CLK(clknet_leaf_211_i_clk),
    .D(_00874_),
    .Q(\mem[88][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14230_ (.CLK(clknet_leaf_210_i_clk),
    .D(_00875_),
    .Q(\mem[88][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14231_ (.CLK(clknet_leaf_188_i_clk),
    .D(_00876_),
    .Q(\mem[88][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14232_ (.CLK(clknet_leaf_209_i_clk),
    .D(_00877_),
    .Q(\mem[88][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14233_ (.CLK(clknet_leaf_188_i_clk),
    .D(_00878_),
    .Q(\mem[88][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14234_ (.CLK(clknet_leaf_208_i_clk),
    .D(_00879_),
    .Q(\mem[88][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14235_ (.CLK(clknet_leaf_208_i_clk),
    .D(_00880_),
    .Q(\mem[88][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14236_ (.CLK(clknet_leaf_178_i_clk),
    .D(_00881_),
    .Q(\mem[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14237_ (.CLK(clknet_leaf_115_i_clk),
    .D(_00882_),
    .Q(\mem[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14238_ (.CLK(clknet_leaf_179_i_clk),
    .D(_00883_),
    .Q(\mem[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14239_ (.CLK(clknet_leaf_115_i_clk),
    .D(_00884_),
    .Q(\mem[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14240_ (.CLK(clknet_leaf_115_i_clk),
    .D(_00885_),
    .Q(\mem[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14241_ (.CLK(clknet_leaf_114_i_clk),
    .D(_00886_),
    .Q(\mem[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14242_ (.CLK(clknet_leaf_118_i_clk),
    .D(_00887_),
    .Q(\mem[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14243_ (.CLK(clknet_leaf_115_i_clk),
    .D(_00888_),
    .Q(\mem[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14244_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00889_),
    .Q(\mem[8][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14245_ (.CLK(clknet_leaf_119_i_clk),
    .D(_00890_),
    .Q(\mem[8][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14246_ (.CLK(clknet_leaf_175_i_clk),
    .D(_00891_),
    .Q(\mem[8][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14247_ (.CLK(clknet_leaf_175_i_clk),
    .D(_00892_),
    .Q(\mem[8][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14248_ (.CLK(clknet_leaf_175_i_clk),
    .D(_00893_),
    .Q(\mem[8][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14249_ (.CLK(clknet_leaf_175_i_clk),
    .D(_00894_),
    .Q(\mem[8][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14250_ (.CLK(clknet_leaf_176_i_clk),
    .D(_00895_),
    .Q(\mem[8][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14251_ (.CLK(clknet_leaf_176_i_clk),
    .D(_00896_),
    .Q(\mem[8][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14252_ (.CLK(clknet_leaf_219_i_clk),
    .D(_00897_),
    .Q(\mem[90][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14253_ (.CLK(clknet_leaf_207_i_clk),
    .D(_00898_),
    .Q(\mem[90][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14254_ (.CLK(clknet_leaf_219_i_clk),
    .D(_00899_),
    .Q(\mem[90][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14255_ (.CLK(clknet_leaf_220_i_clk),
    .D(_00900_),
    .Q(\mem[90][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14256_ (.CLK(clknet_leaf_220_i_clk),
    .D(_00901_),
    .Q(\mem[90][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14257_ (.CLK(clknet_leaf_207_i_clk),
    .D(_00902_),
    .Q(\mem[90][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14258_ (.CLK(clknet_leaf_207_i_clk),
    .D(_00903_),
    .Q(\mem[90][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14259_ (.CLK(clknet_leaf_216_i_clk),
    .D(_00904_),
    .Q(\mem[90][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14260_ (.CLK(clknet_leaf_215_i_clk),
    .D(_00905_),
    .Q(\mem[90][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14261_ (.CLK(clknet_leaf_212_i_clk),
    .D(_00906_),
    .Q(\mem[90][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14262_ (.CLK(clknet_leaf_209_i_clk),
    .D(_00907_),
    .Q(\mem[90][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14263_ (.CLK(clknet_leaf_189_i_clk),
    .D(_00908_),
    .Q(\mem[90][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14264_ (.CLK(clknet_leaf_209_i_clk),
    .D(_00909_),
    .Q(\mem[90][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14265_ (.CLK(clknet_leaf_188_i_clk),
    .D(_00910_),
    .Q(\mem[90][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14266_ (.CLK(clknet_leaf_208_i_clk),
    .D(_00911_),
    .Q(\mem[90][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14267_ (.CLK(clknet_leaf_208_i_clk),
    .D(_00912_),
    .Q(\mem[90][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14268_ (.CLK(clknet_leaf_219_i_clk),
    .D(_00913_),
    .Q(\mem[91][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14269_ (.CLK(clknet_leaf_204_i_clk),
    .D(_00914_),
    .Q(\mem[91][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14270_ (.CLK(clknet_leaf_218_i_clk),
    .D(_00915_),
    .Q(\mem[91][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14271_ (.CLK(clknet_leaf_220_i_clk),
    .D(_00916_),
    .Q(\mem[91][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14272_ (.CLK(clknet_leaf_217_i_clk),
    .D(_00917_),
    .Q(\mem[91][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14273_ (.CLK(clknet_leaf_206_i_clk),
    .D(_00918_),
    .Q(\mem[91][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14274_ (.CLK(clknet_leaf_206_i_clk),
    .D(_00919_),
    .Q(\mem[91][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14275_ (.CLK(clknet_leaf_215_i_clk),
    .D(_00920_),
    .Q(\mem[91][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14276_ (.CLK(clknet_leaf_212_i_clk),
    .D(_00921_),
    .Q(\mem[91][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14277_ (.CLK(clknet_leaf_212_i_clk),
    .D(_00922_),
    .Q(\mem[91][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14278_ (.CLK(clknet_leaf_211_i_clk),
    .D(_00923_),
    .Q(\mem[91][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14279_ (.CLK(clknet_leaf_244_i_clk),
    .D(_00924_),
    .Q(\mem[91][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14280_ (.CLK(clknet_leaf_211_i_clk),
    .D(_00925_),
    .Q(\mem[91][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14281_ (.CLK(clknet_leaf_186_i_clk),
    .D(_00926_),
    .Q(\mem[91][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14282_ (.CLK(clknet_leaf_206_i_clk),
    .D(_00927_),
    .Q(\mem[91][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14283_ (.CLK(clknet_leaf_206_i_clk),
    .D(_00928_),
    .Q(\mem[91][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14284_ (.CLK(clknet_leaf_230_i_clk),
    .D(_00929_),
    .Q(\mem[92][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14285_ (.CLK(clknet_leaf_190_i_clk),
    .D(_00930_),
    .Q(\mem[92][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14286_ (.CLK(clknet_leaf_230_i_clk),
    .D(_00931_),
    .Q(\mem[92][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14287_ (.CLK(clknet_leaf_224_i_clk),
    .D(_00932_),
    .Q(\mem[92][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14288_ (.CLK(clknet_leaf_230_i_clk),
    .D(_00933_),
    .Q(\mem[92][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14289_ (.CLK(clknet_leaf_190_i_clk),
    .D(_00934_),
    .Q(\mem[92][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14290_ (.CLK(clknet_leaf_242_i_clk),
    .D(_00935_),
    .Q(\mem[92][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14291_ (.CLK(clknet_leaf_226_i_clk),
    .D(_00936_),
    .Q(\mem[92][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14292_ (.CLK(clknet_leaf_226_i_clk),
    .D(_00937_),
    .Q(\mem[92][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14293_ (.CLK(clknet_leaf_226_i_clk),
    .D(_00938_),
    .Q(\mem[92][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14294_ (.CLK(clknet_leaf_244_i_clk),
    .D(_00939_),
    .Q(\mem[92][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14295_ (.CLK(clknet_leaf_245_i_clk),
    .D(_00940_),
    .Q(\mem[92][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14296_ (.CLK(clknet_leaf_244_i_clk),
    .D(_00941_),
    .Q(\mem[92][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14297_ (.CLK(clknet_leaf_183_i_clk),
    .D(_00942_),
    .Q(\mem[92][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14298_ (.CLK(clknet_leaf_244_i_clk),
    .D(_00943_),
    .Q(\mem[92][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14299_ (.CLK(clknet_leaf_244_i_clk),
    .D(_00944_),
    .Q(\mem[92][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14300_ (.CLK(clknet_leaf_224_i_clk),
    .D(_00945_),
    .Q(\mem[93][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14301_ (.CLK(clknet_leaf_191_i_clk),
    .D(_00946_),
    .Q(\mem[93][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14302_ (.CLK(clknet_leaf_224_i_clk),
    .D(_00947_),
    .Q(\mem[93][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14303_ (.CLK(clknet_leaf_224_i_clk),
    .D(_00948_),
    .Q(\mem[93][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14304_ (.CLK(clknet_leaf_225_i_clk),
    .D(_00949_),
    .Q(\mem[93][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14305_ (.CLK(clknet_leaf_191_i_clk),
    .D(_00950_),
    .Q(\mem[93][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14306_ (.CLK(clknet_leaf_188_i_clk),
    .D(_00951_),
    .Q(\mem[93][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14307_ (.CLK(clknet_leaf_225_i_clk),
    .D(_00952_),
    .Q(\mem[93][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14308_ (.CLK(clknet_leaf_225_i_clk),
    .D(_00953_),
    .Q(\mem[93][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14309_ (.CLK(clknet_leaf_226_i_clk),
    .D(_00954_),
    .Q(\mem[93][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14310_ (.CLK(clknet_leaf_243_i_clk),
    .D(_00955_),
    .Q(\mem[93][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14311_ (.CLK(clknet_leaf_245_i_clk),
    .D(_00956_),
    .Q(\mem[93][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14312_ (.CLK(clknet_leaf_243_i_clk),
    .D(_00957_),
    .Q(\mem[93][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14313_ (.CLK(clknet_leaf_187_i_clk),
    .D(_00958_),
    .Q(\mem[93][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14314_ (.CLK(clknet_leaf_243_i_clk),
    .D(_00959_),
    .Q(\mem[93][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14315_ (.CLK(clknet_leaf_243_i_clk),
    .D(_00960_),
    .Q(\mem[93][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14316_ (.CLK(clknet_leaf_221_i_clk),
    .D(_00961_),
    .Q(\mem[94][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14317_ (.CLK(clknet_leaf_208_i_clk),
    .D(_00962_),
    .Q(\mem[94][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14318_ (.CLK(clknet_leaf_223_i_clk),
    .D(_00963_),
    .Q(\mem[94][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14319_ (.CLK(clknet_leaf_224_i_clk),
    .D(_00964_),
    .Q(\mem[94][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14320_ (.CLK(clknet_leaf_224_i_clk),
    .D(_00965_),
    .Q(\mem[94][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14321_ (.CLK(clknet_leaf_190_i_clk),
    .D(_00966_),
    .Q(\mem[94][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14322_ (.CLK(clknet_leaf_227_i_clk),
    .D(_00967_),
    .Q(\mem[94][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14323_ (.CLK(clknet_leaf_226_i_clk),
    .D(_00968_),
    .Q(\mem[94][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14324_ (.CLK(clknet_leaf_225_i_clk),
    .D(_00969_),
    .Q(\mem[94][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14325_ (.CLK(clknet_leaf_226_i_clk),
    .D(_00970_),
    .Q(\mem[94][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14326_ (.CLK(clknet_leaf_242_i_clk),
    .D(_00971_),
    .Q(\mem[94][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14327_ (.CLK(clknet_leaf_244_i_clk),
    .D(_00972_),
    .Q(\mem[94][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14328_ (.CLK(clknet_leaf_242_i_clk),
    .D(_00973_),
    .Q(\mem[94][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14329_ (.CLK(clknet_leaf_187_i_clk),
    .D(_00974_),
    .Q(\mem[94][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14330_ (.CLK(clknet_leaf_243_i_clk),
    .D(_00975_),
    .Q(\mem[94][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14331_ (.CLK(clknet_leaf_244_i_clk),
    .D(_00976_),
    .Q(\mem[94][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14332_ (.CLK(clknet_leaf_224_i_clk),
    .D(_00977_),
    .Q(\mem[95][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14333_ (.CLK(clknet_leaf_208_i_clk),
    .D(_00978_),
    .Q(\mem[95][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14334_ (.CLK(clknet_leaf_224_i_clk),
    .D(_00979_),
    .Q(\mem[95][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14335_ (.CLK(clknet_leaf_224_i_clk),
    .D(_00980_),
    .Q(\mem[95][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14336_ (.CLK(clknet_leaf_224_i_clk),
    .D(_00981_),
    .Q(\mem[95][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14337_ (.CLK(clknet_leaf_208_i_clk),
    .D(_00982_),
    .Q(\mem[95][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14338_ (.CLK(clknet_leaf_227_i_clk),
    .D(_00983_),
    .Q(\mem[95][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14339_ (.CLK(clknet_leaf_226_i_clk),
    .D(_00984_),
    .Q(\mem[95][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14340_ (.CLK(clknet_leaf_226_i_clk),
    .D(_00985_),
    .Q(\mem[95][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14341_ (.CLK(clknet_leaf_226_i_clk),
    .D(_00986_),
    .Q(\mem[95][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14342_ (.CLK(clknet_leaf_242_i_clk),
    .D(_00987_),
    .Q(\mem[95][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14343_ (.CLK(clknet_leaf_245_i_clk),
    .D(_00988_),
    .Q(\mem[95][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14344_ (.CLK(clknet_leaf_242_i_clk),
    .D(_00989_),
    .Q(\mem[95][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14345_ (.CLK(clknet_leaf_183_i_clk),
    .D(_00990_),
    .Q(\mem[95][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14346_ (.CLK(clknet_leaf_243_i_clk),
    .D(_00991_),
    .Q(\mem[95][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14347_ (.CLK(clknet_leaf_244_i_clk),
    .D(_00992_),
    .Q(\mem[95][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14348_ (.CLK(clknet_leaf_284_i_clk),
    .D(_00993_),
    .Q(\mem[96][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14349_ (.CLK(clknet_leaf_259_i_clk),
    .D(_00994_),
    .Q(\mem[96][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14350_ (.CLK(clknet_leaf_285_i_clk),
    .D(_00995_),
    .Q(\mem[96][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14351_ (.CLK(clknet_leaf_285_i_clk),
    .D(_00996_),
    .Q(\mem[96][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14352_ (.CLK(clknet_leaf_275_i_clk),
    .D(_00997_),
    .Q(\mem[96][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14353_ (.CLK(clknet_leaf_259_i_clk),
    .D(_00998_),
    .Q(\mem[96][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14354_ (.CLK(clknet_leaf_261_i_clk),
    .D(_00999_),
    .Q(\mem[96][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14355_ (.CLK(clknet_leaf_276_i_clk),
    .D(_01000_),
    .Q(\mem[96][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14356_ (.CLK(clknet_leaf_274_i_clk),
    .D(_01001_),
    .Q(\mem[96][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14357_ (.CLK(clknet_leaf_275_i_clk),
    .D(_01002_),
    .Q(\mem[96][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14358_ (.CLK(clknet_leaf_280_i_clk),
    .D(_01003_),
    .Q(\mem[96][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14359_ (.CLK(clknet_leaf_30_i_clk),
    .D(_01004_),
    .Q(\mem[96][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14360_ (.CLK(clknet_leaf_262_i_clk),
    .D(_01005_),
    .Q(\mem[96][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14361_ (.CLK(clknet_leaf_30_i_clk),
    .D(_01006_),
    .Q(\mem[96][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14362_ (.CLK(clknet_leaf_8_i_clk),
    .D(_01007_),
    .Q(\mem[96][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14363_ (.CLK(clknet_leaf_29_i_clk),
    .D(_01008_),
    .Q(\mem[96][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14364_ (.CLK(clknet_leaf_284_i_clk),
    .D(_01009_),
    .Q(\mem[97][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14365_ (.CLK(clknet_leaf_261_i_clk),
    .D(_01010_),
    .Q(\mem[97][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14366_ (.CLK(clknet_leaf_285_i_clk),
    .D(_01011_),
    .Q(\mem[97][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14367_ (.CLK(clknet_leaf_285_i_clk),
    .D(_01012_),
    .Q(\mem[97][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14368_ (.CLK(clknet_leaf_277_i_clk),
    .D(_01013_),
    .Q(\mem[97][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14369_ (.CLK(clknet_leaf_259_i_clk),
    .D(_01014_),
    .Q(\mem[97][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14370_ (.CLK(clknet_leaf_261_i_clk),
    .D(_01015_),
    .Q(\mem[97][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14371_ (.CLK(clknet_leaf_277_i_clk),
    .D(_01016_),
    .Q(\mem[97][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14372_ (.CLK(clknet_leaf_275_i_clk),
    .D(_01017_),
    .Q(\mem[97][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14373_ (.CLK(clknet_leaf_276_i_clk),
    .D(_01018_),
    .Q(\mem[97][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14374_ (.CLK(clknet_leaf_280_i_clk),
    .D(_01019_),
    .Q(\mem[97][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14375_ (.CLK(clknet_leaf_29_i_clk),
    .D(_01020_),
    .Q(\mem[97][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14376_ (.CLK(clknet_leaf_262_i_clk),
    .D(_01021_),
    .Q(\mem[97][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14377_ (.CLK(clknet_leaf_30_i_clk),
    .D(_01022_),
    .Q(\mem[97][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14378_ (.CLK(clknet_leaf_280_i_clk),
    .D(_01023_),
    .Q(\mem[97][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14379_ (.CLK(clknet_leaf_28_i_clk),
    .D(_01024_),
    .Q(\mem[97][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14380_ (.CLK(clknet_leaf_285_i_clk),
    .D(_01025_),
    .Q(\mem[98][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14381_ (.CLK(clknet_leaf_261_i_clk),
    .D(_01026_),
    .Q(\mem[98][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14382_ (.CLK(clknet_leaf_285_i_clk),
    .D(_01027_),
    .Q(\mem[98][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14383_ (.CLK(clknet_leaf_284_i_clk),
    .D(_01028_),
    .Q(\mem[98][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14384_ (.CLK(clknet_leaf_276_i_clk),
    .D(_01029_),
    .Q(\mem[98][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14385_ (.CLK(clknet_leaf_259_i_clk),
    .D(_01030_),
    .Q(\mem[98][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14386_ (.CLK(clknet_leaf_261_i_clk),
    .D(_01031_),
    .Q(\mem[98][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14387_ (.CLK(clknet_leaf_276_i_clk),
    .D(_01032_),
    .Q(\mem[98][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14388_ (.CLK(clknet_leaf_275_i_clk),
    .D(_01033_),
    .Q(\mem[98][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14389_ (.CLK(clknet_leaf_276_i_clk),
    .D(_01034_),
    .Q(\mem[98][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14390_ (.CLK(clknet_leaf_280_i_clk),
    .D(_01035_),
    .Q(\mem[98][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14391_ (.CLK(clknet_leaf_29_i_clk),
    .D(_01036_),
    .Q(\mem[98][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14392_ (.CLK(clknet_leaf_280_i_clk),
    .D(_01037_),
    .Q(\mem[98][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14393_ (.CLK(clknet_leaf_30_i_clk),
    .D(_01038_),
    .Q(\mem[98][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14394_ (.CLK(clknet_leaf_7_i_clk),
    .D(_01039_),
    .Q(\mem[98][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14395_ (.CLK(clknet_leaf_28_i_clk),
    .D(_01040_),
    .Q(\mem[98][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14396_ (.CLK(clknet_leaf_252_i_clk),
    .D(_01041_),
    .Q(\mem[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14397_ (.CLK(clknet_leaf_252_i_clk),
    .D(_01042_),
    .Q(\mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14398_ (.CLK(clknet_leaf_249_i_clk),
    .D(_01043_),
    .Q(\mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14399_ (.CLK(clknet_leaf_257_i_clk),
    .D(_01044_),
    .Q(\mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14400_ (.CLK(clknet_leaf_253_i_clk),
    .D(_01045_),
    .Q(\mem[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14401_ (.CLK(clknet_leaf_38_i_clk),
    .D(_01046_),
    .Q(\mem[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14402_ (.CLK(clknet_leaf_257_i_clk),
    .D(_01047_),
    .Q(\mem[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14403_ (.CLK(clknet_leaf_253_i_clk),
    .D(_01048_),
    .Q(\mem[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14404_ (.CLK(clknet_leaf_253_i_clk),
    .D(_01049_),
    .Q(\mem[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14405_ (.CLK(clknet_leaf_252_i_clk),
    .D(_01050_),
    .Q(\mem[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14406_ (.CLK(clknet_leaf_251_i_clk),
    .D(_01051_),
    .Q(\mem[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14407_ (.CLK(clknet_leaf_182_i_clk),
    .D(_01052_),
    .Q(\mem[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14408_ (.CLK(clknet_leaf_182_i_clk),
    .D(_01053_),
    .Q(\mem[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14409_ (.CLK(clknet_leaf_181_i_clk),
    .D(_01054_),
    .Q(\mem[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14410_ (.CLK(clknet_leaf_182_i_clk),
    .D(_01055_),
    .Q(\mem[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14411_ (.CLK(clknet_leaf_182_i_clk),
    .D(_01056_),
    .Q(\mem[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14412_ (.CLK(clknet_leaf_284_i_clk),
    .D(_01057_),
    .Q(\mem[100][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14413_ (.CLK(clknet_leaf_263_i_clk),
    .D(_01058_),
    .Q(\mem[100][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14414_ (.CLK(clknet_leaf_283_i_clk),
    .D(_01059_),
    .Q(\mem[100][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14415_ (.CLK(clknet_leaf_277_i_clk),
    .D(_01060_),
    .Q(\mem[100][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14416_ (.CLK(clknet_leaf_277_i_clk),
    .D(_01061_),
    .Q(\mem[100][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14417_ (.CLK(clknet_leaf_265_i_clk),
    .D(_01062_),
    .Q(\mem[100][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14418_ (.CLK(clknet_leaf_261_i_clk),
    .D(_01063_),
    .Q(\mem[100][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14419_ (.CLK(clknet_leaf_279_i_clk),
    .D(_01064_),
    .Q(\mem[100][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14420_ (.CLK(clknet_leaf_278_i_clk),
    .D(_01065_),
    .Q(\mem[100][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14421_ (.CLK(clknet_leaf_279_i_clk),
    .D(_01066_),
    .Q(\mem[100][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14422_ (.CLK(clknet_leaf_279_i_clk),
    .D(_01067_),
    .Q(\mem[100][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14423_ (.CLK(clknet_leaf_260_i_clk),
    .D(_01068_),
    .Q(\mem[100][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14424_ (.CLK(clknet_leaf_263_i_clk),
    .D(_01069_),
    .Q(\mem[100][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14425_ (.CLK(clknet_leaf_31_i_clk),
    .D(_01070_),
    .Q(\mem[100][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14426_ (.CLK(clknet_leaf_262_i_clk),
    .D(_01071_),
    .Q(\mem[100][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14427_ (.CLK(clknet_leaf_29_i_clk),
    .D(_01072_),
    .Q(\mem[100][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14428_ (.CLK(clknet_leaf_283_i_clk),
    .D(_01073_),
    .Q(\mem[101][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14429_ (.CLK(clknet_leaf_263_i_clk),
    .D(_01074_),
    .Q(\mem[101][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14430_ (.CLK(clknet_leaf_281_i_clk),
    .D(_01075_),
    .Q(\mem[101][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14431_ (.CLK(clknet_leaf_284_i_clk),
    .D(_01076_),
    .Q(\mem[101][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14432_ (.CLK(clknet_leaf_278_i_clk),
    .D(_01077_),
    .Q(\mem[101][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14433_ (.CLK(clknet_leaf_265_i_clk),
    .D(_01078_),
    .Q(\mem[101][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14434_ (.CLK(clknet_leaf_263_i_clk),
    .D(_01079_),
    .Q(\mem[101][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14435_ (.CLK(clknet_leaf_279_i_clk),
    .D(_01080_),
    .Q(\mem[101][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14436_ (.CLK(clknet_leaf_279_i_clk),
    .D(_01081_),
    .Q(\mem[101][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14437_ (.CLK(clknet_leaf_281_i_clk),
    .D(_01082_),
    .Q(\mem[101][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14438_ (.CLK(clknet_leaf_279_i_clk),
    .D(_01083_),
    .Q(\mem[101][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14439_ (.CLK(clknet_leaf_31_i_clk),
    .D(_01084_),
    .Q(\mem[101][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14440_ (.CLK(clknet_leaf_279_i_clk),
    .D(_01085_),
    .Q(\mem[101][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14441_ (.CLK(clknet_leaf_32_i_clk),
    .D(_01086_),
    .Q(\mem[101][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14442_ (.CLK(clknet_leaf_262_i_clk),
    .D(_01087_),
    .Q(\mem[101][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14443_ (.CLK(clknet_leaf_29_i_clk),
    .D(_01088_),
    .Q(\mem[101][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14444_ (.CLK(clknet_leaf_283_i_clk),
    .D(_01089_),
    .Q(\mem[102][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14445_ (.CLK(clknet_leaf_263_i_clk),
    .D(_01090_),
    .Q(\mem[102][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14446_ (.CLK(clknet_leaf_281_i_clk),
    .D(_01091_),
    .Q(\mem[102][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14447_ (.CLK(clknet_leaf_284_i_clk),
    .D(_01092_),
    .Q(\mem[102][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14448_ (.CLK(clknet_leaf_277_i_clk),
    .D(_01093_),
    .Q(\mem[102][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14449_ (.CLK(clknet_leaf_265_i_clk),
    .D(_01094_),
    .Q(\mem[102][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14450_ (.CLK(clknet_leaf_262_i_clk),
    .D(_01095_),
    .Q(\mem[102][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14451_ (.CLK(clknet_leaf_281_i_clk),
    .D(_01096_),
    .Q(\mem[102][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14452_ (.CLK(clknet_leaf_279_i_clk),
    .D(_01097_),
    .Q(\mem[102][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14453_ (.CLK(clknet_leaf_281_i_clk),
    .D(_01098_),
    .Q(\mem[102][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14454_ (.CLK(clknet_leaf_280_i_clk),
    .D(_01099_),
    .Q(\mem[102][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14455_ (.CLK(clknet_leaf_31_i_clk),
    .D(_01100_),
    .Q(\mem[102][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14456_ (.CLK(clknet_leaf_262_i_clk),
    .D(_01101_),
    .Q(\mem[102][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14457_ (.CLK(clknet_leaf_31_i_clk),
    .D(_01102_),
    .Q(\mem[102][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14458_ (.CLK(clknet_leaf_262_i_clk),
    .D(_01103_),
    .Q(\mem[102][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14459_ (.CLK(clknet_leaf_28_i_clk),
    .D(_01104_),
    .Q(\mem[102][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14460_ (.CLK(clknet_leaf_283_i_clk),
    .D(_01105_),
    .Q(\mem[103][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14461_ (.CLK(clknet_leaf_263_i_clk),
    .D(_01106_),
    .Q(\mem[103][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14462_ (.CLK(clknet_leaf_281_i_clk),
    .D(_01107_),
    .Q(\mem[103][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14463_ (.CLK(clknet_leaf_284_i_clk),
    .D(_01108_),
    .Q(\mem[103][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14464_ (.CLK(clknet_leaf_277_i_clk),
    .D(_01109_),
    .Q(\mem[103][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14465_ (.CLK(clknet_leaf_265_i_clk),
    .D(_01110_),
    .Q(\mem[103][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14466_ (.CLK(clknet_leaf_262_i_clk),
    .D(_01111_),
    .Q(\mem[103][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14467_ (.CLK(clknet_leaf_281_i_clk),
    .D(_01112_),
    .Q(\mem[103][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14468_ (.CLK(clknet_leaf_279_i_clk),
    .D(_01113_),
    .Q(\mem[103][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14469_ (.CLK(clknet_leaf_281_i_clk),
    .D(_01114_),
    .Q(\mem[103][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14470_ (.CLK(clknet_leaf_279_i_clk),
    .D(_01115_),
    .Q(\mem[103][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14471_ (.CLK(clknet_leaf_261_i_clk),
    .D(_01116_),
    .Q(\mem[103][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14472_ (.CLK(clknet_leaf_279_i_clk),
    .D(_01117_),
    .Q(\mem[103][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14473_ (.CLK(clknet_leaf_32_i_clk),
    .D(_01118_),
    .Q(\mem[103][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14474_ (.CLK(clknet_leaf_262_i_clk),
    .D(_01119_),
    .Q(\mem[103][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14475_ (.CLK(clknet_leaf_29_i_clk),
    .D(_01120_),
    .Q(\mem[103][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14476_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01121_),
    .Q(\mem[104][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14477_ (.CLK(clknet_leaf_36_i_clk),
    .D(_01122_),
    .Q(\mem[104][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14478_ (.CLK(clknet_leaf_32_i_clk),
    .D(_01123_),
    .Q(\mem[104][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14479_ (.CLK(clknet_leaf_32_i_clk),
    .D(_01124_),
    .Q(\mem[104][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14480_ (.CLK(clknet_leaf_32_i_clk),
    .D(_01125_),
    .Q(\mem[104][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14481_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01126_),
    .Q(\mem[104][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14482_ (.CLK(clknet_leaf_35_i_clk),
    .D(_01127_),
    .Q(\mem[104][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14483_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01128_),
    .Q(\mem[104][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14484_ (.CLK(clknet_leaf_35_i_clk),
    .D(_01129_),
    .Q(\mem[104][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14485_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01130_),
    .Q(\mem[104][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14486_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01131_),
    .Q(\mem[104][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14487_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01132_),
    .Q(\mem[104][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14488_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01133_),
    .Q(\mem[104][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14489_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01134_),
    .Q(\mem[104][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14490_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01135_),
    .Q(\mem[104][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14491_ (.CLK(clknet_leaf_40_i_clk),
    .D(_01136_),
    .Q(\mem[104][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14492_ (.CLK(clknet_leaf_23_i_clk),
    .D(_01137_),
    .Q(\mem[105][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14493_ (.CLK(clknet_leaf_36_i_clk),
    .D(_01138_),
    .Q(\mem[105][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14494_ (.CLK(clknet_leaf_24_i_clk),
    .D(_01139_),
    .Q(\mem[105][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14495_ (.CLK(clknet_leaf_33_i_clk),
    .D(_01140_),
    .Q(\mem[105][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14496_ (.CLK(clknet_leaf_32_i_clk),
    .D(_01141_),
    .Q(\mem[105][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14497_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01142_),
    .Q(\mem[105][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14498_ (.CLK(clknet_leaf_35_i_clk),
    .D(_01143_),
    .Q(\mem[105][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14499_ (.CLK(clknet_leaf_23_i_clk),
    .D(_01144_),
    .Q(\mem[105][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14500_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01145_),
    .Q(\mem[105][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14501_ (.CLK(clknet_leaf_33_i_clk),
    .D(_01146_),
    .Q(\mem[105][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14502_ (.CLK(clknet_leaf_44_i_clk),
    .D(_01147_),
    .Q(\mem[105][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14503_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01148_),
    .Q(\mem[105][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14504_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01149_),
    .Q(\mem[105][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14505_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01150_),
    .Q(\mem[105][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14506_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01151_),
    .Q(\mem[105][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14507_ (.CLK(clknet_leaf_43_i_clk),
    .D(_01152_),
    .Q(\mem[105][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14508_ (.CLK(clknet_leaf_24_i_clk),
    .D(_01153_),
    .Q(\mem[106][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14509_ (.CLK(clknet_leaf_35_i_clk),
    .D(_01154_),
    .Q(\mem[106][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14510_ (.CLK(clknet_leaf_25_i_clk),
    .D(_01155_),
    .Q(\mem[106][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14511_ (.CLK(clknet_leaf_24_i_clk),
    .D(_01156_),
    .Q(\mem[106][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14512_ (.CLK(clknet_leaf_33_i_clk),
    .D(_01157_),
    .Q(\mem[106][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14513_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01158_),
    .Q(\mem[106][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14514_ (.CLK(clknet_leaf_35_i_clk),
    .D(_01159_),
    .Q(\mem[106][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14515_ (.CLK(clknet_leaf_23_i_clk),
    .D(_01160_),
    .Q(\mem[106][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14516_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01161_),
    .Q(\mem[106][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14517_ (.CLK(clknet_leaf_24_i_clk),
    .D(_01162_),
    .Q(\mem[106][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14518_ (.CLK(clknet_leaf_43_i_clk),
    .D(_01163_),
    .Q(\mem[106][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14519_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01164_),
    .Q(\mem[106][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14520_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01165_),
    .Q(\mem[106][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14521_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01166_),
    .Q(\mem[106][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14522_ (.CLK(clknet_leaf_43_i_clk),
    .D(_01167_),
    .Q(\mem[106][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14523_ (.CLK(clknet_leaf_53_i_clk),
    .D(_01168_),
    .Q(\mem[106][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14524_ (.CLK(clknet_leaf_22_i_clk),
    .D(_01169_),
    .Q(\mem[107][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14525_ (.CLK(clknet_leaf_36_i_clk),
    .D(_01170_),
    .Q(\mem[107][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14526_ (.CLK(clknet_leaf_25_i_clk),
    .D(_01171_),
    .Q(\mem[107][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14527_ (.CLK(clknet_leaf_25_i_clk),
    .D(_01172_),
    .Q(\mem[107][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14528_ (.CLK(clknet_leaf_33_i_clk),
    .D(_01173_),
    .Q(\mem[107][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14529_ (.CLK(clknet_leaf_37_i_clk),
    .D(_01174_),
    .Q(\mem[107][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14530_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01175_),
    .Q(\mem[107][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14531_ (.CLK(clknet_leaf_23_i_clk),
    .D(_01176_),
    .Q(\mem[107][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14532_ (.CLK(clknet_leaf_34_i_clk),
    .D(_01177_),
    .Q(\mem[107][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14533_ (.CLK(clknet_leaf_23_i_clk),
    .D(_01178_),
    .Q(\mem[107][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14534_ (.CLK(clknet_leaf_44_i_clk),
    .D(_01179_),
    .Q(\mem[107][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14535_ (.CLK(clknet_leaf_35_i_clk),
    .D(_01180_),
    .Q(\mem[107][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14536_ (.CLK(clknet_leaf_44_i_clk),
    .D(_01181_),
    .Q(\mem[107][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14537_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01182_),
    .Q(\mem[107][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14538_ (.CLK(clknet_leaf_42_i_clk),
    .D(_01183_),
    .Q(\mem[107][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14539_ (.CLK(clknet_leaf_43_i_clk),
    .D(_01184_),
    .Q(\mem[107][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14540_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01185_),
    .Q(\mem[108][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14541_ (.CLK(clknet_leaf_110_i_clk),
    .D(_01186_),
    .Q(\mem[108][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14542_ (.CLK(clknet_leaf_51_i_clk),
    .D(_01187_),
    .Q(\mem[108][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14543_ (.CLK(clknet_leaf_52_i_clk),
    .D(_01188_),
    .Q(\mem[108][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14544_ (.CLK(clknet_leaf_45_i_clk),
    .D(_01189_),
    .Q(\mem[108][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14545_ (.CLK(clknet_leaf_110_i_clk),
    .D(_01190_),
    .Q(\mem[108][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14546_ (.CLK(clknet_leaf_52_i_clk),
    .D(_01191_),
    .Q(\mem[108][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14547_ (.CLK(clknet_leaf_45_i_clk),
    .D(_01192_),
    .Q(\mem[108][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14548_ (.CLK(clknet_leaf_45_i_clk),
    .D(_01193_),
    .Q(\mem[108][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14549_ (.CLK(clknet_leaf_50_i_clk),
    .D(_01194_),
    .Q(\mem[108][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14550_ (.CLK(clknet_leaf_46_i_clk),
    .D(_01195_),
    .Q(\mem[108][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14551_ (.CLK(clknet_leaf_46_i_clk),
    .D(_01196_),
    .Q(\mem[108][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14552_ (.CLK(clknet_leaf_47_i_clk),
    .D(_01197_),
    .Q(\mem[108][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14553_ (.CLK(clknet_leaf_106_i_clk),
    .D(_01198_),
    .Q(\mem[108][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14554_ (.CLK(clknet_leaf_105_i_clk),
    .D(_01199_),
    .Q(\mem[108][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14555_ (.CLK(clknet_leaf_47_i_clk),
    .D(_01200_),
    .Q(\mem[108][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14556_ (.CLK(clknet_leaf_179_i_clk),
    .D(_01201_),
    .Q(\mem[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14557_ (.CLK(clknet_leaf_116_i_clk),
    .D(_01202_),
    .Q(\mem[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14558_ (.CLK(clknet_leaf_125_i_clk),
    .D(_01203_),
    .Q(\mem[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14559_ (.CLK(clknet_leaf_125_i_clk),
    .D(_01204_),
    .Q(\mem[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14560_ (.CLK(clknet_leaf_117_i_clk),
    .D(_01205_),
    .Q(\mem[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14561_ (.CLK(clknet_leaf_114_i_clk),
    .D(_01206_),
    .Q(\mem[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14562_ (.CLK(clknet_leaf_125_i_clk),
    .D(_01207_),
    .Q(\mem[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14563_ (.CLK(clknet_leaf_118_i_clk),
    .D(_01208_),
    .Q(\mem[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14564_ (.CLK(clknet_leaf_122_i_clk),
    .D(_01209_),
    .Q(\mem[10][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14565_ (.CLK(clknet_leaf_122_i_clk),
    .D(_01210_),
    .Q(\mem[10][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14566_ (.CLK(clknet_leaf_141_i_clk),
    .D(_01211_),
    .Q(\mem[10][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14567_ (.CLK(clknet_leaf_143_i_clk),
    .D(_01212_),
    .Q(\mem[10][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14568_ (.CLK(clknet_leaf_143_i_clk),
    .D(_01213_),
    .Q(\mem[10][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14569_ (.CLK(clknet_leaf_119_i_clk),
    .D(_01214_),
    .Q(\mem[10][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14570_ (.CLK(clknet_leaf_142_i_clk),
    .D(_01215_),
    .Q(\mem[10][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14571_ (.CLK(clknet_leaf_142_i_clk),
    .D(_01216_),
    .Q(\mem[10][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14572_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01217_),
    .Q(\mem[110][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14573_ (.CLK(clknet_leaf_46_i_clk),
    .D(_01218_),
    .Q(\mem[110][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14574_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01219_),
    .Q(\mem[110][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14575_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01220_),
    .Q(\mem[110][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14576_ (.CLK(clknet_leaf_50_i_clk),
    .D(_01221_),
    .Q(\mem[110][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14577_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01222_),
    .Q(\mem[110][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14578_ (.CLK(clknet_leaf_52_i_clk),
    .D(_01223_),
    .Q(\mem[110][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14579_ (.CLK(clknet_leaf_52_i_clk),
    .D(_01224_),
    .Q(\mem[110][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14580_ (.CLK(clknet_leaf_45_i_clk),
    .D(_01225_),
    .Q(\mem[110][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14581_ (.CLK(clknet_leaf_50_i_clk),
    .D(_01226_),
    .Q(\mem[110][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14582_ (.CLK(clknet_leaf_47_i_clk),
    .D(_01227_),
    .Q(\mem[110][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14583_ (.CLK(clknet_leaf_46_i_clk),
    .D(_01228_),
    .Q(\mem[110][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14584_ (.CLK(clknet_leaf_47_i_clk),
    .D(_01229_),
    .Q(\mem[110][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14585_ (.CLK(clknet_leaf_106_i_clk),
    .D(_01230_),
    .Q(\mem[110][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14586_ (.CLK(clknet_leaf_47_i_clk),
    .D(_01231_),
    .Q(\mem[110][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14587_ (.CLK(clknet_leaf_47_i_clk),
    .D(_01232_),
    .Q(\mem[110][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14588_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01233_),
    .Q(\mem[111][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14589_ (.CLK(clknet_leaf_46_i_clk),
    .D(_01234_),
    .Q(\mem[111][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14590_ (.CLK(clknet_leaf_55_i_clk),
    .D(_01235_),
    .Q(\mem[111][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14591_ (.CLK(clknet_leaf_51_i_clk),
    .D(_01236_),
    .Q(\mem[111][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14592_ (.CLK(clknet_leaf_50_i_clk),
    .D(_01237_),
    .Q(\mem[111][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14593_ (.CLK(clknet_leaf_41_i_clk),
    .D(_01238_),
    .Q(\mem[111][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14594_ (.CLK(clknet_leaf_52_i_clk),
    .D(_01239_),
    .Q(\mem[111][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14595_ (.CLK(clknet_leaf_52_i_clk),
    .D(_01240_),
    .Q(\mem[111][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14596_ (.CLK(clknet_leaf_45_i_clk),
    .D(_01241_),
    .Q(\mem[111][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14597_ (.CLK(clknet_leaf_52_i_clk),
    .D(_01242_),
    .Q(\mem[111][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14598_ (.CLK(clknet_leaf_46_i_clk),
    .D(_01243_),
    .Q(\mem[111][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14599_ (.CLK(clknet_leaf_46_i_clk),
    .D(_01244_),
    .Q(\mem[111][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14600_ (.CLK(clknet_leaf_47_i_clk),
    .D(_01245_),
    .Q(\mem[111][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14601_ (.CLK(clknet_leaf_105_i_clk),
    .D(_01246_),
    .Q(\mem[111][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14602_ (.CLK(clknet_leaf_105_i_clk),
    .D(_01247_),
    .Q(\mem[111][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14603_ (.CLK(clknet_leaf_47_i_clk),
    .D(_01248_),
    .Q(\mem[111][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14604_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01249_),
    .Q(\mem[112][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14605_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01250_),
    .Q(\mem[112][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14606_ (.CLK(clknet_leaf_131_i_clk),
    .D(_01251_),
    .Q(\mem[112][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14607_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01252_),
    .Q(\mem[112][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14608_ (.CLK(clknet_leaf_131_i_clk),
    .D(_01253_),
    .Q(\mem[112][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14609_ (.CLK(clknet_leaf_128_i_clk),
    .D(_01254_),
    .Q(\mem[112][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14610_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01255_),
    .Q(\mem[112][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14611_ (.CLK(clknet_leaf_132_i_clk),
    .D(_01256_),
    .Q(\mem[112][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14612_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01257_),
    .Q(\mem[112][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14613_ (.CLK(clknet_leaf_132_i_clk),
    .D(_01258_),
    .Q(\mem[112][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14614_ (.CLK(clknet_leaf_145_i_clk),
    .D(_01259_),
    .Q(\mem[112][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14615_ (.CLK(clknet_leaf_144_i_clk),
    .D(_01260_),
    .Q(\mem[112][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14616_ (.CLK(clknet_leaf_146_i_clk),
    .D(_01261_),
    .Q(\mem[112][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14617_ (.CLK(clknet_leaf_137_i_clk),
    .D(_01262_),
    .Q(\mem[112][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14618_ (.CLK(clknet_leaf_145_i_clk),
    .D(_01263_),
    .Q(\mem[112][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14619_ (.CLK(clknet_leaf_146_i_clk),
    .D(_01264_),
    .Q(\mem[112][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14620_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01265_),
    .Q(\mem[113][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14621_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01266_),
    .Q(\mem[113][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14622_ (.CLK(clknet_leaf_131_i_clk),
    .D(_01267_),
    .Q(\mem[113][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14623_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01268_),
    .Q(\mem[113][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14624_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01269_),
    .Q(\mem[113][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14625_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01270_),
    .Q(\mem[113][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14626_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01271_),
    .Q(\mem[113][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14627_ (.CLK(clknet_leaf_132_i_clk),
    .D(_01272_),
    .Q(\mem[113][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14628_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01273_),
    .Q(\mem[113][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14629_ (.CLK(clknet_leaf_132_i_clk),
    .D(_01274_),
    .Q(\mem[113][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14630_ (.CLK(clknet_leaf_144_i_clk),
    .D(_01275_),
    .Q(\mem[113][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14631_ (.CLK(clknet_leaf_144_i_clk),
    .D(_01276_),
    .Q(\mem[113][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14632_ (.CLK(clknet_leaf_145_i_clk),
    .D(_01277_),
    .Q(\mem[113][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14633_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01278_),
    .Q(\mem[113][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14634_ (.CLK(clknet_leaf_145_i_clk),
    .D(_01279_),
    .Q(\mem[113][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14635_ (.CLK(clknet_leaf_146_i_clk),
    .D(_01280_),
    .Q(\mem[113][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14636_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01281_),
    .Q(\mem[114][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14637_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01282_),
    .Q(\mem[114][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14638_ (.CLK(clknet_leaf_131_i_clk),
    .D(_01283_),
    .Q(\mem[114][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14639_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01284_),
    .Q(\mem[114][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14640_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01285_),
    .Q(\mem[114][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14641_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01286_),
    .Q(\mem[114][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14642_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01287_),
    .Q(\mem[114][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14643_ (.CLK(clknet_leaf_131_i_clk),
    .D(_01288_),
    .Q(\mem[114][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14644_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01289_),
    .Q(\mem[114][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14645_ (.CLK(clknet_leaf_132_i_clk),
    .D(_01290_),
    .Q(\mem[114][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14646_ (.CLK(clknet_leaf_144_i_clk),
    .D(_01291_),
    .Q(\mem[114][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14647_ (.CLK(clknet_leaf_135_i_clk),
    .D(_01292_),
    .Q(\mem[114][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14648_ (.CLK(clknet_leaf_146_i_clk),
    .D(_01293_),
    .Q(\mem[114][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14649_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01294_),
    .Q(\mem[114][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14650_ (.CLK(clknet_leaf_145_i_clk),
    .D(_01295_),
    .Q(\mem[114][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14651_ (.CLK(clknet_leaf_142_i_clk),
    .D(_01296_),
    .Q(\mem[114][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14652_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01297_),
    .Q(\mem[115][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14653_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01298_),
    .Q(\mem[115][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14654_ (.CLK(clknet_leaf_131_i_clk),
    .D(_01299_),
    .Q(\mem[115][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14655_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01300_),
    .Q(\mem[115][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14656_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01301_),
    .Q(\mem[115][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14657_ (.CLK(clknet_leaf_128_i_clk),
    .D(_01302_),
    .Q(\mem[115][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14658_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01303_),
    .Q(\mem[115][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14659_ (.CLK(clknet_leaf_131_i_clk),
    .D(_01304_),
    .Q(\mem[115][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14660_ (.CLK(clknet_leaf_132_i_clk),
    .D(_01305_),
    .Q(\mem[115][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14661_ (.CLK(clknet_leaf_132_i_clk),
    .D(_01306_),
    .Q(\mem[115][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14662_ (.CLK(clknet_leaf_144_i_clk),
    .D(_01307_),
    .Q(\mem[115][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14663_ (.CLK(clknet_leaf_135_i_clk),
    .D(_01308_),
    .Q(\mem[115][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14664_ (.CLK(clknet_leaf_145_i_clk),
    .D(_01309_),
    .Q(\mem[115][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14665_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01310_),
    .Q(\mem[115][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14666_ (.CLK(clknet_leaf_145_i_clk),
    .D(_01311_),
    .Q(\mem[115][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14667_ (.CLK(clknet_leaf_146_i_clk),
    .D(_01312_),
    .Q(\mem[115][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14668_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01313_),
    .Q(\mem[116][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14669_ (.CLK(clknet_leaf_101_i_clk),
    .D(_01314_),
    .Q(\mem[116][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14670_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01315_),
    .Q(\mem[116][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14671_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01316_),
    .Q(\mem[116][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14672_ (.CLK(clknet_leaf_95_i_clk),
    .D(_01317_),
    .Q(\mem[116][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14673_ (.CLK(clknet_leaf_100_i_clk),
    .D(_01318_),
    .Q(\mem[116][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14674_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01319_),
    .Q(\mem[116][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14675_ (.CLK(clknet_leaf_132_i_clk),
    .D(_01320_),
    .Q(\mem[116][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14676_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01321_),
    .Q(\mem[116][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14677_ (.CLK(clknet_leaf_137_i_clk),
    .D(_01322_),
    .Q(\mem[116][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14678_ (.CLK(clknet_leaf_147_i_clk),
    .D(_01323_),
    .Q(\mem[116][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14679_ (.CLK(clknet_leaf_135_i_clk),
    .D(_01324_),
    .Q(\mem[116][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14680_ (.CLK(clknet_leaf_147_i_clk),
    .D(_01325_),
    .Q(\mem[116][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14681_ (.CLK(clknet_leaf_138_i_clk),
    .D(_01326_),
    .Q(\mem[116][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14682_ (.CLK(clknet_leaf_148_i_clk),
    .D(_01327_),
    .Q(\mem[116][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14683_ (.CLK(clknet_leaf_150_i_clk),
    .D(_01328_),
    .Q(\mem[116][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14684_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01329_),
    .Q(\mem[117][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14685_ (.CLK(clknet_leaf_101_i_clk),
    .D(_01330_),
    .Q(\mem[117][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14686_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01331_),
    .Q(\mem[117][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14687_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01332_),
    .Q(\mem[117][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14688_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01333_),
    .Q(\mem[117][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14689_ (.CLK(clknet_leaf_101_i_clk),
    .D(_01334_),
    .Q(\mem[117][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14690_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01335_),
    .Q(\mem[117][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14691_ (.CLK(clknet_leaf_131_i_clk),
    .D(_01336_),
    .Q(\mem[117][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14692_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01337_),
    .Q(\mem[117][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14693_ (.CLK(clknet_leaf_134_i_clk),
    .D(_01338_),
    .Q(\mem[117][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14694_ (.CLK(clknet_leaf_148_i_clk),
    .D(_01339_),
    .Q(\mem[117][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14695_ (.CLK(clknet_leaf_135_i_clk),
    .D(_01340_),
    .Q(\mem[117][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14696_ (.CLK(clknet_leaf_147_i_clk),
    .D(_01341_),
    .Q(\mem[117][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14697_ (.CLK(clknet_leaf_138_i_clk),
    .D(_01342_),
    .Q(\mem[117][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14698_ (.CLK(clknet_leaf_148_i_clk),
    .D(_01343_),
    .Q(\mem[117][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14699_ (.CLK(clknet_leaf_151_i_clk),
    .D(_01344_),
    .Q(\mem[117][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14700_ (.CLK(clknet_leaf_89_i_clk),
    .D(_01345_),
    .Q(\mem[118][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14701_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01346_),
    .Q(\mem[118][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14702_ (.CLK(clknet_leaf_90_i_clk),
    .D(_01347_),
    .Q(\mem[118][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14703_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01348_),
    .Q(\mem[118][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14704_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01349_),
    .Q(\mem[118][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14705_ (.CLK(clknet_leaf_101_i_clk),
    .D(_01350_),
    .Q(\mem[118][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14706_ (.CLK(clknet_leaf_101_i_clk),
    .D(_01351_),
    .Q(\mem[118][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14707_ (.CLK(clknet_leaf_130_i_clk),
    .D(_01352_),
    .Q(\mem[118][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14708_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01353_),
    .Q(\mem[118][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14709_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01354_),
    .Q(\mem[118][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14710_ (.CLK(clknet_leaf_145_i_clk),
    .D(_01355_),
    .Q(\mem[118][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14711_ (.CLK(clknet_leaf_134_i_clk),
    .D(_01356_),
    .Q(\mem[118][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14712_ (.CLK(clknet_leaf_146_i_clk),
    .D(_01357_),
    .Q(\mem[118][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14713_ (.CLK(clknet_leaf_124_i_clk),
    .D(_01358_),
    .Q(\mem[118][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14714_ (.CLK(clknet_leaf_148_i_clk),
    .D(_01359_),
    .Q(\mem[118][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14715_ (.CLK(clknet_leaf_146_i_clk),
    .D(_01360_),
    .Q(\mem[118][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14716_ (.CLK(clknet_leaf_115_i_clk),
    .D(_01361_),
    .Q(\mem[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14717_ (.CLK(clknet_leaf_116_i_clk),
    .D(_01362_),
    .Q(\mem[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14718_ (.CLK(clknet_leaf_117_i_clk),
    .D(_01363_),
    .Q(\mem[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14719_ (.CLK(clknet_leaf_126_i_clk),
    .D(_01364_),
    .Q(\mem[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14720_ (.CLK(clknet_leaf_116_i_clk),
    .D(_01365_),
    .Q(\mem[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14721_ (.CLK(clknet_leaf_114_i_clk),
    .D(_01366_),
    .Q(\mem[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14722_ (.CLK(clknet_leaf_126_i_clk),
    .D(_01367_),
    .Q(\mem[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14723_ (.CLK(clknet_leaf_117_i_clk),
    .D(_01368_),
    .Q(\mem[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14724_ (.CLK(clknet_leaf_120_i_clk),
    .D(_01369_),
    .Q(\mem[11][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14725_ (.CLK(clknet_leaf_122_i_clk),
    .D(_01370_),
    .Q(\mem[11][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14726_ (.CLK(clknet_leaf_140_i_clk),
    .D(_01371_),
    .Q(\mem[11][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14727_ (.CLK(clknet_leaf_136_i_clk),
    .D(_01372_),
    .Q(\mem[11][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14728_ (.CLK(clknet_leaf_141_i_clk),
    .D(_01373_),
    .Q(\mem[11][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14729_ (.CLK(clknet_leaf_120_i_clk),
    .D(_01374_),
    .Q(\mem[11][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14730_ (.CLK(clknet_leaf_141_i_clk),
    .D(_01375_),
    .Q(\mem[11][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14731_ (.CLK(clknet_leaf_142_i_clk),
    .D(_01376_),
    .Q(\mem[11][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14732_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01377_),
    .Q(\mem[120][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14733_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01378_),
    .Q(\mem[120][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14734_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01379_),
    .Q(\mem[120][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14735_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01380_),
    .Q(\mem[120][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14736_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01381_),
    .Q(\mem[120][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14737_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01382_),
    .Q(\mem[120][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14738_ (.CLK(clknet_leaf_96_i_clk),
    .D(_01383_),
    .Q(\mem[120][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14739_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01384_),
    .Q(\mem[120][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14740_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01385_),
    .Q(\mem[120][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14741_ (.CLK(clknet_leaf_134_i_clk),
    .D(_01386_),
    .Q(\mem[120][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14742_ (.CLK(clknet_leaf_148_i_clk),
    .D(_01387_),
    .Q(\mem[120][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14743_ (.CLK(clknet_leaf_135_i_clk),
    .D(_01388_),
    .Q(\mem[120][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14744_ (.CLK(clknet_leaf_149_i_clk),
    .D(_01389_),
    .Q(\mem[120][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14745_ (.CLK(clknet_leaf_137_i_clk),
    .D(_01390_),
    .Q(\mem[120][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14746_ (.CLK(clknet_leaf_149_i_clk),
    .D(_01391_),
    .Q(\mem[120][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14747_ (.CLK(clknet_leaf_149_i_clk),
    .D(_01392_),
    .Q(\mem[120][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14748_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01393_),
    .Q(\mem[121][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14749_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01394_),
    .Q(\mem[121][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14750_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01395_),
    .Q(\mem[121][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14751_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01396_),
    .Q(\mem[121][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14752_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01397_),
    .Q(\mem[121][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14753_ (.CLK(clknet_leaf_101_i_clk),
    .D(_01398_),
    .Q(\mem[121][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14754_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01399_),
    .Q(\mem[121][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14755_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01400_),
    .Q(\mem[121][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14756_ (.CLK(clknet_leaf_134_i_clk),
    .D(_01401_),
    .Q(\mem[121][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14757_ (.CLK(clknet_leaf_134_i_clk),
    .D(_01402_),
    .Q(\mem[121][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14758_ (.CLK(clknet_leaf_148_i_clk),
    .D(_01403_),
    .Q(\mem[121][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14759_ (.CLK(clknet_leaf_134_i_clk),
    .D(_01404_),
    .Q(\mem[121][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14760_ (.CLK(clknet_leaf_149_i_clk),
    .D(_01405_),
    .Q(\mem[121][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14761_ (.CLK(clknet_leaf_137_i_clk),
    .D(_01406_),
    .Q(\mem[121][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14762_ (.CLK(clknet_leaf_149_i_clk),
    .D(_01407_),
    .Q(\mem[121][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14763_ (.CLK(clknet_leaf_149_i_clk),
    .D(_01408_),
    .Q(\mem[121][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14764_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01409_),
    .Q(\mem[122][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14765_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01410_),
    .Q(\mem[122][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14766_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01411_),
    .Q(\mem[122][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14767_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01412_),
    .Q(\mem[122][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14768_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01413_),
    .Q(\mem[122][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14769_ (.CLK(clknet_leaf_101_i_clk),
    .D(_01414_),
    .Q(\mem[122][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14770_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01415_),
    .Q(\mem[122][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14771_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01416_),
    .Q(\mem[122][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14772_ (.CLK(clknet_leaf_132_i_clk),
    .D(_01417_),
    .Q(\mem[122][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14773_ (.CLK(clknet_leaf_134_i_clk),
    .D(_01418_),
    .Q(\mem[122][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14774_ (.CLK(clknet_leaf_148_i_clk),
    .D(_01419_),
    .Q(\mem[122][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14775_ (.CLK(clknet_leaf_134_i_clk),
    .D(_01420_),
    .Q(\mem[122][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14776_ (.CLK(clknet_leaf_149_i_clk),
    .D(_01421_),
    .Q(\mem[122][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14777_ (.CLK(clknet_leaf_133_i_clk),
    .D(_01422_),
    .Q(\mem[122][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14778_ (.CLK(clknet_leaf_148_i_clk),
    .D(_01423_),
    .Q(\mem[122][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14779_ (.CLK(clknet_leaf_150_i_clk),
    .D(_01424_),
    .Q(\mem[122][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14780_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01425_),
    .Q(\mem[123][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14781_ (.CLK(clknet_leaf_88_i_clk),
    .D(_01426_),
    .Q(\mem[123][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14782_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01427_),
    .Q(\mem[123][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14783_ (.CLK(clknet_leaf_92_i_clk),
    .D(_01428_),
    .Q(\mem[123][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14784_ (.CLK(clknet_leaf_91_i_clk),
    .D(_01429_),
    .Q(\mem[123][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14785_ (.CLK(clknet_leaf_93_i_clk),
    .D(_01430_),
    .Q(\mem[123][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14786_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01431_),
    .Q(\mem[123][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14787_ (.CLK(clknet_leaf_94_i_clk),
    .D(_01432_),
    .Q(\mem[123][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14788_ (.CLK(clknet_leaf_132_i_clk),
    .D(_01433_),
    .Q(\mem[123][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14789_ (.CLK(clknet_leaf_134_i_clk),
    .D(_01434_),
    .Q(\mem[123][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14790_ (.CLK(clknet_leaf_148_i_clk),
    .D(_01435_),
    .Q(\mem[123][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14791_ (.CLK(clknet_leaf_134_i_clk),
    .D(_01436_),
    .Q(\mem[123][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14792_ (.CLK(clknet_leaf_149_i_clk),
    .D(_01437_),
    .Q(\mem[123][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14793_ (.CLK(clknet_leaf_137_i_clk),
    .D(_01438_),
    .Q(\mem[123][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14794_ (.CLK(clknet_leaf_148_i_clk),
    .D(_01439_),
    .Q(\mem[123][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14795_ (.CLK(clknet_leaf_150_i_clk),
    .D(_01440_),
    .Q(\mem[123][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14796_ (.CLK(clknet_leaf_99_i_clk),
    .D(_01441_),
    .Q(\mem[124][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14797_ (.CLK(clknet_leaf_108_i_clk),
    .D(_01442_),
    .Q(\mem[124][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14798_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01443_),
    .Q(\mem[124][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14799_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01444_),
    .Q(\mem[124][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14800_ (.CLK(clknet_leaf_127_i_clk),
    .D(_01445_),
    .Q(\mem[124][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14801_ (.CLK(clknet_leaf_99_i_clk),
    .D(_01446_),
    .Q(\mem[124][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14802_ (.CLK(clknet_leaf_126_i_clk),
    .D(_01447_),
    .Q(\mem[124][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14803_ (.CLK(clknet_leaf_127_i_clk),
    .D(_01448_),
    .Q(\mem[124][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14804_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01449_),
    .Q(\mem[124][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14805_ (.CLK(clknet_leaf_123_i_clk),
    .D(_01450_),
    .Q(\mem[124][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14806_ (.CLK(clknet_leaf_143_i_clk),
    .D(_01451_),
    .Q(\mem[124][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14807_ (.CLK(clknet_leaf_138_i_clk),
    .D(_01452_),
    .Q(\mem[124][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14808_ (.CLK(clknet_leaf_143_i_clk),
    .D(_01453_),
    .Q(\mem[124][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14809_ (.CLK(clknet_leaf_124_i_clk),
    .D(_01454_),
    .Q(\mem[124][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14810_ (.CLK(clknet_leaf_143_i_clk),
    .D(_01455_),
    .Q(\mem[124][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14811_ (.CLK(clknet_leaf_135_i_clk),
    .D(_01456_),
    .Q(\mem[124][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14812_ (.CLK(clknet_leaf_99_i_clk),
    .D(_01457_),
    .Q(\mem[125][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14813_ (.CLK(clknet_leaf_108_i_clk),
    .D(_01458_),
    .Q(\mem[125][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14814_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01459_),
    .Q(\mem[125][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14815_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01460_),
    .Q(\mem[125][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14816_ (.CLK(clknet_leaf_127_i_clk),
    .D(_01461_),
    .Q(\mem[125][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14817_ (.CLK(clknet_leaf_126_i_clk),
    .D(_01462_),
    .Q(\mem[125][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14818_ (.CLK(clknet_leaf_126_i_clk),
    .D(_01463_),
    .Q(\mem[125][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14819_ (.CLK(clknet_leaf_127_i_clk),
    .D(_01464_),
    .Q(\mem[125][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14820_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01465_),
    .Q(\mem[125][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14821_ (.CLK(clknet_leaf_124_i_clk),
    .D(_01466_),
    .Q(\mem[125][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14822_ (.CLK(clknet_leaf_144_i_clk),
    .D(_01467_),
    .Q(\mem[125][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14823_ (.CLK(clknet_leaf_138_i_clk),
    .D(_01468_),
    .Q(\mem[125][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14824_ (.CLK(clknet_leaf_143_i_clk),
    .D(_01469_),
    .Q(\mem[125][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14825_ (.CLK(clknet_leaf_125_i_clk),
    .D(_01470_),
    .Q(\mem[125][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14826_ (.CLK(clknet_leaf_135_i_clk),
    .D(_01471_),
    .Q(\mem[125][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14827_ (.CLK(clknet_leaf_135_i_clk),
    .D(_01472_),
    .Q(\mem[125][15] ));
 sky130_fd_sc_hd__dfxtp_1 _14828_ (.CLK(clknet_leaf_100_i_clk),
    .D(_01473_),
    .Q(\mem[126][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14829_ (.CLK(clknet_leaf_100_i_clk),
    .D(_01474_),
    .Q(\mem[126][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14830_ (.CLK(clknet_leaf_100_i_clk),
    .D(_01475_),
    .Q(\mem[126][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14831_ (.CLK(clknet_leaf_97_i_clk),
    .D(_01476_),
    .Q(\mem[126][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14832_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01477_),
    .Q(\mem[126][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14833_ (.CLK(clknet_leaf_99_i_clk),
    .D(_01478_),
    .Q(\mem[126][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14834_ (.CLK(clknet_leaf_127_i_clk),
    .D(_01479_),
    .Q(\mem[126][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14835_ (.CLK(clknet_leaf_98_i_clk),
    .D(_01480_),
    .Q(\mem[126][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14836_ (.CLK(clknet_leaf_128_i_clk),
    .D(_01481_),
    .Q(\mem[126][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14837_ (.CLK(clknet_leaf_129_i_clk),
    .D(_01482_),
    .Q(\mem[126][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14838_ (.CLK(clknet_leaf_144_i_clk),
    .D(_01483_),
    .Q(\mem[126][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14839_ (.CLK(clknet_leaf_138_i_clk),
    .D(_01484_),
    .Q(\mem[126][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14840_ (.CLK(clknet_leaf_143_i_clk),
    .D(_01485_),
    .Q(\mem[126][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14841_ (.CLK(clknet_leaf_125_i_clk),
    .D(_01486_),
    .Q(\mem[126][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14842_ (.CLK(clknet_leaf_135_i_clk),
    .D(_01487_),
    .Q(\mem[126][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14843_ (.CLK(clknet_leaf_136_i_clk),
    .D(_01488_),
    .Q(\mem[126][15] ));
 sky130_fd_sc_hd__dfxtp_2 _14844_ (.CLK(clknet_leaf_251_i_clk),
    .D(_00000_),
    .Q(net25));
 sky130_fd_sc_hd__dfxtp_4 _14845_ (.CLK(clknet_leaf_112_i_clk),
    .D(_00007_),
    .Q(net32));
 sky130_fd_sc_hd__dfxtp_2 _14846_ (.CLK(clknet_leaf_251_i_clk),
    .D(_00008_),
    .Q(net33));
 sky130_fd_sc_hd__dfxtp_2 _14847_ (.CLK(clknet_leaf_252_i_clk),
    .D(_00009_),
    .Q(net34));
 sky130_fd_sc_hd__dfxtp_2 _14848_ (.CLK(clknet_leaf_251_i_clk),
    .D(_00010_),
    .Q(net35));
 sky130_fd_sc_hd__dfxtp_2 _14849_ (.CLK(clknet_leaf_112_i_clk),
    .D(_00011_),
    .Q(net36));
 sky130_fd_sc_hd__dfxtp_2 _14850_ (.CLK(clknet_leaf_182_i_clk),
    .D(_00012_),
    .Q(net37));
 sky130_fd_sc_hd__dfxtp_2 _14851_ (.CLK(clknet_leaf_181_i_clk),
    .D(_00013_),
    .Q(net38));
 sky130_fd_sc_hd__dfxtp_2 _14852_ (.CLK(clknet_leaf_180_i_clk),
    .D(_00014_),
    .Q(net39));
 sky130_fd_sc_hd__dfxtp_2 _14853_ (.CLK(clknet_leaf_180_i_clk),
    .D(_00015_),
    .Q(net40));
 sky130_fd_sc_hd__dfxtp_2 _14854_ (.CLK(clknet_leaf_169_i_clk),
    .D(_00001_),
    .Q(net26));
 sky130_fd_sc_hd__dfxtp_2 _14855_ (.CLK(clknet_leaf_180_i_clk),
    .D(_00002_),
    .Q(net27));
 sky130_fd_sc_hd__dfxtp_2 _14856_ (.CLK(clknet_leaf_169_i_clk),
    .D(_00003_),
    .Q(net28));
 sky130_fd_sc_hd__dfxtp_2 _14857_ (.CLK(clknet_leaf_112_i_clk),
    .D(_00004_),
    .Q(net29));
 sky130_fd_sc_hd__dfxtp_2 _14858_ (.CLK(clknet_leaf_169_i_clk),
    .D(_00005_),
    .Q(net30));
 sky130_fd_sc_hd__dfxtp_2 _14859_ (.CLK(clknet_leaf_177_i_clk),
    .D(_00006_),
    .Q(net31));
 sky130_fd_sc_hd__dfxtp_1 _14860_ (.CLK(clknet_leaf_115_i_clk),
    .D(_01489_),
    .Q(\mem[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 _14861_ (.CLK(clknet_leaf_116_i_clk),
    .D(_01490_),
    .Q(\mem[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 _14862_ (.CLK(clknet_leaf_125_i_clk),
    .D(_01491_),
    .Q(\mem[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 _14863_ (.CLK(clknet_leaf_117_i_clk),
    .D(_01492_),
    .Q(\mem[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 _14864_ (.CLK(clknet_leaf_117_i_clk),
    .D(_01493_),
    .Q(\mem[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 _14865_ (.CLK(clknet_leaf_115_i_clk),
    .D(_01494_),
    .Q(\mem[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 _14866_ (.CLK(clknet_leaf_125_i_clk),
    .D(_01495_),
    .Q(\mem[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 _14867_ (.CLK(clknet_leaf_118_i_clk),
    .D(_01496_),
    .Q(\mem[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 _14868_ (.CLK(clknet_leaf_120_i_clk),
    .D(_01497_),
    .Q(\mem[9][8] ));
 sky130_fd_sc_hd__dfxtp_1 _14869_ (.CLK(clknet_leaf_122_i_clk),
    .D(_01498_),
    .Q(\mem[9][9] ));
 sky130_fd_sc_hd__dfxtp_1 _14870_ (.CLK(clknet_leaf_141_i_clk),
    .D(_01499_),
    .Q(\mem[9][10] ));
 sky130_fd_sc_hd__dfxtp_1 _14871_ (.CLK(clknet_leaf_143_i_clk),
    .D(_01500_),
    .Q(\mem[9][11] ));
 sky130_fd_sc_hd__dfxtp_1 _14872_ (.CLK(clknet_leaf_141_i_clk),
    .D(_01501_),
    .Q(\mem[9][12] ));
 sky130_fd_sc_hd__dfxtp_1 _14873_ (.CLK(clknet_leaf_119_i_clk),
    .D(_01502_),
    .Q(\mem[9][13] ));
 sky130_fd_sc_hd__dfxtp_1 _14874_ (.CLK(clknet_leaf_141_i_clk),
    .D(_01503_),
    .Q(\mem[9][14] ));
 sky130_fd_sc_hd__dfxtp_1 _14875_ (.CLK(clknet_leaf_142_i_clk),
    .D(_01504_),
    .Q(\mem[9][15] ));
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(i_addr[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(i_addr[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input3 (.A(i_addr[2]),
    .X(net3));
 sky130_fd_sc_hd__buf_8 input4 (.A(i_addr[3]),
    .X(net4));
 sky130_fd_sc_hd__buf_4 input5 (.A(i_addr[4]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(i_addr[5]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(i_addr[6]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_4 input8 (.A(i_data[0]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input9 (.A(i_data[10]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(i_data[11]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(i_data[12]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(i_data[13]),
    .X(net12));
 sky130_fd_sc_hd__dlymetal6s2s_1 input13 (.A(i_data[14]),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 input14 (.A(i_data[15]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(i_data[1]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 input16 (.A(i_data[2]),
    .X(net16));
 sky130_fd_sc_hd__buf_2 input17 (.A(i_data[3]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 input18 (.A(i_data[4]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 input19 (.A(i_data[5]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 input20 (.A(i_data[6]),
    .X(net20));
 sky130_fd_sc_hd__buf_2 input21 (.A(i_data[7]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(i_data[8]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 input23 (.A(i_data[9]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(i_we),
    .X(net24));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(o_data[0]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(o_data[10]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(o_data[11]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(o_data[12]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(o_data[13]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(o_data[14]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(o_data[15]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(o_data[1]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(o_data[2]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(o_data[3]));
 sky130_fd_sc_hd__buf_2 output35 (.A(net35),
    .X(o_data[4]));
 sky130_fd_sc_hd__buf_2 output36 (.A(net36),
    .X(o_data[5]));
 sky130_fd_sc_hd__buf_2 output37 (.A(net37),
    .X(o_data[6]));
 sky130_fd_sc_hd__buf_2 output38 (.A(net38),
    .X(o_data[7]));
 sky130_fd_sc_hd__buf_2 output39 (.A(net39),
    .X(o_data[8]));
 sky130_fd_sc_hd__buf_2 output40 (.A(net40),
    .X(o_data[9]));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_i_clk (.A(clknet_5_0_0_i_clk),
    .X(clknet_leaf_0_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_i_clk (.A(clknet_5_0_0_i_clk),
    .X(clknet_leaf_1_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_i_clk (.A(clknet_5_0_0_i_clk),
    .X(clknet_leaf_2_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_i_clk (.A(clknet_5_0_0_i_clk),
    .X(clknet_leaf_3_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_i_clk (.A(clknet_5_0_0_i_clk),
    .X(clknet_leaf_4_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_i_clk (.A(clknet_5_0_0_i_clk),
    .X(clknet_leaf_5_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_i_clk (.A(clknet_5_1_0_i_clk),
    .X(clknet_leaf_6_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_i_clk (.A(clknet_5_1_0_i_clk),
    .X(clknet_leaf_7_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_i_clk (.A(clknet_5_1_0_i_clk),
    .X(clknet_leaf_8_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_i_clk (.A(clknet_5_3_0_i_clk),
    .X(clknet_leaf_9_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_i_clk (.A(clknet_5_3_0_i_clk),
    .X(clknet_leaf_10_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_i_clk (.A(clknet_5_2_0_i_clk),
    .X(clknet_leaf_11_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_i_clk (.A(clknet_5_2_0_i_clk),
    .X(clknet_leaf_12_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_i_clk (.A(clknet_5_2_0_i_clk),
    .X(clknet_leaf_13_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_i_clk (.A(clknet_5_2_0_i_clk),
    .X(clknet_leaf_14_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_i_clk (.A(clknet_5_2_0_i_clk),
    .X(clknet_leaf_15_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_i_clk (.A(clknet_5_2_0_i_clk),
    .X(clknet_leaf_16_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_i_clk (.A(clknet_5_2_0_i_clk),
    .X(clknet_leaf_17_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_i_clk (.A(clknet_5_2_0_i_clk),
    .X(clknet_leaf_18_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_i_clk (.A(clknet_5_2_0_i_clk),
    .X(clknet_leaf_19_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_i_clk (.A(clknet_5_2_0_i_clk),
    .X(clknet_leaf_20_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_i_clk (.A(clknet_5_3_0_i_clk),
    .X(clknet_leaf_21_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_i_clk (.A(clknet_5_3_0_i_clk),
    .X(clknet_leaf_22_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_i_clk (.A(clknet_5_3_0_i_clk),
    .X(clknet_leaf_23_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_i_clk (.A(clknet_5_3_0_i_clk),
    .X(clknet_leaf_24_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_i_clk (.A(clknet_5_3_0_i_clk),
    .X(clknet_leaf_25_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_i_clk (.A(clknet_5_3_0_i_clk),
    .X(clknet_leaf_26_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_i_clk (.A(clknet_5_3_0_i_clk),
    .X(clknet_leaf_27_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_i_clk (.A(clknet_5_3_0_i_clk),
    .X(clknet_leaf_28_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_i_clk (.A(clknet_5_6_0_i_clk),
    .X(clknet_leaf_29_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_i_clk (.A(clknet_5_6_0_i_clk),
    .X(clknet_leaf_30_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_i_clk (.A(clknet_5_6_0_i_clk),
    .X(clknet_leaf_31_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_i_clk (.A(clknet_5_6_0_i_clk),
    .X(clknet_leaf_32_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_i_clk (.A(clknet_5_6_0_i_clk),
    .X(clknet_leaf_33_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_i_clk (.A(clknet_5_6_0_i_clk),
    .X(clknet_leaf_34_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_i_clk (.A(clknet_5_6_0_i_clk),
    .X(clknet_leaf_35_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_i_clk (.A(clknet_5_7_0_i_clk),
    .X(clknet_leaf_36_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_i_clk (.A(clknet_5_7_0_i_clk),
    .X(clknet_leaf_37_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_i_clk (.A(clknet_5_7_0_i_clk),
    .X(clknet_leaf_38_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_i_clk (.A(clknet_5_13_0_i_clk),
    .X(clknet_leaf_39_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_i_clk (.A(clknet_5_13_0_i_clk),
    .X(clknet_leaf_40_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_i_clk (.A(clknet_5_12_0_i_clk),
    .X(clknet_leaf_41_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_i_clk (.A(clknet_5_12_0_i_clk),
    .X(clknet_leaf_42_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_i_clk (.A(clknet_5_12_0_i_clk),
    .X(clknet_leaf_43_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_i_clk (.A(clknet_5_12_0_i_clk),
    .X(clknet_leaf_44_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_i_clk (.A(clknet_5_12_0_i_clk),
    .X(clknet_leaf_45_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_i_clk (.A(clknet_5_12_0_i_clk),
    .X(clknet_leaf_46_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_i_clk (.A(clknet_5_12_0_i_clk),
    .X(clknet_leaf_47_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_i_clk (.A(clknet_5_9_0_i_clk),
    .X(clknet_leaf_48_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_i_clk (.A(clknet_5_9_0_i_clk),
    .X(clknet_leaf_49_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_50_i_clk (.A(clknet_5_9_0_i_clk),
    .X(clknet_leaf_50_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_i_clk (.A(clknet_5_9_0_i_clk),
    .X(clknet_leaf_51_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_52_i_clk (.A(clknet_5_9_0_i_clk),
    .X(clknet_leaf_52_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_i_clk (.A(clknet_5_9_0_i_clk),
    .X(clknet_leaf_53_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_i_clk (.A(clknet_5_9_0_i_clk),
    .X(clknet_leaf_54_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_i_clk (.A(clknet_5_8_0_i_clk),
    .X(clknet_leaf_55_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_i_clk (.A(clknet_5_8_0_i_clk),
    .X(clknet_leaf_56_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_i_clk (.A(clknet_5_8_0_i_clk),
    .X(clknet_leaf_57_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_i_clk (.A(clknet_5_8_0_i_clk),
    .X(clknet_leaf_58_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_i_clk (.A(clknet_5_8_0_i_clk),
    .X(clknet_leaf_59_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_i_clk (.A(clknet_5_8_0_i_clk),
    .X(clknet_leaf_60_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_61_i_clk (.A(clknet_5_8_0_i_clk),
    .X(clknet_leaf_61_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_i_clk (.A(clknet_5_8_0_i_clk),
    .X(clknet_leaf_62_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_i_clk (.A(clknet_5_8_0_i_clk),
    .X(clknet_leaf_63_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_64_i_clk (.A(clknet_5_8_0_i_clk),
    .X(clknet_leaf_64_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_i_clk (.A(clknet_5_8_0_i_clk),
    .X(clknet_leaf_65_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_i_clk (.A(clknet_5_9_0_i_clk),
    .X(clknet_leaf_66_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_i_clk (.A(clknet_5_9_0_i_clk),
    .X(clknet_leaf_67_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_68_i_clk (.A(clknet_5_9_0_i_clk),
    .X(clknet_leaf_68_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_i_clk (.A(clknet_5_9_0_i_clk),
    .X(clknet_leaf_69_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_i_clk (.A(clknet_5_11_0_i_clk),
    .X(clknet_leaf_70_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_71_i_clk (.A(clknet_5_11_0_i_clk),
    .X(clknet_leaf_71_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_i_clk (.A(clknet_5_10_0_i_clk),
    .X(clknet_leaf_72_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_i_clk (.A(clknet_5_10_0_i_clk),
    .X(clknet_leaf_73_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_i_clk (.A(clknet_5_10_0_i_clk),
    .X(clknet_leaf_74_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_i_clk (.A(clknet_5_10_0_i_clk),
    .X(clknet_leaf_75_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_i_clk (.A(clknet_5_10_0_i_clk),
    .X(clknet_leaf_76_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_i_clk (.A(clknet_5_10_0_i_clk),
    .X(clknet_leaf_77_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_i_clk (.A(clknet_5_10_0_i_clk),
    .X(clknet_leaf_78_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_i_clk (.A(clknet_5_11_0_i_clk),
    .X(clknet_leaf_79_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_i_clk (.A(clknet_5_11_0_i_clk),
    .X(clknet_leaf_80_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_i_clk (.A(clknet_5_11_0_i_clk),
    .X(clknet_leaf_81_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_i_clk (.A(clknet_5_11_0_i_clk),
    .X(clknet_leaf_82_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_i_clk (.A(clknet_5_11_0_i_clk),
    .X(clknet_leaf_83_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_i_clk (.A(clknet_5_11_0_i_clk),
    .X(clknet_leaf_84_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_i_clk (.A(clknet_5_11_0_i_clk),
    .X(clknet_leaf_85_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_i_clk (.A(clknet_5_14_0_i_clk),
    .X(clknet_leaf_86_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_i_clk (.A(clknet_5_14_0_i_clk),
    .X(clknet_leaf_87_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_i_clk (.A(clknet_5_14_0_i_clk),
    .X(clknet_leaf_88_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_i_clk (.A(clknet_5_14_0_i_clk),
    .X(clknet_leaf_89_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_i_clk (.A(clknet_5_14_0_i_clk),
    .X(clknet_leaf_90_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_i_clk (.A(clknet_5_14_0_i_clk),
    .X(clknet_leaf_91_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_i_clk (.A(clknet_5_14_0_i_clk),
    .X(clknet_leaf_92_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_i_clk (.A(clknet_5_15_0_i_clk),
    .X(clknet_leaf_93_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_i_clk (.A(clknet_5_15_0_i_clk),
    .X(clknet_leaf_94_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_i_clk (.A(clknet_5_15_0_i_clk),
    .X(clknet_leaf_95_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_i_clk (.A(clknet_5_15_0_i_clk),
    .X(clknet_leaf_96_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_i_clk (.A(clknet_5_15_0_i_clk),
    .X(clknet_leaf_97_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_98_i_clk (.A(clknet_5_15_0_i_clk),
    .X(clknet_leaf_98_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_i_clk (.A(clknet_5_15_0_i_clk),
    .X(clknet_leaf_99_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_i_clk (.A(clknet_5_15_0_i_clk),
    .X(clknet_leaf_100_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_101_i_clk (.A(clknet_5_14_0_i_clk),
    .X(clknet_leaf_101_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_i_clk (.A(clknet_5_14_0_i_clk),
    .X(clknet_leaf_102_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_i_clk (.A(clknet_5_14_0_i_clk),
    .X(clknet_leaf_103_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_i_clk (.A(clknet_5_12_0_i_clk),
    .X(clknet_leaf_104_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_i_clk (.A(clknet_5_12_0_i_clk),
    .X(clknet_leaf_105_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_i_clk (.A(clknet_5_13_0_i_clk),
    .X(clknet_leaf_106_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_i_clk (.A(clknet_5_13_0_i_clk),
    .X(clknet_leaf_107_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_108_i_clk (.A(clknet_5_13_0_i_clk),
    .X(clknet_leaf_108_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_i_clk (.A(clknet_5_13_0_i_clk),
    .X(clknet_leaf_109_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_i_clk (.A(clknet_5_13_0_i_clk),
    .X(clknet_leaf_110_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_i_clk (.A(clknet_5_13_0_i_clk),
    .X(clknet_leaf_111_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_i_clk (.A(clknet_5_13_0_i_clk),
    .X(clknet_leaf_112_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_i_clk (.A(clknet_5_24_0_i_clk),
    .X(clknet_leaf_113_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_i_clk (.A(clknet_5_24_0_i_clk),
    .X(clknet_leaf_114_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_i_clk (.A(clknet_5_24_0_i_clk),
    .X(clknet_leaf_115_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_i_clk (.A(clknet_5_24_0_i_clk),
    .X(clknet_leaf_116_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_i_clk (.A(clknet_5_24_0_i_clk),
    .X(clknet_leaf_117_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_i_clk (.A(clknet_5_24_0_i_clk),
    .X(clknet_leaf_118_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_119_i_clk (.A(clknet_5_25_0_i_clk),
    .X(clknet_leaf_119_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_i_clk (.A(clknet_5_25_0_i_clk),
    .X(clknet_leaf_120_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_121_i_clk (.A(clknet_5_27_0_i_clk),
    .X(clknet_leaf_121_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_i_clk (.A(clknet_5_27_0_i_clk),
    .X(clknet_leaf_122_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_i_clk (.A(clknet_5_27_0_i_clk),
    .X(clknet_leaf_123_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_i_clk (.A(clknet_5_26_0_i_clk),
    .X(clknet_leaf_124_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_125_i_clk (.A(clknet_5_26_0_i_clk),
    .X(clknet_leaf_125_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_i_clk (.A(clknet_5_26_0_i_clk),
    .X(clknet_leaf_126_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_i_clk (.A(clknet_5_26_0_i_clk),
    .X(clknet_leaf_127_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_i_clk (.A(clknet_5_26_0_i_clk),
    .X(clknet_leaf_128_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_129_i_clk (.A(clknet_5_26_0_i_clk),
    .X(clknet_leaf_129_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_130_i_clk (.A(clknet_5_26_0_i_clk),
    .X(clknet_leaf_130_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_131_i_clk (.A(clknet_5_26_0_i_clk),
    .X(clknet_leaf_131_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_132_i_clk (.A(clknet_5_26_0_i_clk),
    .X(clknet_leaf_132_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_133_i_clk (.A(clknet_5_27_0_i_clk),
    .X(clknet_leaf_133_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_134_i_clk (.A(clknet_5_27_0_i_clk),
    .X(clknet_leaf_134_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_135_i_clk (.A(clknet_5_27_0_i_clk),
    .X(clknet_leaf_135_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_136_i_clk (.A(clknet_5_27_0_i_clk),
    .X(clknet_leaf_136_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_137_i_clk (.A(clknet_5_27_0_i_clk),
    .X(clknet_leaf_137_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_138_i_clk (.A(clknet_5_27_0_i_clk),
    .X(clknet_leaf_138_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_139_i_clk (.A(clknet_5_27_0_i_clk),
    .X(clknet_leaf_139_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_140_i_clk (.A(clknet_5_30_0_i_clk),
    .X(clknet_leaf_140_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_141_i_clk (.A(clknet_5_30_0_i_clk),
    .X(clknet_leaf_141_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_142_i_clk (.A(clknet_5_30_0_i_clk),
    .X(clknet_leaf_142_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_143_i_clk (.A(clknet_5_30_0_i_clk),
    .X(clknet_leaf_143_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_144_i_clk (.A(clknet_5_30_0_i_clk),
    .X(clknet_leaf_144_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_145_i_clk (.A(clknet_5_30_0_i_clk),
    .X(clknet_leaf_145_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_146_i_clk (.A(clknet_5_30_0_i_clk),
    .X(clknet_leaf_146_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_147_i_clk (.A(clknet_5_31_0_i_clk),
    .X(clknet_leaf_147_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_148_i_clk (.A(clknet_5_31_0_i_clk),
    .X(clknet_leaf_148_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_149_i_clk (.A(clknet_5_31_0_i_clk),
    .X(clknet_leaf_149_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_150_i_clk (.A(clknet_5_31_0_i_clk),
    .X(clknet_leaf_150_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_151_i_clk (.A(clknet_5_31_0_i_clk),
    .X(clknet_leaf_151_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_152_i_clk (.A(clknet_5_31_0_i_clk),
    .X(clknet_leaf_152_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_153_i_clk (.A(clknet_5_31_0_i_clk),
    .X(clknet_leaf_153_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_154_i_clk (.A(clknet_5_31_0_i_clk),
    .X(clknet_leaf_154_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_155_i_clk (.A(clknet_5_31_0_i_clk),
    .X(clknet_leaf_155_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_156_i_clk (.A(clknet_5_30_0_i_clk),
    .X(clknet_leaf_156_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_157_i_clk (.A(clknet_5_30_0_i_clk),
    .X(clknet_leaf_157_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_158_i_clk (.A(clknet_5_28_0_i_clk),
    .X(clknet_leaf_158_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_159_i_clk (.A(clknet_5_28_0_i_clk),
    .X(clknet_leaf_159_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_160_i_clk (.A(clknet_5_29_0_i_clk),
    .X(clknet_leaf_160_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_161_i_clk (.A(clknet_5_29_0_i_clk),
    .X(clknet_leaf_161_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_162_i_clk (.A(clknet_5_29_0_i_clk),
    .X(clknet_leaf_162_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_163_i_clk (.A(clknet_5_29_0_i_clk),
    .X(clknet_leaf_163_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_164_i_clk (.A(clknet_5_29_0_i_clk),
    .X(clknet_leaf_164_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_165_i_clk (.A(clknet_5_29_0_i_clk),
    .X(clknet_leaf_165_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_166_i_clk (.A(clknet_5_29_0_i_clk),
    .X(clknet_leaf_166_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_167_i_clk (.A(clknet_5_29_0_i_clk),
    .X(clknet_leaf_167_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_168_i_clk (.A(clknet_5_28_0_i_clk),
    .X(clknet_leaf_168_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_169_i_clk (.A(clknet_5_28_0_i_clk),
    .X(clknet_leaf_169_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_170_i_clk (.A(clknet_5_28_0_i_clk),
    .X(clknet_leaf_170_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_171_i_clk (.A(clknet_5_28_0_i_clk),
    .X(clknet_leaf_171_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_172_i_clk (.A(clknet_5_28_0_i_clk),
    .X(clknet_leaf_172_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_173_i_clk (.A(clknet_5_25_0_i_clk),
    .X(clknet_leaf_173_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_174_i_clk (.A(clknet_5_25_0_i_clk),
    .X(clknet_leaf_174_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_175_i_clk (.A(clknet_5_25_0_i_clk),
    .X(clknet_leaf_175_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_176_i_clk (.A(clknet_5_25_0_i_clk),
    .X(clknet_leaf_176_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_177_i_clk (.A(clknet_5_25_0_i_clk),
    .X(clknet_leaf_177_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_178_i_clk (.A(clknet_5_25_0_i_clk),
    .X(clknet_leaf_178_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_179_i_clk (.A(clknet_5_24_0_i_clk),
    .X(clknet_leaf_179_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_180_i_clk (.A(clknet_5_24_0_i_clk),
    .X(clknet_leaf_180_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_181_i_clk (.A(clknet_5_18_0_i_clk),
    .X(clknet_leaf_181_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_182_i_clk (.A(clknet_5_18_0_i_clk),
    .X(clknet_leaf_182_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_183_i_clk (.A(clknet_5_19_0_i_clk),
    .X(clknet_leaf_183_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_184_i_clk (.A(clknet_5_19_0_i_clk),
    .X(clknet_leaf_184_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_185_i_clk (.A(clknet_5_19_0_i_clk),
    .X(clknet_leaf_185_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_186_i_clk (.A(clknet_5_19_0_i_clk),
    .X(clknet_leaf_186_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_187_i_clk (.A(clknet_5_19_0_i_clk),
    .X(clknet_leaf_187_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_188_i_clk (.A(clknet_5_19_0_i_clk),
    .X(clknet_leaf_188_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_189_i_clk (.A(clknet_5_19_0_i_clk),
    .X(clknet_leaf_189_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_190_i_clk (.A(clknet_5_22_0_i_clk),
    .X(clknet_leaf_190_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_191_i_clk (.A(clknet_5_22_0_i_clk),
    .X(clknet_leaf_191_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_192_i_clk (.A(clknet_5_22_0_i_clk),
    .X(clknet_leaf_192_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_193_i_clk (.A(clknet_5_22_0_i_clk),
    .X(clknet_leaf_193_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_194_i_clk (.A(clknet_5_22_0_i_clk),
    .X(clknet_leaf_194_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_195_i_clk (.A(clknet_5_22_0_i_clk),
    .X(clknet_leaf_195_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_196_i_clk (.A(clknet_5_22_0_i_clk),
    .X(clknet_leaf_196_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_197_i_clk (.A(clknet_5_23_0_i_clk),
    .X(clknet_leaf_197_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_198_i_clk (.A(clknet_5_23_0_i_clk),
    .X(clknet_leaf_198_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_199_i_clk (.A(clknet_5_23_0_i_clk),
    .X(clknet_leaf_199_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_200_i_clk (.A(clknet_5_23_0_i_clk),
    .X(clknet_leaf_200_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_201_i_clk (.A(clknet_5_23_0_i_clk),
    .X(clknet_leaf_201_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_202_i_clk (.A(clknet_5_23_0_i_clk),
    .X(clknet_leaf_202_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_203_i_clk (.A(clknet_5_23_0_i_clk),
    .X(clknet_leaf_203_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_204_i_clk (.A(clknet_5_23_0_i_clk),
    .X(clknet_leaf_204_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_205_i_clk (.A(clknet_5_23_0_i_clk),
    .X(clknet_leaf_205_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_206_i_clk (.A(clknet_5_23_0_i_clk),
    .X(clknet_leaf_206_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_207_i_clk (.A(clknet_5_22_0_i_clk),
    .X(clknet_leaf_207_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_208_i_clk (.A(clknet_5_22_0_i_clk),
    .X(clknet_leaf_208_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_209_i_clk (.A(clknet_5_20_0_i_clk),
    .X(clknet_leaf_209_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_210_i_clk (.A(clknet_5_20_0_i_clk),
    .X(clknet_leaf_210_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_211_i_clk (.A(clknet_5_21_0_i_clk),
    .X(clknet_leaf_211_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_212_i_clk (.A(clknet_5_21_0_i_clk),
    .X(clknet_leaf_212_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_213_i_clk (.A(clknet_5_21_0_i_clk),
    .X(clknet_leaf_213_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_214_i_clk (.A(clknet_5_21_0_i_clk),
    .X(clknet_leaf_214_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_215_i_clk (.A(clknet_5_21_0_i_clk),
    .X(clknet_leaf_215_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_216_i_clk (.A(clknet_5_21_0_i_clk),
    .X(clknet_leaf_216_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_217_i_clk (.A(clknet_5_21_0_i_clk),
    .X(clknet_leaf_217_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_218_i_clk (.A(clknet_5_21_0_i_clk),
    .X(clknet_leaf_218_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_219_i_clk (.A(clknet_5_21_0_i_clk),
    .X(clknet_leaf_219_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_220_i_clk (.A(clknet_5_21_0_i_clk),
    .X(clknet_leaf_220_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_221_i_clk (.A(clknet_5_20_0_i_clk),
    .X(clknet_leaf_221_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_222_i_clk (.A(clknet_5_20_0_i_clk),
    .X(clknet_leaf_222_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_223_i_clk (.A(clknet_5_20_0_i_clk),
    .X(clknet_leaf_223_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_224_i_clk (.A(clknet_5_20_0_i_clk),
    .X(clknet_leaf_224_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_225_i_clk (.A(clknet_5_20_0_i_clk),
    .X(clknet_leaf_225_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_226_i_clk (.A(clknet_5_20_0_i_clk),
    .X(clknet_leaf_226_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_227_i_clk (.A(clknet_5_17_0_i_clk),
    .X(clknet_leaf_227_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_228_i_clk (.A(clknet_5_17_0_i_clk),
    .X(clknet_leaf_228_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_229_i_clk (.A(clknet_5_17_0_i_clk),
    .X(clknet_leaf_229_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_230_i_clk (.A(clknet_5_17_0_i_clk),
    .X(clknet_leaf_230_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_231_i_clk (.A(clknet_5_17_0_i_clk),
    .X(clknet_leaf_231_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_232_i_clk (.A(clknet_5_17_0_i_clk),
    .X(clknet_leaf_232_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_233_i_clk (.A(clknet_5_17_0_i_clk),
    .X(clknet_leaf_233_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_234_i_clk (.A(clknet_5_16_0_i_clk),
    .X(clknet_leaf_234_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_235_i_clk (.A(clknet_5_16_0_i_clk),
    .X(clknet_leaf_235_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_236_i_clk (.A(clknet_5_16_0_i_clk),
    .X(clknet_leaf_236_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_237_i_clk (.A(clknet_5_16_0_i_clk),
    .X(clknet_leaf_237_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_238_i_clk (.A(clknet_5_16_0_i_clk),
    .X(clknet_leaf_238_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_239_i_clk (.A(clknet_5_16_0_i_clk),
    .X(clknet_leaf_239_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_240_i_clk (.A(clknet_5_16_0_i_clk),
    .X(clknet_leaf_240_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_241_i_clk (.A(clknet_5_16_0_i_clk),
    .X(clknet_leaf_241_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_242_i_clk (.A(clknet_5_17_0_i_clk),
    .X(clknet_leaf_242_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_243_i_clk (.A(clknet_5_19_0_i_clk),
    .X(clknet_leaf_243_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_244_i_clk (.A(clknet_5_19_0_i_clk),
    .X(clknet_leaf_244_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_245_i_clk (.A(clknet_5_19_0_i_clk),
    .X(clknet_leaf_245_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_246_i_clk (.A(clknet_5_18_0_i_clk),
    .X(clknet_leaf_246_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_247_i_clk (.A(clknet_5_18_0_i_clk),
    .X(clknet_leaf_247_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_248_i_clk (.A(clknet_5_18_0_i_clk),
    .X(clknet_leaf_248_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_249_i_clk (.A(clknet_5_18_0_i_clk),
    .X(clknet_leaf_249_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_250_i_clk (.A(clknet_5_18_0_i_clk),
    .X(clknet_leaf_250_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_251_i_clk (.A(clknet_5_18_0_i_clk),
    .X(clknet_leaf_251_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_252_i_clk (.A(clknet_5_7_0_i_clk),
    .X(clknet_leaf_252_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_253_i_clk (.A(clknet_5_7_0_i_clk),
    .X(clknet_leaf_253_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_254_i_clk (.A(clknet_5_7_0_i_clk),
    .X(clknet_leaf_254_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_255_i_clk (.A(clknet_5_7_0_i_clk),
    .X(clknet_leaf_255_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_256_i_clk (.A(clknet_5_7_0_i_clk),
    .X(clknet_leaf_256_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_257_i_clk (.A(clknet_5_7_0_i_clk),
    .X(clknet_leaf_257_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_258_i_clk (.A(clknet_5_7_0_i_clk),
    .X(clknet_leaf_258_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_259_i_clk (.A(clknet_5_7_0_i_clk),
    .X(clknet_leaf_259_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_260_i_clk (.A(clknet_5_6_0_i_clk),
    .X(clknet_leaf_260_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_261_i_clk (.A(clknet_5_6_0_i_clk),
    .X(clknet_leaf_261_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_262_i_clk (.A(clknet_5_4_0_i_clk),
    .X(clknet_leaf_262_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_263_i_clk (.A(clknet_5_4_0_i_clk),
    .X(clknet_leaf_263_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_264_i_clk (.A(clknet_5_5_0_i_clk),
    .X(clknet_leaf_264_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_265_i_clk (.A(clknet_5_5_0_i_clk),
    .X(clknet_leaf_265_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_266_i_clk (.A(clknet_5_5_0_i_clk),
    .X(clknet_leaf_266_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_267_i_clk (.A(clknet_5_5_0_i_clk),
    .X(clknet_leaf_267_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_268_i_clk (.A(clknet_5_5_0_i_clk),
    .X(clknet_leaf_268_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_269_i_clk (.A(clknet_5_5_0_i_clk),
    .X(clknet_leaf_269_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_270_i_clk (.A(clknet_5_5_0_i_clk),
    .X(clknet_leaf_270_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_271_i_clk (.A(clknet_5_5_0_i_clk),
    .X(clknet_leaf_271_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_272_i_clk (.A(clknet_5_5_0_i_clk),
    .X(clknet_leaf_272_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_273_i_clk (.A(clknet_5_4_0_i_clk),
    .X(clknet_leaf_273_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_274_i_clk (.A(clknet_5_4_0_i_clk),
    .X(clknet_leaf_274_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_275_i_clk (.A(clknet_5_4_0_i_clk),
    .X(clknet_leaf_275_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_276_i_clk (.A(clknet_5_4_0_i_clk),
    .X(clknet_leaf_276_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_277_i_clk (.A(clknet_5_4_0_i_clk),
    .X(clknet_leaf_277_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_278_i_clk (.A(clknet_5_4_0_i_clk),
    .X(clknet_leaf_278_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_279_i_clk (.A(clknet_5_4_0_i_clk),
    .X(clknet_leaf_279_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_280_i_clk (.A(clknet_5_1_0_i_clk),
    .X(clknet_leaf_280_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_281_i_clk (.A(clknet_5_1_0_i_clk),
    .X(clknet_leaf_281_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_282_i_clk (.A(clknet_5_1_0_i_clk),
    .X(clknet_leaf_282_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_283_i_clk (.A(clknet_5_1_0_i_clk),
    .X(clknet_leaf_283_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_284_i_clk (.A(clknet_5_1_0_i_clk),
    .X(clknet_leaf_284_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_285_i_clk (.A(clknet_5_1_0_i_clk),
    .X(clknet_leaf_285_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_286_i_clk (.A(clknet_5_1_0_i_clk),
    .X(clknet_leaf_286_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_287_i_clk (.A(clknet_5_0_0_i_clk),
    .X(clknet_leaf_287_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_288_i_clk (.A(clknet_5_0_0_i_clk),
    .X(clknet_leaf_288_i_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_i_clk (.A(i_clk),
    .X(clknet_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_1_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_0_1_i_clk (.A(clknet_1_0_0_i_clk),
    .X(clknet_1_0_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_0_i_clk (.A(clknet_0_i_clk),
    .X(clknet_1_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_1_1_1_i_clk (.A(clknet_1_1_0_i_clk),
    .X(clknet_1_1_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_i_clk (.A(clknet_1_0_1_i_clk),
    .X(clknet_2_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_1_i_clk (.A(clknet_2_0_0_i_clk),
    .X(clknet_2_0_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_i_clk (.A(clknet_1_0_1_i_clk),
    .X(clknet_2_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_1_i_clk (.A(clknet_2_1_0_i_clk),
    .X(clknet_2_1_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_i_clk (.A(clknet_1_1_1_i_clk),
    .X(clknet_2_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_1_i_clk (.A(clknet_2_2_0_i_clk),
    .X(clknet_2_2_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_i_clk (.A(clknet_1_1_1_i_clk),
    .X(clknet_2_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_1_i_clk (.A(clknet_2_3_0_i_clk),
    .X(clknet_2_3_1_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_i_clk (.A(clknet_2_0_1_i_clk),
    .X(clknet_3_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_i_clk (.A(clknet_2_0_1_i_clk),
    .X(clknet_3_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_i_clk (.A(clknet_2_1_1_i_clk),
    .X(clknet_3_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_i_clk (.A(clknet_2_1_1_i_clk),
    .X(clknet_3_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_i_clk (.A(clknet_2_2_1_i_clk),
    .X(clknet_3_4_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_i_clk (.A(clknet_2_2_1_i_clk),
    .X(clknet_3_5_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_i_clk (.A(clknet_2_3_1_i_clk),
    .X(clknet_3_6_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_i_clk (.A(clknet_2_3_1_i_clk),
    .X(clknet_3_7_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_0_0_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_4_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_1_0_i_clk (.A(clknet_3_0_0_i_clk),
    .X(clknet_4_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_2_0_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_4_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_3_0_i_clk (.A(clknet_3_1_0_i_clk),
    .X(clknet_4_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_4_0_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_4_4_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_5_0_i_clk (.A(clknet_3_2_0_i_clk),
    .X(clknet_4_5_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_6_0_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_4_6_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_7_0_i_clk (.A(clknet_3_3_0_i_clk),
    .X(clknet_4_7_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_8_0_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_4_8_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_9_0_i_clk (.A(clknet_3_4_0_i_clk),
    .X(clknet_4_9_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_10_0_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_4_10_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_11_0_i_clk (.A(clknet_3_5_0_i_clk),
    .X(clknet_4_11_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_12_0_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_4_12_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_13_0_i_clk (.A(clknet_3_6_0_i_clk),
    .X(clknet_4_13_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_14_0_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_4_14_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_4_15_0_i_clk (.A(clknet_3_7_0_i_clk),
    .X(clknet_4_15_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_0_0_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_5_0_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_1_0_i_clk (.A(clknet_4_0_0_i_clk),
    .X(clknet_5_1_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_2_0_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_5_2_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_3_0_i_clk (.A(clknet_4_1_0_i_clk),
    .X(clknet_5_3_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_4_0_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_5_4_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_5_0_i_clk (.A(clknet_4_2_0_i_clk),
    .X(clknet_5_5_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_6_0_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_5_6_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_7_0_i_clk (.A(clknet_4_3_0_i_clk),
    .X(clknet_5_7_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_8_0_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_5_8_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_9_0_i_clk (.A(clknet_4_4_0_i_clk),
    .X(clknet_5_9_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_10_0_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_5_10_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_11_0_i_clk (.A(clknet_4_5_0_i_clk),
    .X(clknet_5_11_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_12_0_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_5_12_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_13_0_i_clk (.A(clknet_4_6_0_i_clk),
    .X(clknet_5_13_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_14_0_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_5_14_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_15_0_i_clk (.A(clknet_4_7_0_i_clk),
    .X(clknet_5_15_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_16_0_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_5_16_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_17_0_i_clk (.A(clknet_4_8_0_i_clk),
    .X(clknet_5_17_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_18_0_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_5_18_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_19_0_i_clk (.A(clknet_4_9_0_i_clk),
    .X(clknet_5_19_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_20_0_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_5_20_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_21_0_i_clk (.A(clknet_4_10_0_i_clk),
    .X(clknet_5_21_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_22_0_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_5_22_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_23_0_i_clk (.A(clknet_4_11_0_i_clk),
    .X(clknet_5_23_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_24_0_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_5_24_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_25_0_i_clk (.A(clknet_4_12_0_i_clk),
    .X(clknet_5_25_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_26_0_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_5_26_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_27_0_i_clk (.A(clknet_4_13_0_i_clk),
    .X(clknet_5_27_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_28_0_i_clk (.A(clknet_4_14_0_i_clk),
    .X(clknet_5_28_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_29_0_i_clk (.A(clknet_4_14_0_i_clk),
    .X(clknet_5_29_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_30_0_i_clk (.A(clknet_4_15_0_i_clk),
    .X(clknet_5_30_0_i_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_5_31_0_i_clk (.A(clknet_4_15_0_i_clk),
    .X(clknet_5_31_0_i_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\mem[42][7] ),
    .X(net41));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\mem[12][13] ),
    .X(net42));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\mem[120][4] ),
    .X(net43));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\mem[12][5] ),
    .X(net44));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\mem[9][5] ),
    .X(net45));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\mem[84][6] ),
    .X(net46));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\mem[97][12] ),
    .X(net47));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\mem[37][5] ),
    .X(net48));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\mem[76][5] ),
    .X(net49));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\mem[97][7] ),
    .X(net50));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\mem[37][6] ),
    .X(net51));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\mem[10][1] ),
    .X(net52));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\mem[33][14] ),
    .X(net53));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\mem[4][14] ),
    .X(net54));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\mem[68][4] ),
    .X(net55));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\mem[15][13] ),
    .X(net56));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\mem[97][11] ),
    .X(net57));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\mem[28][11] ),
    .X(net58));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\mem[20][2] ),
    .X(net59));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\mem[12][8] ),
    .X(net60));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\mem[68][11] ),
    .X(net61));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\mem[10][5] ),
    .X(net62));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\mem[35][13] ),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\mem[37][8] ),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\mem[76][8] ),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\mem[82][2] ),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\mem[76][15] ),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\mem[35][0] ),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\mem[68][10] ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\mem[20][8] ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\mem[84][7] ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\mem[48][14] ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\mem[12][12] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\mem[18][10] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\mem[68][9] ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\mem[113][1] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\mem[112][1] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\mem[72][13] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\mem[100][4] ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\mem[112][5] ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\mem[112][6] ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\mem[48][5] ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\mem[96][9] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\mem[41][12] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\mem[76][11] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\mem[48][0] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\mem[44][5] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\mem[28][15] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\mem[52][1] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\mem[114][13] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\mem[76][9] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\mem[12][6] ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\mem[8][7] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\mem[100][1] ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\mem[116][6] ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\mem[50][13] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\mem[104][5] ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\mem[112][10] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\mem[37][2] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\mem[12][4] ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\mem[20][1] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\mem[8][4] ),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\mem[37][1] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\mem[41][4] ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\mem[76][12] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\mem[20][4] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\mem[76][7] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\mem[72][8] ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\mem[74][10] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\mem[72][4] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\mem[113][10] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\mem[20][10] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\mem[33][12] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\mem[68][12] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\mem[84][8] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\mem[84][4] ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\mem[28][10] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\mem[37][3] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\mem[48][11] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\mem[74][14] ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\mem[82][4] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\mem[84][1] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\mem[35][14] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\mem[12][10] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\mem[50][8] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\mem[20][7] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\mem[84][13] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\mem[4][0] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\mem[20][11] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\mem[97][4] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\mem[104][4] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\mem[38][2] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\mem[45][3] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\mem[12][11] ),
    .X(net134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\mem[20][6] ),
    .X(net135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\mem[82][3] ),
    .X(net136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\mem[28][0] ),
    .X(net137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\mem[76][4] ),
    .X(net138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\mem[48][12] ),
    .X(net139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\mem[12][9] ),
    .X(net140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\mem[113][2] ),
    .X(net141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\mem[36][15] ),
    .X(net142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\mem[5][5] ),
    .X(net143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\mem[68][5] ),
    .X(net144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\mem[114][12] ),
    .X(net145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\mem[28][12] ),
    .X(net146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\mem[112][3] ),
    .X(net147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\mem[68][1] ),
    .X(net148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\mem[68][15] ),
    .X(net149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\mem[110][10] ),
    .X(net150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\mem[56][7] ),
    .X(net151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\mem[12][3] ),
    .X(net152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\mem[96][11] ),
    .X(net153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\mem[98][4] ),
    .X(net154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\mem[97][1] ),
    .X(net155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\mem[48][1] ),
    .X(net156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\mem[72][15] ),
    .X(net157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\mem[68][8] ),
    .X(net158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\mem[116][14] ),
    .X(net159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\mem[8][2] ),
    .X(net160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\mem[20][12] ),
    .X(net161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\mem[72][12] ),
    .X(net162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\mem[56][13] ),
    .X(net163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\mem[42][6] ),
    .X(net164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\mem[84][15] ),
    .X(net165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\mem[76][13] ),
    .X(net166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\mem[35][15] ),
    .X(net167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\mem[97][14] ),
    .X(net168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\mem[112][4] ),
    .X(net169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(\mem[4][11] ),
    .X(net170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\mem[74][0] ),
    .X(net171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\mem[52][11] ),
    .X(net172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(\mem[113][7] ),
    .X(net173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\mem[40][6] ),
    .X(net174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\mem[98][2] ),
    .X(net175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\mem[40][7] ),
    .X(net176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\mem[74][15] ),
    .X(net177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(\mem[44][0] ),
    .X(net178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\mem[42][0] ),
    .X(net179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\mem[10][6] ),
    .X(net180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(\mem[37][14] ),
    .X(net181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(\mem[72][14] ),
    .X(net182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\mem[48][8] ),
    .X(net183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\mem[68][6] ),
    .X(net184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\mem[20][3] ),
    .X(net185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(\mem[115][5] ),
    .X(net186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\mem[72][9] ),
    .X(net187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\mem[37][0] ),
    .X(net188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(\mem[74][11] ),
    .X(net189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\mem[76][10] ),
    .X(net190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\mem[20][15] ),
    .X(net191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(\mem[116][7] ),
    .X(net192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\mem[33][9] ),
    .X(net193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\mem[120][7] ),
    .X(net194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\mem[68][13] ),
    .X(net195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\mem[35][1] ),
    .X(net196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\mem[12][2] ),
    .X(net197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\mem[40][2] ),
    .X(net198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\mem[10][11] ),
    .X(net199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\mem[50][10] ),
    .X(net200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\mem[114][15] ),
    .X(net201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\mem[21][1] ),
    .X(net202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\mem[114][14] ),
    .X(net203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\mem[82][10] ),
    .X(net204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\mem[20][14] ),
    .X(net205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\mem[28][2] ),
    .X(net206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\mem[33][1] ),
    .X(net207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\mem[32][5] ),
    .X(net208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\mem[10][4] ),
    .X(net209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\mem[98][15] ),
    .X(net210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\mem[37][7] ),
    .X(net211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\mem[4][4] ),
    .X(net212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\mem[26][1] ),
    .X(net213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\mem[105][14] ),
    .X(net214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\mem[113][9] ),
    .X(net215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\mem[84][9] ),
    .X(net216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\mem[82][15] ),
    .X(net217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\mem[100][11] ),
    .X(net218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\mem[24][13] ),
    .X(net219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\mem[2][4] ),
    .X(net220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\mem[124][3] ),
    .X(net221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\mem[0][13] ),
    .X(net222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\mem[33][11] ),
    .X(net223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\mem[15][10] ),
    .X(net224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\mem[41][3] ),
    .X(net225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\mem[4][3] ),
    .X(net226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\mem[109][14] ),
    .X(net227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\mem[84][3] ),
    .X(net228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\mem[84][11] ),
    .X(net229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\mem[72][7] ),
    .X(net230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\mem[97][13] ),
    .X(net231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\mem[40][3] ),
    .X(net232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\mem[32][2] ),
    .X(net233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\mem[41][8] ),
    .X(net234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\mem[35][5] ),
    .X(net235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\mem[41][9] ),
    .X(net236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\mem[113][4] ),
    .X(net237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\mem[49][10] ),
    .X(net238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\mem[48][9] ),
    .X(net239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\mem[114][7] ),
    .X(net240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\mem[4][5] ),
    .X(net241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\mem[74][3] ),
    .X(net242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\mem[48][6] ),
    .X(net243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\mem[72][11] ),
    .X(net244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\mem[41][15] ),
    .X(net245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\mem[119][11] ),
    .X(net246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\mem[42][3] ),
    .X(net247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\mem[8][5] ),
    .X(net248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\mem[10][12] ),
    .X(net249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\mem[32][1] ),
    .X(net250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\mem[98][9] ),
    .X(net251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\mem[10][8] ),
    .X(net252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\mem[117][12] ),
    .X(net253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\mem[36][12] ),
    .X(net254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\mem[112][9] ),
    .X(net255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\mem[2][13] ),
    .X(net256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\mem[106][5] ),
    .X(net257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\mem[56][11] ),
    .X(net258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\mem[96][3] ),
    .X(net259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\mem[74][6] ),
    .X(net260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\mem[50][6] ),
    .X(net261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\mem[36][9] ),
    .X(net262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\mem[21][14] ),
    .X(net263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(\mem[114][8] ),
    .X(net264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(\mem[38][13] ),
    .X(net265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\mem[48][13] ),
    .X(net266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\mem[37][9] ),
    .X(net267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\mem[82][0] ),
    .X(net268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\mem[41][13] ),
    .X(net269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\mem[4][7] ),
    .X(net270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\mem[16][4] ),
    .X(net271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\mem[40][9] ),
    .X(net272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\mem[25][4] ),
    .X(net273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\mem[88][4] ),
    .X(net274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(\mem[39][6] ),
    .X(net275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(\mem[28][13] ),
    .X(net276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\mem[28][7] ),
    .X(net277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\mem[102][2] ),
    .X(net278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\mem[19][13] ),
    .X(net279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\mem[61][4] ),
    .X(net280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\mem[41][1] ),
    .X(net281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\mem[45][6] ),
    .X(net282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\mem[38][9] ),
    .X(net283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\mem[121][13] ),
    .X(net284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\mem[10][2] ),
    .X(net285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\mem[114][2] ),
    .X(net286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\mem[42][10] ),
    .X(net287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\mem[56][12] ),
    .X(net288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\mem[82][14] ),
    .X(net289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\mem[36][11] ),
    .X(net290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\mem[92][13] ),
    .X(net291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\mem[35][6] ),
    .X(net292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\mem[12][1] ),
    .X(net293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\mem[100][8] ),
    .X(net294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\mem[113][12] ),
    .X(net295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\mem[34][13] ),
    .X(net296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\mem[112][8] ),
    .X(net297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\mem[50][11] ),
    .X(net298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\mem[36][6] ),
    .X(net299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\mem[28][9] ),
    .X(net300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(\mem[42][8] ),
    .X(net301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\mem[33][0] ),
    .X(net302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\mem[120][10] ),
    .X(net303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\mem[47][10] ),
    .X(net304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\mem[8][8] ),
    .X(net305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\mem[17][10] ),
    .X(net306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\mem[127][15] ),
    .X(net307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\mem[114][9] ),
    .X(net308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(\mem[4][12] ),
    .X(net309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\mem[102][0] ),
    .X(net310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\mem[35][9] ),
    .X(net311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\mem[104][1] ),
    .X(net312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\mem[104][11] ),
    .X(net313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\mem[84][0] ),
    .X(net314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\mem[113][6] ),
    .X(net315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\mem[19][5] ),
    .X(net316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\mem[82][7] ),
    .X(net317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\mem[8][9] ),
    .X(net318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\mem[106][1] ),
    .X(net319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(\mem[50][5] ),
    .X(net320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(\mem[116][0] ),
    .X(net321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\mem[119][15] ),
    .X(net322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\mem[41][14] ),
    .X(net323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\mem[12][15] ),
    .X(net324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\mem[105][5] ),
    .X(net325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(\mem[50][12] ),
    .X(net326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\mem[74][2] ),
    .X(net327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\mem[10][10] ),
    .X(net328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\mem[114][4] ),
    .X(net329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\mem[55][8] ),
    .X(net330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\mem[64][2] ),
    .X(net331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(\mem[108][8] ),
    .X(net332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\mem[14][5] ),
    .X(net333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\mem[38][11] ),
    .X(net334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\mem[28][14] ),
    .X(net335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\mem[20][0] ),
    .X(net336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(\mem[44][15] ),
    .X(net337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\mem[42][5] ),
    .X(net338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\mem[52][14] ),
    .X(net339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(\mem[118][3] ),
    .X(net340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\mem[5][15] ),
    .X(net341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\mem[56][2] ),
    .X(net342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\mem[6][1] ),
    .X(net343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\mem[38][3] ),
    .X(net344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(\mem[100][2] ),
    .X(net345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\mem[92][2] ),
    .X(net346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\mem[52][15] ),
    .X(net347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\mem[125][3] ),
    .X(net348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\mem[56][10] ),
    .X(net349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(\mem[38][4] ),
    .X(net350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\mem[48][2] ),
    .X(net351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\mem[52][8] ),
    .X(net352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(\mem[97][15] ),
    .X(net353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\mem[34][3] ),
    .X(net354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\mem[72][1] ),
    .X(net355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\mem[64][13] ),
    .X(net356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\mem[1][10] ),
    .X(net357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\mem[97][0] ),
    .X(net358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\mem[84][12] ),
    .X(net359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(\mem[113][3] ),
    .X(net360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\mem[36][2] ),
    .X(net361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\mem[50][15] ),
    .X(net362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\mem[50][0] ),
    .X(net363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\mem[120][8] ),
    .X(net364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\mem[114][0] ),
    .X(net365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\mem[40][13] ),
    .X(net366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\mem[120][5] ),
    .X(net367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\mem[113][14] ),
    .X(net368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\mem[48][4] ),
    .X(net369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(\mem[26][5] ),
    .X(net370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(\mem[50][1] ),
    .X(net371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\mem[36][7] ),
    .X(net372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(\mem[76][6] ),
    .X(net373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(\mem[37][11] ),
    .X(net374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\mem[8][6] ),
    .X(net375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\mem[32][3] ),
    .X(net376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\mem[1][13] ),
    .X(net377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\mem[38][0] ),
    .X(net378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\mem[0][1] ),
    .X(net379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\mem[112][2] ),
    .X(net380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\mem[45][12] ),
    .X(net381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\mem[45][9] ),
    .X(net382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\mem[103][2] ),
    .X(net383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\mem[48][7] ),
    .X(net384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\mem[120][11] ),
    .X(net385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\mem[98][3] ),
    .X(net386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\mem[2][1] ),
    .X(net387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\mem[26][13] ),
    .X(net388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\mem[40][0] ),
    .X(net389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\mem[33][10] ),
    .X(net390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\mem[97][9] ),
    .X(net391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(\mem[4][10] ),
    .X(net392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\mem[61][7] ),
    .X(net393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\mem[45][15] ),
    .X(net394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\mem[20][13] ),
    .X(net395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\mem[120][14] ),
    .X(net396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\mem[21][2] ),
    .X(net397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\mem[42][9] ),
    .X(net398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\mem[12][7] ),
    .X(net399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\mem[41][10] ),
    .X(net400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\mem[10][7] ),
    .X(net401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\mem[44][12] ),
    .X(net402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\mem[53][7] ),
    .X(net403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\mem[50][14] ),
    .X(net404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\mem[96][4] ),
    .X(net405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\mem[68][7] ),
    .X(net406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\mem[126][11] ),
    .X(net407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\mem[113][0] ),
    .X(net408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\mem[73][0] ),
    .X(net409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\mem[125][14] ),
    .X(net410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\mem[52][13] ),
    .X(net411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\mem[38][1] ),
    .X(net412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\mem[114][11] ),
    .X(net413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\mem[113][13] ),
    .X(net414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\mem[4][2] ),
    .X(net415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\mem[33][5] ),
    .X(net416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\mem[37][10] ),
    .X(net417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\mem[73][7] ),
    .X(net418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\mem[37][4] ),
    .X(net419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\mem[113][11] ),
    .X(net420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\mem[107][4] ),
    .X(net421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\mem[76][3] ),
    .X(net422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\mem[121][0] ),
    .X(net423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\mem[61][11] ),
    .X(net424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\mem[92][3] ),
    .X(net425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\mem[116][12] ),
    .X(net426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\mem[97][8] ),
    .X(net427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\mem[38][6] ),
    .X(net428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\mem[96][8] ),
    .X(net429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\mem[112][7] ),
    .X(net430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(\mem[98][6] ),
    .X(net431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\mem[32][12] ),
    .X(net432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\mem[18][5] ),
    .X(net433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\mem[37][13] ),
    .X(net434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\mem[32][15] ),
    .X(net435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\mem[125][5] ),
    .X(net436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\mem[35][3] ),
    .X(net437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\mem[100][0] ),
    .X(net438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(\mem[82][5] ),
    .X(net439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(\mem[88][10] ),
    .X(net440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\mem[18][9] ),
    .X(net441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\mem[88][12] ),
    .X(net442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\mem[2][6] ),
    .X(net443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\mem[2][0] ),
    .X(net444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\mem[102][7] ),
    .X(net445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\mem[82][8] ),
    .X(net446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\mem[109][4] ),
    .X(net447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(\mem[113][15] ),
    .X(net448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\mem[123][13] ),
    .X(net449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(\mem[76][14] ),
    .X(net450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\mem[48][3] ),
    .X(net451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\mem[1][11] ),
    .X(net452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\mem[33][6] ),
    .X(net453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\mem[50][9] ),
    .X(net454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\mem[68][14] ),
    .X(net455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\mem[82][1] ),
    .X(net456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\mem[5][4] ),
    .X(net457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\mem[81][1] ),
    .X(net458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\mem[52][3] ),
    .X(net459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(\mem[18][0] ),
    .X(net460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\mem[0][3] ),
    .X(net461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(\mem[52][4] ),
    .X(net462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\mem[21][13] ),
    .X(net463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(\mem[41][11] ),
    .X(net464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\mem[20][9] ),
    .X(net465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(\mem[69][15] ),
    .X(net466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\mem[101][3] ),
    .X(net467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(\mem[16][10] ),
    .X(net468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\mem[40][12] ),
    .X(net469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\mem[1][6] ),
    .X(net470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\mem[38][12] ),
    .X(net471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(\mem[36][3] ),
    .X(net472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\mem[112][14] ),
    .X(net473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\mem[124][11] ),
    .X(net474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\mem[55][9] ),
    .X(net475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\mem[100][3] ),
    .X(net476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\mem[40][14] ),
    .X(net477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\mem[98][1] ),
    .X(net478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\mem[66][12] ),
    .X(net479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\mem[114][3] ),
    .X(net480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\mem[35][10] ),
    .X(net481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\mem[109][5] ),
    .X(net482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\mem[41][7] ),
    .X(net483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(\mem[33][8] ),
    .X(net484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\mem[18][12] ),
    .X(net485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\mem[105][11] ),
    .X(net486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\mem[44][14] ),
    .X(net487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(\mem[82][12] ),
    .X(net488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\mem[4][9] ),
    .X(net489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\mem[18][13] ),
    .X(net490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\mem[2][9] ),
    .X(net491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\mem[24][1] ),
    .X(net492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\mem[34][9] ),
    .X(net493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\mem[107][1] ),
    .X(net494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\mem[82][13] ),
    .X(net495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\mem[45][5] ),
    .X(net496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\mem[42][11] ),
    .X(net497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\mem[32][10] ),
    .X(net498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\mem[112][15] ),
    .X(net499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\mem[84][10] ),
    .X(net500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\mem[92][10] ),
    .X(net501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\mem[115][1] ),
    .X(net502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\mem[45][11] ),
    .X(net503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\mem[56][9] ),
    .X(net504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\mem[103][6] ),
    .X(net505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\mem[117][3] ),
    .X(net506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\mem[2][5] ),
    .X(net507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\mem[59][12] ),
    .X(net508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\mem[116][3] ),
    .X(net509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\mem[98][14] ),
    .X(net510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\mem[110][8] ),
    .X(net511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\mem[96][10] ),
    .X(net512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\mem[40][11] ),
    .X(net513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\mem[126][5] ),
    .X(net514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\mem[61][0] ),
    .X(net515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\mem[116][1] ),
    .X(net516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\mem[99][8] ),
    .X(net517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\mem[59][6] ),
    .X(net518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\mem[119][10] ),
    .X(net519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\mem[8][14] ),
    .X(net520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\mem[0][4] ),
    .X(net521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\mem[98][0] ),
    .X(net522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\mem[109][0] ),
    .X(net523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\mem[44][11] ),
    .X(net524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\mem[74][4] ),
    .X(net525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\mem[116][13] ),
    .X(net526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\mem[15][5] ),
    .X(net527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\mem[116][15] ),
    .X(net528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\mem[112][0] ),
    .X(net529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\mem[81][11] ),
    .X(net530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\mem[32][9] ),
    .X(net531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\mem[69][5] ),
    .X(net532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\mem[46][10] ),
    .X(net533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\mem[47][6] ),
    .X(net534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\mem[17][8] ),
    .X(net535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\mem[44][10] ),
    .X(net536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\mem[107][12] ),
    .X(net537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\mem[54][6] ),
    .X(net538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\mem[41][0] ),
    .X(net539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(\mem[113][5] ),
    .X(net540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\mem[96][13] ),
    .X(net541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(\mem[9][4] ),
    .X(net542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\mem[96][6] ),
    .X(net543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(\mem[55][13] ),
    .X(net544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\mem[107][5] ),
    .X(net545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\mem[47][4] ),
    .X(net546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\mem[5][3] ),
    .X(net547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\mem[53][5] ),
    .X(net548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\mem[122][12] ),
    .X(net549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\mem[0][14] ),
    .X(net550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\mem[99][6] ),
    .X(net551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\mem[2][8] ),
    .X(net552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\mem[124][5] ),
    .X(net553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\mem[13][1] ),
    .X(net554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\mem[10][9] ),
    .X(net555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(\mem[1][5] ),
    .X(net556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\mem[48][10] ),
    .X(net557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\mem[116][5] ),
    .X(net558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\mem[54][2] ),
    .X(net559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(\mem[100][6] ),
    .X(net560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\mem[109][8] ),
    .X(net561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(\mem[34][1] ),
    .X(net562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\mem[119][1] ),
    .X(net563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\mem[106][12] ),
    .X(net564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\mem[45][2] ),
    .X(net565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(\mem[122][14] ),
    .X(net566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\mem[121][3] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(\mem[126][13] ),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\mem[125][6] ),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(\mem[57][11] ),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\mem[57][15] ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(\mem[37][15] ),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\mem[116][9] ),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(\mem[9][9] ),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\mem[58][7] ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(\mem[35][2] ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\mem[67][11] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(\mem[80][15] ),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\mem[33][2] ),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(\mem[51][15] ),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\mem[4][8] ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(\mem[96][2] ),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\mem[21][3] ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(\mem[110][2] ),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\mem[10][3] ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(\mem[107][9] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\mem[19][7] ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(\mem[57][10] ),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(\mem[44][9] ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(\mem[120][13] ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\mem[100][14] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(\mem[117][0] ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\mem[100][15] ),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(\mem[73][13] ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\mem[28][1] ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(\mem[108][13] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\mem[96][15] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(\mem[43][15] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\mem[32][13] ),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(\mem[101][11] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\mem[114][10] ),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(\mem[114][6] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\mem[43][8] ),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(\mem[52][7] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\mem[127][6] ),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(\mem[56][6] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\mem[0][15] ),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(\mem[92][4] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\mem[60][12] ),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(\mem[53][9] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\mem[101][13] ),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(\mem[2][11] ),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\mem[4][13] ),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(\mem[110][14] ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\mem[61][9] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(\mem[45][0] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\mem[98][11] ),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(\mem[56][14] ),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\mem[100][7] ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(\mem[115][11] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\mem[96][0] ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(\mem[126][15] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\mem[112][13] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(\mem[124][13] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\mem[106][3] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(\mem[34][7] ),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\mem[107][11] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(\mem[96][7] ),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\mem[37][12] ),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(\mem[69][12] ),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(\mem[116][4] ),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(\mem[92][1] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\mem[127][7] ),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(\mem[58][11] ),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\mem[112][11] ),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(\mem[81][8] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\mem[124][8] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(\mem[61][1] ),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\mem[38][7] ),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(\mem[121][5] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\mem[126][10] ),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(\mem[65][2] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\mem[104][9] ),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(\mem[21][4] ),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\mem[105][0] ),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(\mem[43][0] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\mem[26][9] ),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(\mem[5][11] ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\mem[43][9] ),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(\mem[5][9] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\mem[18][14] ),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(\mem[70][15] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\mem[44][13] ),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(\mem[17][6] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\mem[16][11] ),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(\mem[113][8] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\mem[36][0] ),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(\mem[21][12] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\mem[40][8] ),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(\mem[15][1] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\mem[124][1] ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(\mem[101][9] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\mem[26][3] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(\mem[92][15] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\mem[76][0] ),
    .X(net665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(\mem[39][4] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\mem[125][10] ),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(\mem[74][13] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\mem[112][12] ),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(\mem[16][2] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\mem[66][1] ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(\mem[96][1] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\mem[70][13] ),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(\mem[114][1] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\mem[117][2] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(\mem[24][5] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\mem[125][15] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(\mem[46][6] ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\mem[72][5] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(\mem[16][7] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\mem[33][4] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(\mem[0][10] ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\mem[117][15] ),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(\mem[100][12] ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\mem[34][5] ),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(\mem[115][6] ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(\mem[62][4] ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(\mem[108][5] ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\mem[57][6] ),
    .X(net689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(\mem[99][15] ),
    .X(net690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold651 (.A(\mem[53][8] ),
    .X(net691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold652 (.A(\mem[49][11] ),
    .X(net692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold653 (.A(\mem[108][7] ),
    .X(net693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold654 (.A(\mem[81][7] ),
    .X(net694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold655 (.A(\mem[2][2] ),
    .X(net695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold656 (.A(\mem[58][12] ),
    .X(net696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold657 (.A(\mem[107][3] ),
    .X(net697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold658 (.A(\mem[0][2] ),
    .X(net698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold659 (.A(\mem[9][14] ),
    .X(net699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold660 (.A(\mem[121][11] ),
    .X(net700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold661 (.A(\mem[102][12] ),
    .X(net701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold662 (.A(\mem[103][14] ),
    .X(net702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold663 (.A(\mem[92][6] ),
    .X(net703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold664 (.A(\mem[73][12] ),
    .X(net704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold665 (.A(\mem[18][15] ),
    .X(net705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold666 (.A(\mem[122][15] ),
    .X(net706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold667 (.A(\mem[106][9] ),
    .X(net707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold668 (.A(\mem[73][14] ),
    .X(net708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold669 (.A(\mem[4][6] ),
    .X(net709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold670 (.A(\mem[98][8] ),
    .X(net710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold671 (.A(\mem[56][1] ),
    .X(net711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold672 (.A(\mem[60][8] ),
    .X(net712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold673 (.A(\mem[109][7] ),
    .X(net713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold674 (.A(\mem[50][7] ),
    .X(net714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold675 (.A(\mem[99][4] ),
    .X(net715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold676 (.A(\mem[116][11] ),
    .X(net716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold677 (.A(\mem[55][5] ),
    .X(net717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold678 (.A(\mem[118][12] ),
    .X(net718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold679 (.A(\mem[0][5] ),
    .X(net719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold680 (.A(\mem[62][7] ),
    .X(net720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold681 (.A(\mem[33][13] ),
    .X(net721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold682 (.A(\mem[35][11] ),
    .X(net722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold683 (.A(\mem[64][7] ),
    .X(net723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold684 (.A(\mem[88][7] ),
    .X(net724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold685 (.A(\mem[4][15] ),
    .X(net725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold686 (.A(\mem[51][2] ),
    .X(net726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold687 (.A(\mem[122][5] ),
    .X(net727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold688 (.A(\mem[118][13] ),
    .X(net728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold689 (.A(\mem[115][14] ),
    .X(net729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold690 (.A(\mem[45][7] ),
    .X(net730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold691 (.A(\mem[63][7] ),
    .X(net731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold692 (.A(\mem[40][1] ),
    .X(net732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold693 (.A(\mem[92][14] ),
    .X(net733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold694 (.A(\mem[41][6] ),
    .X(net734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold695 (.A(\mem[114][5] ),
    .X(net735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold696 (.A(\mem[84][14] ),
    .X(net736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold697 (.A(\mem[92][5] ),
    .X(net737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold698 (.A(\mem[51][4] ),
    .X(net738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold699 (.A(\mem[39][15] ),
    .X(net739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold700 (.A(\mem[122][7] ),
    .X(net740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold701 (.A(\mem[45][1] ),
    .X(net741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold702 (.A(\mem[60][10] ),
    .X(net742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold703 (.A(\mem[42][15] ),
    .X(net743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold704 (.A(\mem[119][13] ),
    .X(net744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold705 (.A(\mem[53][6] ),
    .X(net745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold706 (.A(\mem[67][5] ),
    .X(net746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold707 (.A(\mem[52][6] ),
    .X(net747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold708 (.A(\mem[52][9] ),
    .X(net748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold709 (.A(\mem[32][14] ),
    .X(net749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold710 (.A(\mem[8][1] ),
    .X(net750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold711 (.A(\mem[111][12] ),
    .X(net751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold712 (.A(\mem[63][14] ),
    .X(net752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold713 (.A(\mem[25][7] ),
    .X(net753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold714 (.A(\mem[102][10] ),
    .X(net754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold715 (.A(\mem[21][11] ),
    .X(net755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold716 (.A(\mem[52][12] ),
    .X(net756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold717 (.A(\mem[121][7] ),
    .X(net757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold718 (.A(\mem[41][2] ),
    .X(net758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold719 (.A(\mem[44][1] ),
    .X(net759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold720 (.A(\mem[100][9] ),
    .X(net760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold721 (.A(\mem[67][12] ),
    .X(net761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold722 (.A(\mem[73][9] ),
    .X(net762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold723 (.A(\mem[119][5] ),
    .X(net763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold724 (.A(\mem[61][5] ),
    .X(net764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold725 (.A(\mem[53][3] ),
    .X(net765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold726 (.A(\mem[11][1] ),
    .X(net766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold727 (.A(\mem[4][1] ),
    .X(net767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold728 (.A(\mem[110][3] ),
    .X(net768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold729 (.A(\mem[35][7] ),
    .X(net769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold730 (.A(\mem[124][4] ),
    .X(net770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold731 (.A(\mem[111][4] ),
    .X(net771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold732 (.A(\mem[51][13] ),
    .X(net772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold733 (.A(\mem[96][14] ),
    .X(net773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold734 (.A(\mem[120][6] ),
    .X(net774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold735 (.A(\mem[36][5] ),
    .X(net775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold736 (.A(\mem[63][1] ),
    .X(net776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold737 (.A(\mem[103][15] ),
    .X(net777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold738 (.A(\mem[127][8] ),
    .X(net778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold739 (.A(\mem[19][1] ),
    .X(net779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold740 (.A(\mem[66][13] ),
    .X(net780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold741 (.A(\mem[74][5] ),
    .X(net781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold742 (.A(\mem[90][7] ),
    .X(net782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold743 (.A(\mem[77][9] ),
    .X(net783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold744 (.A(\mem[107][10] ),
    .X(net784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold745 (.A(\mem[24][3] ),
    .X(net785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold746 (.A(\mem[43][14] ),
    .X(net786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold747 (.A(\mem[1][2] ),
    .X(net787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold748 (.A(\mem[67][10] ),
    .X(net788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold749 (.A(\mem[127][4] ),
    .X(net789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold750 (.A(\mem[101][4] ),
    .X(net790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold751 (.A(\mem[125][2] ),
    .X(net791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold752 (.A(\mem[115][10] ),
    .X(net792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold753 (.A(\mem[64][15] ),
    .X(net793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold754 (.A(\mem[25][3] ),
    .X(net794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold755 (.A(\mem[42][4] ),
    .X(net795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold756 (.A(\mem[124][7] ),
    .X(net796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold757 (.A(\mem[105][15] ),
    .X(net797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold758 (.A(\mem[70][10] ),
    .X(net798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold759 (.A(\mem[61][6] ),
    .X(net799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold760 (.A(\mem[121][14] ),
    .X(net800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold761 (.A(\mem[33][3] ),
    .X(net801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold762 (.A(\mem[26][0] ),
    .X(net802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold763 (.A(\mem[15][11] ),
    .X(net803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold764 (.A(\mem[53][11] ),
    .X(net804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold765 (.A(\mem[34][10] ),
    .X(net805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold766 (.A(\mem[120][2] ),
    .X(net806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold767 (.A(\mem[109][15] ),
    .X(net807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold768 (.A(\mem[9][13] ),
    .X(net808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold769 (.A(\mem[67][15] ),
    .X(net809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold770 (.A(\mem[15][9] ),
    .X(net810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold771 (.A(\mem[56][8] ),
    .X(net811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold772 (.A(\mem[62][11] ),
    .X(net812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold773 (.A(\mem[121][4] ),
    .X(net813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold774 (.A(\mem[31][12] ),
    .X(net814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold775 (.A(\mem[9][1] ),
    .X(net815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold776 (.A(\mem[9][15] ),
    .X(net816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold777 (.A(\mem[39][9] ),
    .X(net817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold778 (.A(\mem[118][7] ),
    .X(net818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold779 (.A(\mem[52][5] ),
    .X(net819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold780 (.A(\mem[50][3] ),
    .X(net820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold781 (.A(\mem[74][12] ),
    .X(net821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold782 (.A(\mem[27][13] ),
    .X(net822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold783 (.A(\mem[103][13] ),
    .X(net823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold784 (.A(\mem[29][6] ),
    .X(net824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold785 (.A(\mem[116][2] ),
    .X(net825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold786 (.A(\mem[2][7] ),
    .X(net826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold787 (.A(\mem[32][0] ),
    .X(net827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold788 (.A(\mem[18][2] ),
    .X(net828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold789 (.A(\mem[64][8] ),
    .X(net829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold790 (.A(\mem[15][12] ),
    .X(net830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold791 (.A(\mem[94][14] ),
    .X(net831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold792 (.A(\mem[19][10] ),
    .X(net832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold793 (.A(\mem[100][10] ),
    .X(net833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold794 (.A(\mem[65][4] ),
    .X(net834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold795 (.A(\mem[56][4] ),
    .X(net835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold796 (.A(\mem[115][0] ),
    .X(net836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold797 (.A(\mem[127][0] ),
    .X(net837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold798 (.A(\mem[77][15] ),
    .X(net838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold799 (.A(\mem[84][2] ),
    .X(net839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold800 (.A(\mem[44][4] ),
    .X(net840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold801 (.A(\mem[64][3] ),
    .X(net841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold802 (.A(\mem[105][12] ),
    .X(net842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold803 (.A(\mem[53][0] ),
    .X(net843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold804 (.A(\mem[81][4] ),
    .X(net844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold805 (.A(\mem[44][7] ),
    .X(net845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold806 (.A(\mem[26][7] ),
    .X(net846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold807 (.A(\mem[108][9] ),
    .X(net847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold808 (.A(\mem[82][11] ),
    .X(net848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold809 (.A(\mem[45][8] ),
    .X(net849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold810 (.A(\mem[40][5] ),
    .X(net850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold811 (.A(\mem[118][8] ),
    .X(net851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold812 (.A(\mem[17][1] ),
    .X(net852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold813 (.A(\mem[6][7] ),
    .X(net853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold814 (.A(\mem[101][14] ),
    .X(net854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold815 (.A(\mem[46][3] ),
    .X(net855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold816 (.A(\mem[46][8] ),
    .X(net856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold817 (.A(\mem[110][13] ),
    .X(net857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold818 (.A(\mem[57][7] ),
    .X(net858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold819 (.A(\mem[57][3] ),
    .X(net859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold820 (.A(\mem[64][11] ),
    .X(net860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold821 (.A(\mem[98][7] ),
    .X(net861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold822 (.A(\mem[57][4] ),
    .X(net862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold823 (.A(\mem[121][15] ),
    .X(net863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold824 (.A(\mem[28][3] ),
    .X(net864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold825 (.A(\mem[81][0] ),
    .X(net865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold826 (.A(\mem[5][12] ),
    .X(net866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold827 (.A(\mem[111][11] ),
    .X(net867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold828 (.A(\mem[124][12] ),
    .X(net868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold829 (.A(\mem[103][10] ),
    .X(net869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold830 (.A(\mem[22][6] ),
    .X(net870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold831 (.A(\mem[19][9] ),
    .X(net871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold832 (.A(\mem[110][9] ),
    .X(net872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold833 (.A(\mem[17][15] ),
    .X(net873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold834 (.A(\mem[81][15] ),
    .X(net874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold835 (.A(\mem[22][1] ),
    .X(net875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold836 (.A(\mem[54][12] ),
    .X(net876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold837 (.A(\mem[106][11] ),
    .X(net877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold838 (.A(\mem[122][3] ),
    .X(net878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold839 (.A(\mem[25][1] ),
    .X(net879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold840 (.A(\mem[47][15] ),
    .X(net880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold841 (.A(\mem[102][13] ),
    .X(net881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold842 (.A(\mem[18][11] ),
    .X(net882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold843 (.A(\mem[54][3] ),
    .X(net883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold844 (.A(\mem[103][4] ),
    .X(net884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold845 (.A(\mem[59][9] ),
    .X(net885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold846 (.A(\mem[35][4] ),
    .X(net886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold847 (.A(\mem[61][15] ),
    .X(net887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold848 (.A(\mem[122][11] ),
    .X(net888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold849 (.A(\mem[2][15] ),
    .X(net889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold850 (.A(\mem[66][11] ),
    .X(net890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold851 (.A(\mem[105][9] ),
    .X(net891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold852 (.A(\mem[57][2] ),
    .X(net892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold853 (.A(\mem[123][1] ),
    .X(net893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold854 (.A(\mem[21][15] ),
    .X(net894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold855 (.A(\mem[35][8] ),
    .X(net895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold856 (.A(\mem[0][0] ),
    .X(net896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold857 (.A(\mem[15][7] ),
    .X(net897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold858 (.A(\mem[111][1] ),
    .X(net898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold859 (.A(\mem[81][12] ),
    .X(net899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold860 (.A(\mem[107][7] ),
    .X(net900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold861 (.A(\mem[1][14] ),
    .X(net901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold862 (.A(\mem[18][1] ),
    .X(net902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold863 (.A(\mem[73][11] ),
    .X(net903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold864 (.A(\mem[44][2] ),
    .X(net904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold865 (.A(\mem[47][7] ),
    .X(net905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold866 (.A(\mem[43][13] ),
    .X(net906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold867 (.A(\mem[42][2] ),
    .X(net907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold868 (.A(\mem[46][0] ),
    .X(net908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold869 (.A(\mem[19][14] ),
    .X(net909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold870 (.A(\mem[89][7] ),
    .X(net910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold871 (.A(\mem[57][8] ),
    .X(net911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold872 (.A(\mem[6][15] ),
    .X(net912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold873 (.A(\mem[99][9] ),
    .X(net913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold874 (.A(\mem[10][14] ),
    .X(net914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold875 (.A(\mem[92][9] ),
    .X(net915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold876 (.A(\mem[26][10] ),
    .X(net916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold877 (.A(\mem[99][10] ),
    .X(net917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold878 (.A(\mem[107][6] ),
    .X(net918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold879 (.A(\mem[123][6] ),
    .X(net919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold880 (.A(\mem[100][13] ),
    .X(net920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold881 (.A(\mem[88][11] ),
    .X(net921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold882 (.A(\mem[111][3] ),
    .X(net922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold883 (.A(\mem[63][0] ),
    .X(net923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold884 (.A(\mem[127][9] ),
    .X(net924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold885 (.A(\mem[64][5] ),
    .X(net925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold886 (.A(\mem[22][7] ),
    .X(net926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold887 (.A(\mem[51][9] ),
    .X(net927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold888 (.A(\mem[96][12] ),
    .X(net928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold889 (.A(\mem[80][5] ),
    .X(net929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold890 (.A(\mem[126][4] ),
    .X(net930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold891 (.A(\mem[103][12] ),
    .X(net931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold892 (.A(\mem[1][3] ),
    .X(net932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold893 (.A(\mem[25][2] ),
    .X(net933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold894 (.A(\mem[63][12] ),
    .X(net934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold895 (.A(\mem[108][15] ),
    .X(net935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold896 (.A(\mem[17][12] ),
    .X(net936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold897 (.A(\mem[61][8] ),
    .X(net937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold898 (.A(\mem[0][9] ),
    .X(net938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold899 (.A(\mem[77][13] ),
    .X(net939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold900 (.A(\mem[99][1] ),
    .X(net940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold901 (.A(\mem[53][2] ),
    .X(net941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold902 (.A(\mem[55][10] ),
    .X(net942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold903 (.A(\mem[26][6] ),
    .X(net943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold904 (.A(\mem[111][15] ),
    .X(net944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold905 (.A(\mem[109][1] ),
    .X(net945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold906 (.A(\mem[66][8] ),
    .X(net946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold907 (.A(\mem[116][10] ),
    .X(net947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold908 (.A(\mem[88][8] ),
    .X(net948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold909 (.A(\mem[7][13] ),
    .X(net949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold910 (.A(\mem[45][4] ),
    .X(net950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold911 (.A(\mem[115][13] ),
    .X(net951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold912 (.A(\mem[13][12] ),
    .X(net952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold913 (.A(\mem[36][8] ),
    .X(net953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold914 (.A(\mem[48][15] ),
    .X(net954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold915 (.A(\mem[126][8] ),
    .X(net955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold916 (.A(\mem[1][1] ),
    .X(net956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold917 (.A(\mem[53][1] ),
    .X(net957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold918 (.A(\mem[115][2] ),
    .X(net958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold919 (.A(\mem[64][4] ),
    .X(net959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold920 (.A(\mem[28][4] ),
    .X(net960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold921 (.A(\mem[16][14] ),
    .X(net961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold922 (.A(\mem[101][15] ),
    .X(net962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold923 (.A(\mem[92][12] ),
    .X(net963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold924 (.A(\mem[103][5] ),
    .X(net964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold925 (.A(\mem[108][3] ),
    .X(net965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold926 (.A(\mem[117][9] ),
    .X(net966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold927 (.A(\mem[60][3] ),
    .X(net967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold928 (.A(\mem[70][11] ),
    .X(net968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold929 (.A(\mem[70][14] ),
    .X(net969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold930 (.A(\mem[115][3] ),
    .X(net970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold931 (.A(\mem[34][11] ),
    .X(net971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold932 (.A(\mem[105][6] ),
    .X(net972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold933 (.A(\mem[57][5] ),
    .X(net973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold934 (.A(\mem[54][0] ),
    .X(net974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold935 (.A(\mem[89][13] ),
    .X(net975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold936 (.A(\mem[36][10] ),
    .X(net976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold937 (.A(\mem[39][5] ),
    .X(net977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold938 (.A(\mem[57][13] ),
    .X(net978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold939 (.A(\mem[59][1] ),
    .X(net979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold940 (.A(\mem[21][8] ),
    .X(net980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold941 (.A(\mem[21][5] ),
    .X(net981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold942 (.A(\mem[51][10] ),
    .X(net982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold943 (.A(\mem[65][10] ),
    .X(net983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold944 (.A(\mem[103][0] ),
    .X(net984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold945 (.A(\mem[38][8] ),
    .X(net985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold946 (.A(\mem[46][13] ),
    .X(net986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold947 (.A(\mem[16][5] ),
    .X(net987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold948 (.A(\mem[65][6] ),
    .X(net988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold949 (.A(\mem[1][0] ),
    .X(net989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold950 (.A(\mem[52][2] ),
    .X(net990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold951 (.A(\mem[123][11] ),
    .X(net991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold952 (.A(\mem[6][12] ),
    .X(net992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold953 (.A(\mem[9][6] ),
    .X(net993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold954 (.A(\mem[9][7] ),
    .X(net994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold955 (.A(\mem[47][0] ),
    .X(net995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold956 (.A(\mem[64][14] ),
    .X(net996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold957 (.A(\mem[5][14] ),
    .X(net997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold958 (.A(\mem[1][9] ),
    .X(net998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold959 (.A(\mem[36][1] ),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold960 (.A(\mem[102][4] ),
    .X(net1000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold961 (.A(\mem[47][8] ),
    .X(net1001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold962 (.A(\mem[54][10] ),
    .X(net1002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold963 (.A(\mem[69][14] ),
    .X(net1003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold964 (.A(\mem[63][3] ),
    .X(net1004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold965 (.A(\mem[55][0] ),
    .X(net1005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold966 (.A(\mem[110][11] ),
    .X(net1006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold967 (.A(\mem[105][2] ),
    .X(net1007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold968 (.A(\mem[118][2] ),
    .X(net1008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold969 (.A(\mem[127][2] ),
    .X(net1009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold970 (.A(\mem[15][4] ),
    .X(net1010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold971 (.A(\mem[10][15] ),
    .X(net1011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold972 (.A(\mem[22][0] ),
    .X(net1012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold973 (.A(\mem[126][9] ),
    .X(net1013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold974 (.A(\mem[96][5] ),
    .X(net1014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold975 (.A(\mem[16][8] ),
    .X(net1015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold976 (.A(\mem[107][2] ),
    .X(net1016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold977 (.A(\mem[110][4] ),
    .X(net1017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold978 (.A(\mem[117][11] ),
    .X(net1018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold979 (.A(\mem[50][4] ),
    .X(net1019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold980 (.A(\mem[110][12] ),
    .X(net1020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold981 (.A(\mem[127][3] ),
    .X(net1021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold982 (.A(\mem[16][9] ),
    .X(net1022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold983 (.A(\mem[5][6] ),
    .X(net1023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold984 (.A(\mem[9][3] ),
    .X(net1024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold985 (.A(\mem[13][5] ),
    .X(net1025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold986 (.A(\mem[0][12] ),
    .X(net1026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold987 (.A(\mem[36][14] ),
    .X(net1027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold988 (.A(\mem[123][12] ),
    .X(net1028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold989 (.A(\mem[17][2] ),
    .X(net1029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold990 (.A(\mem[103][1] ),
    .X(net1030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold991 (.A(\mem[127][12] ),
    .X(net1031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold992 (.A(\mem[57][14] ),
    .X(net1032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold993 (.A(\mem[77][6] ),
    .X(net1033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold994 (.A(\mem[47][3] ),
    .X(net1034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold995 (.A(\mem[125][13] ),
    .X(net1035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold996 (.A(\mem[0][6] ),
    .X(net1036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold997 (.A(\mem[115][8] ),
    .X(net1037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold998 (.A(\mem[56][0] ),
    .X(net1038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold999 (.A(\mem[106][15] ),
    .X(net1039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1000 (.A(\mem[32][4] ),
    .X(net1040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1001 (.A(\mem[53][12] ),
    .X(net1041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1002 (.A(\mem[51][7] ),
    .X(net1042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1003 (.A(\mem[25][9] ),
    .X(net1043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1004 (.A(\mem[74][7] ),
    .X(net1044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1005 (.A(\mem[38][5] ),
    .X(net1045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1006 (.A(\mem[76][2] ),
    .X(net1046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1007 (.A(\mem[69][6] ),
    .X(net1047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1008 (.A(\mem[118][1] ),
    .X(net1048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1009 (.A(\mem[17][7] ),
    .X(net1049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1010 (.A(\mem[82][6] ),
    .X(net1050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1011 (.A(\mem[120][3] ),
    .X(net1051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1012 (.A(\mem[109][3] ),
    .X(net1052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1013 (.A(\mem[119][0] ),
    .X(net1053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1014 (.A(\mem[32][7] ),
    .X(net1054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1015 (.A(\mem[24][4] ),
    .X(net1055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1016 (.A(\mem[58][1] ),
    .X(net1056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1017 (.A(\mem[9][8] ),
    .X(net1057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1018 (.A(\mem[18][3] ),
    .X(net1058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1019 (.A(\mem[99][2] ),
    .X(net1059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1020 (.A(\mem[84][5] ),
    .X(net1060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1021 (.A(\mem[65][1] ),
    .X(net1061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1022 (.A(\mem[59][0] ),
    .X(net1062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1023 (.A(\mem[123][3] ),
    .X(net1063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1024 (.A(\mem[42][13] ),
    .X(net1064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1025 (.A(\mem[118][6] ),
    .X(net1065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1026 (.A(\mem[6][11] ),
    .X(net1066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1027 (.A(\mem[104][12] ),
    .X(net1067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1028 (.A(\mem[98][10] ),
    .X(net1068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1029 (.A(\mem[73][3] ),
    .X(net1069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1030 (.A(\mem[106][10] ),
    .X(net1070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1031 (.A(\mem[65][7] ),
    .X(net1071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1032 (.A(\mem[70][4] ),
    .X(net1072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1033 (.A(\mem[60][4] ),
    .X(net1073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1034 (.A(\mem[73][15] ),
    .X(net1074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1035 (.A(\mem[115][7] ),
    .X(net1075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1036 (.A(\mem[40][4] ),
    .X(net1076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1037 (.A(\mem[21][10] ),
    .X(net1077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1038 (.A(\mem[74][8] ),
    .X(net1078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1039 (.A(\mem[15][6] ),
    .X(net1079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1040 (.A(\mem[102][15] ),
    .X(net1080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1041 (.A(\mem[32][6] ),
    .X(net1081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1042 (.A(\mem[59][11] ),
    .X(net1082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1043 (.A(\mem[8][12] ),
    .X(net1083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1044 (.A(\mem[57][9] ),
    .X(net1084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1045 (.A(\mem[34][4] ),
    .X(net1085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1046 (.A(\mem[43][12] ),
    .X(net1086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1047 (.A(\mem[70][0] ),
    .X(net1087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1048 (.A(\mem[34][6] ),
    .X(net1088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1049 (.A(\mem[38][14] ),
    .X(net1089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1050 (.A(\mem[99][3] ),
    .X(net1090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1051 (.A(\mem[88][14] ),
    .X(net1091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1052 (.A(\mem[97][2] ),
    .X(net1092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1053 (.A(\mem[34][14] ),
    .X(net1093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1054 (.A(\mem[16][0] ),
    .X(net1094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1055 (.A(\mem[105][10] ),
    .X(net1095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1056 (.A(\mem[23][7] ),
    .X(net1096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1057 (.A(\mem[1][8] ),
    .X(net1097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1058 (.A(\mem[102][11] ),
    .X(net1098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1059 (.A(\mem[38][10] ),
    .X(net1099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1060 (.A(\mem[25][0] ),
    .X(net1100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1061 (.A(\mem[5][13] ),
    .X(net1101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1062 (.A(\mem[59][4] ),
    .X(net1102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1063 (.A(\mem[92][7] ),
    .X(net1103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1064 (.A(\mem[13][9] ),
    .X(net1104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1065 (.A(\mem[88][6] ),
    .X(net1105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1066 (.A(\mem[121][2] ),
    .X(net1106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1067 (.A(\mem[36][13] ),
    .X(net1107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1068 (.A(\mem[85][8] ),
    .X(net1108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1069 (.A(\mem[24][7] ),
    .X(net1109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1070 (.A(\mem[18][7] ),
    .X(net1110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1071 (.A(\mem[65][8] ),
    .X(net1111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1072 (.A(\mem[66][0] ),
    .X(net1112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1073 (.A(\mem[24][8] ),
    .X(net1113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1074 (.A(\mem[12][14] ),
    .X(net1114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1075 (.A(\mem[122][1] ),
    .X(net1115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1076 (.A(\mem[119][8] ),
    .X(net1116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1077 (.A(\mem[81][2] ),
    .X(net1117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1078 (.A(\mem[117][6] ),
    .X(net1118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1079 (.A(\mem[73][10] ),
    .X(net1119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1080 (.A(\mem[111][10] ),
    .X(net1120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1081 (.A(\mem[97][3] ),
    .X(net1121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1082 (.A(\mem[90][9] ),
    .X(net1122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1083 (.A(\mem[54][5] ),
    .X(net1123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1084 (.A(\mem[52][0] ),
    .X(net1124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1085 (.A(\mem[46][7] ),
    .X(net1125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1086 (.A(\mem[27][2] ),
    .X(net1126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1087 (.A(\mem[22][12] ),
    .X(net1127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1088 (.A(\mem[70][1] ),
    .X(net1128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1089 (.A(\mem[65][9] ),
    .X(net1129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1090 (.A(\mem[24][15] ),
    .X(net1130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1091 (.A(\mem[122][0] ),
    .X(net1131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1092 (.A(\mem[118][0] ),
    .X(net1132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1093 (.A(\mem[124][2] ),
    .X(net1133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1094 (.A(\mem[123][8] ),
    .X(net1134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1095 (.A(\mem[5][8] ),
    .X(net1135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1096 (.A(\mem[125][1] ),
    .X(net1136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1097 (.A(\mem[72][10] ),
    .X(net1137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1098 (.A(\mem[16][13] ),
    .X(net1138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1099 (.A(\mem[54][11] ),
    .X(net1139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1100 (.A(\mem[70][8] ),
    .X(net1140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1101 (.A(\mem[57][12] ),
    .X(net1141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1102 (.A(\mem[102][8] ),
    .X(net1142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1103 (.A(\mem[105][1] ),
    .X(net1143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1104 (.A(\mem[103][7] ),
    .X(net1144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1105 (.A(\mem[117][4] ),
    .X(net1145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1106 (.A(\mem[47][12] ),
    .X(net1146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1107 (.A(\mem[43][6] ),
    .X(net1147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1108 (.A(\mem[51][11] ),
    .X(net1148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1109 (.A(\mem[67][6] ),
    .X(net1149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1110 (.A(\mem[7][3] ),
    .X(net1150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1111 (.A(\mem[119][2] ),
    .X(net1151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1112 (.A(\mem[22][15] ),
    .X(net1152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1113 (.A(\mem[80][3] ),
    .X(net1153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1114 (.A(\mem[53][4] ),
    .X(net1154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1115 (.A(\mem[77][2] ),
    .X(net1155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1116 (.A(\mem[97][6] ),
    .X(net1156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1117 (.A(\mem[90][12] ),
    .X(net1157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1118 (.A(\mem[116][8] ),
    .X(net1158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1119 (.A(\mem[111][9] ),
    .X(net1159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1120 (.A(\mem[106][6] ),
    .X(net1160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1121 (.A(\mem[89][10] ),
    .X(net1161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1122 (.A(\mem[2][12] ),
    .X(net1162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1123 (.A(\mem[29][5] ),
    .X(net1163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1124 (.A(\mem[15][15] ),
    .X(net1164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1125 (.A(\mem[56][5] ),
    .X(net1165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1126 (.A(\mem[70][7] ),
    .X(net1166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1127 (.A(\mem[94][5] ),
    .X(net1167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1128 (.A(\mem[43][11] ),
    .X(net1168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1129 (.A(\mem[120][12] ),
    .X(net1169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1130 (.A(\mem[88][0] ),
    .X(net1170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1131 (.A(\mem[54][14] ),
    .X(net1171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1132 (.A(\mem[124][10] ),
    .X(net1172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1133 (.A(\mem[17][11] ),
    .X(net1173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1134 (.A(\mem[95][13] ),
    .X(net1174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1135 (.A(\mem[7][14] ),
    .X(net1175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1136 (.A(\mem[60][15] ),
    .X(net1176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1137 (.A(\mem[26][4] ),
    .X(net1177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1138 (.A(\mem[88][2] ),
    .X(net1178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1139 (.A(\mem[109][11] ),
    .X(net1179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1140 (.A(\mem[6][13] ),
    .X(net1180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1141 (.A(\mem[97][10] ),
    .X(net1181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1142 (.A(\mem[17][3] ),
    .X(net1182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1143 (.A(\mem[64][0] ),
    .X(net1183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1144 (.A(\mem[39][3] ),
    .X(net1184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1145 (.A(\mem[119][7] ),
    .X(net1185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1146 (.A(\mem[16][12] ),
    .X(net1186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1147 (.A(\mem[101][8] ),
    .X(net1187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1148 (.A(\mem[79][4] ),
    .X(net1188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1149 (.A(\mem[59][3] ),
    .X(net1189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1150 (.A(\mem[46][4] ),
    .X(net1190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1151 (.A(\mem[81][10] ),
    .X(net1191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1152 (.A(\mem[61][3] ),
    .X(net1192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1153 (.A(\mem[108][14] ),
    .X(net1193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1154 (.A(\mem[124][15] ),
    .X(net1194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1155 (.A(\mem[46][12] ),
    .X(net1195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1156 (.A(\mem[89][0] ),
    .X(net1196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1157 (.A(\mem[61][14] ),
    .X(net1197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1158 (.A(\mem[107][8] ),
    .X(net1198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1159 (.A(\mem[33][15] ),
    .X(net1199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1160 (.A(\mem[88][3] ),
    .X(net1200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1161 (.A(\mem[124][14] ),
    .X(net1201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1162 (.A(\mem[123][5] ),
    .X(net1202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1163 (.A(\mem[127][13] ),
    .X(net1203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1164 (.A(\mem[118][9] ),
    .X(net1204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1165 (.A(\mem[90][4] ),
    .X(net1205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1166 (.A(\mem[105][13] ),
    .X(net1206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1167 (.A(\mem[69][11] ),
    .X(net1207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1168 (.A(\mem[70][3] ),
    .X(net1208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1169 (.A(\mem[80][0] ),
    .X(net1209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1170 (.A(\mem[125][11] ),
    .X(net1210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1171 (.A(\mem[76][1] ),
    .X(net1211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1172 (.A(\mem[64][10] ),
    .X(net1212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1173 (.A(\mem[79][5] ),
    .X(net1213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1174 (.A(\mem[126][6] ),
    .X(net1214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1175 (.A(\mem[62][5] ),
    .X(net1215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1176 (.A(\mem[85][7] ),
    .X(net1216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1177 (.A(\mem[74][9] ),
    .X(net1217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1178 (.A(\mem[11][9] ),
    .X(net1218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1179 (.A(\mem[16][3] ),
    .X(net1219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1180 (.A(\mem[109][2] ),
    .X(net1220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1181 (.A(\mem[39][13] ),
    .X(net1221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1182 (.A(\mem[60][1] ),
    .X(net1222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1183 (.A(\mem[36][4] ),
    .X(net1223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1184 (.A(\mem[106][14] ),
    .X(net1224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1185 (.A(\mem[21][9] ),
    .X(net1225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1186 (.A(\mem[121][6] ),
    .X(net1226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1187 (.A(\mem[59][15] ),
    .X(net1227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1188 (.A(\mem[62][12] ),
    .X(net1228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1189 (.A(\mem[30][14] ),
    .X(net1229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1190 (.A(\mem[15][2] ),
    .X(net1230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1191 (.A(\mem[92][8] ),
    .X(net1231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1192 (.A(\mem[73][5] ),
    .X(net1232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1193 (.A(\mem[5][7] ),
    .X(net1233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1194 (.A(\mem[39][1] ),
    .X(net1234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1195 (.A(\mem[108][1] ),
    .X(net1235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1196 (.A(\mem[60][7] ),
    .X(net1236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1197 (.A(\mem[117][1] ),
    .X(net1237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1198 (.A(\mem[93][6] ),
    .X(net1238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1199 (.A(\mem[55][7] ),
    .X(net1239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1200 (.A(\mem[31][6] ),
    .X(net1240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1201 (.A(\mem[93][7] ),
    .X(net1241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1202 (.A(\mem[103][9] ),
    .X(net1242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1203 (.A(\mem[73][2] ),
    .X(net1243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1204 (.A(\mem[108][2] ),
    .X(net1244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1205 (.A(\mem[98][12] ),
    .X(net1245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1206 (.A(\mem[64][9] ),
    .X(net1246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1207 (.A(\mem[47][9] ),
    .X(net1247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1208 (.A(\mem[8][0] ),
    .X(net1248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1209 (.A(\mem[67][1] ),
    .X(net1249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1210 (.A(\mem[125][8] ),
    .X(net1250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1211 (.A(\mem[110][1] ),
    .X(net1251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1212 (.A(\mem[26][14] ),
    .X(net1252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1213 (.A(\mem[118][15] ),
    .X(net1253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1214 (.A(\mem[46][1] ),
    .X(net1254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1215 (.A(\mem[127][1] ),
    .X(net1255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1216 (.A(\mem[105][7] ),
    .X(net1256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1217 (.A(\mem[32][11] ),
    .X(net1257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1218 (.A(\mem[62][10] ),
    .X(net1258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1219 (.A(\mem[67][13] ),
    .X(net1259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1220 (.A(\mem[42][1] ),
    .X(net1260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1221 (.A(\mem[111][14] ),
    .X(net1261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1222 (.A(\mem[125][9] ),
    .X(net1262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1223 (.A(\mem[119][9] ),
    .X(net1263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1224 (.A(\mem[88][15] ),
    .X(net1264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1225 (.A(\mem[1][15] ),
    .X(net1265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1226 (.A(\mem[110][5] ),
    .X(net1266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1227 (.A(\mem[81][14] ),
    .X(net1267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1228 (.A(\mem[62][3] ),
    .X(net1268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1229 (.A(\mem[126][7] ),
    .X(net1269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1230 (.A(\mem[77][12] ),
    .X(net1270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1231 (.A(\mem[67][14] ),
    .X(net1271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1232 (.A(\mem[24][9] ),
    .X(net1272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1233 (.A(\mem[23][1] ),
    .X(net1273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1234 (.A(\mem[88][13] ),
    .X(net1274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1235 (.A(\mem[78][12] ),
    .X(net1275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1236 (.A(\mem[53][13] ),
    .X(net1276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1237 (.A(\mem[78][15] ),
    .X(net1277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1238 (.A(\mem[101][10] ),
    .X(net1278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1239 (.A(\mem[34][8] ),
    .X(net1279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1240 (.A(\mem[101][12] ),
    .X(net1280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1241 (.A(\mem[108][4] ),
    .X(net1281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1242 (.A(\mem[103][3] ),
    .X(net1282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1243 (.A(\mem[22][10] ),
    .X(net1283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1244 (.A(\mem[122][10] ),
    .X(net1284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1245 (.A(\mem[90][10] ),
    .X(net1285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1246 (.A(\mem[126][3] ),
    .X(net1286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1247 (.A(\mem[108][12] ),
    .X(net1287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1248 (.A(\mem[67][9] ),
    .X(net1288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1249 (.A(\mem[51][1] ),
    .X(net1289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1250 (.A(\mem[0][7] ),
    .X(net1290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1251 (.A(\mem[15][14] ),
    .X(net1291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1252 (.A(\mem[22][4] ),
    .X(net1292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1253 (.A(\mem[6][9] ),
    .X(net1293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1254 (.A(\mem[64][6] ),
    .X(net1294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1255 (.A(\mem[63][8] ),
    .X(net1295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1256 (.A(\mem[51][3] ),
    .X(net1296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1257 (.A(\mem[5][10] ),
    .X(net1297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1258 (.A(\mem[125][0] ),
    .X(net1298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1259 (.A(\mem[66][15] ),
    .X(net1299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1260 (.A(\mem[34][0] ),
    .X(net1300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1261 (.A(\mem[60][2] ),
    .X(net1301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1262 (.A(\mem[63][9] ),
    .X(net1302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1263 (.A(\mem[60][5] ),
    .X(net1303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1264 (.A(\mem[107][15] ),
    .X(net1304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1265 (.A(\mem[19][6] ),
    .X(net1305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1266 (.A(\mem[28][5] ),
    .X(net1306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1267 (.A(\mem[81][9] ),
    .X(net1307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1268 (.A(\mem[14][1] ),
    .X(net1308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1269 (.A(\mem[107][0] ),
    .X(net1309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1270 (.A(\mem[87][4] ),
    .X(net1310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1271 (.A(\mem[13][6] ),
    .X(net1311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1272 (.A(\mem[10][13] ),
    .X(net1312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1273 (.A(\mem[66][9] ),
    .X(net1313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1274 (.A(\mem[57][0] ),
    .X(net1314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1275 (.A(\mem[26][15] ),
    .X(net1315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1276 (.A(\mem[91][15] ),
    .X(net1316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1277 (.A(\mem[79][6] ),
    .X(net1317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1278 (.A(\mem[19][15] ),
    .X(net1318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1279 (.A(\mem[59][13] ),
    .X(net1319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1280 (.A(\mem[70][6] ),
    .X(net1320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1281 (.A(\mem[70][2] ),
    .X(net1321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1282 (.A(\mem[73][6] ),
    .X(net1322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1283 (.A(\mem[103][8] ),
    .X(net1323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1284 (.A(\mem[22][13] ),
    .X(net1324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1285 (.A(\mem[13][3] ),
    .X(net1325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1286 (.A(\mem[107][13] ),
    .X(net1326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1287 (.A(\mem[46][15] ),
    .X(net1327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1288 (.A(\mem[74][1] ),
    .X(net1328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1289 (.A(\mem[31][2] ),
    .X(net1329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1290 (.A(\mem[16][1] ),
    .X(net1330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1291 (.A(\mem[40][10] ),
    .X(net1331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1292 (.A(\mem[104][10] ),
    .X(net1332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1293 (.A(\mem[115][12] ),
    .X(net1333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1294 (.A(\mem[7][4] ),
    .X(net1334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1295 (.A(\mem[79][7] ),
    .X(net1335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1296 (.A(\mem[25][11] ),
    .X(net1336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1297 (.A(\mem[62][9] ),
    .X(net1337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1298 (.A(\mem[105][8] ),
    .X(net1338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1299 (.A(\mem[126][14] ),
    .X(net1339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1300 (.A(\mem[123][14] ),
    .X(net1340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1301 (.A(\mem[117][10] ),
    .X(net1341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1302 (.A(\mem[63][5] ),
    .X(net1342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1303 (.A(\mem[95][0] ),
    .X(net1343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1304 (.A(\mem[119][14] ),
    .X(net1344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1305 (.A(\mem[8][10] ),
    .X(net1345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1306 (.A(\mem[106][7] ),
    .X(net1346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1307 (.A(\mem[25][5] ),
    .X(net1347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1308 (.A(\mem[13][0] ),
    .X(net1348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1309 (.A(\mem[100][5] ),
    .X(net1349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1310 (.A(\mem[43][2] ),
    .X(net1350));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1311 (.A(\mem[6][14] ),
    .X(net1351));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1312 (.A(\mem[46][5] ),
    .X(net1352));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1313 (.A(\mem[65][0] ),
    .X(net1353));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1314 (.A(\mem[122][2] ),
    .X(net1354));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1315 (.A(\mem[17][0] ),
    .X(net1355));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1316 (.A(\mem[22][3] ),
    .X(net1356));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1317 (.A(\mem[123][0] ),
    .X(net1357));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1318 (.A(\mem[66][10] ),
    .X(net1358));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1319 (.A(\mem[122][13] ),
    .X(net1359));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1320 (.A(\mem[124][6] ),
    .X(net1360));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1321 (.A(\mem[57][1] ),
    .X(net1361));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1322 (.A(\mem[87][11] ),
    .X(net1362));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1323 (.A(\mem[104][3] ),
    .X(net1363));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1324 (.A(\mem[44][6] ),
    .X(net1364));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1325 (.A(\mem[121][8] ),
    .X(net1365));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1326 (.A(\mem[60][0] ),
    .X(net1366));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1327 (.A(\mem[14][13] ),
    .X(net1367));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1328 (.A(\mem[64][12] ),
    .X(net1368));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1329 (.A(\mem[119][3] ),
    .X(net1369));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1330 (.A(\mem[127][14] ),
    .X(net1370));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1331 (.A(\mem[59][5] ),
    .X(net1371));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1332 (.A(\mem[42][12] ),
    .X(net1372));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1333 (.A(\mem[6][8] ),
    .X(net1373));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1334 (.A(\mem[101][7] ),
    .X(net1374));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1335 (.A(\mem[93][13] ),
    .X(net1375));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1336 (.A(\mem[127][10] ),
    .X(net1376));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1337 (.A(\mem[58][15] ),
    .X(net1377));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1338 (.A(\mem[93][2] ),
    .X(net1378));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1339 (.A(\mem[111][7] ),
    .X(net1379));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1340 (.A(\mem[29][9] ),
    .X(net1380));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1341 (.A(\mem[118][10] ),
    .X(net1381));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1342 (.A(\mem[32][8] ),
    .X(net1382));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1343 (.A(\mem[99][5] ),
    .X(net1383));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1344 (.A(\mem[31][7] ),
    .X(net1384));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1345 (.A(\mem[14][10] ),
    .X(net1385));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1346 (.A(\mem[121][9] ),
    .X(net1386));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1347 (.A(\mem[22][8] ),
    .X(net1387));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1348 (.A(\mem[31][11] ),
    .X(net1388));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1349 (.A(\mem[122][8] ),
    .X(net1389));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1350 (.A(\mem[86][10] ),
    .X(net1390));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1351 (.A(\mem[59][8] ),
    .X(net1391));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1352 (.A(\mem[22][11] ),
    .X(net1392));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1353 (.A(\mem[43][7] ),
    .X(net1393));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1354 (.A(\mem[60][11] ),
    .X(net1394));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1355 (.A(\mem[118][11] ),
    .X(net1395));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1356 (.A(\mem[109][6] ),
    .X(net1396));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1357 (.A(\mem[9][11] ),
    .X(net1397));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1358 (.A(\mem[16][6] ),
    .X(net1398));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1359 (.A(\mem[123][15] ),
    .X(net1399));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1360 (.A(\mem[29][1] ),
    .X(net1400));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1361 (.A(\mem[103][11] ),
    .X(net1401));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1362 (.A(\mem[60][14] ),
    .X(net1402));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1363 (.A(\mem[39][11] ),
    .X(net1403));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1364 (.A(\mem[43][4] ),
    .X(net1404));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1365 (.A(\mem[5][2] ),
    .X(net1405));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1366 (.A(\mem[14][6] ),
    .X(net1406));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1367 (.A(\mem[61][13] ),
    .X(net1407));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1368 (.A(\mem[106][2] ),
    .X(net1408));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1369 (.A(\mem[107][14] ),
    .X(net1409));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1370 (.A(\mem[91][3] ),
    .X(net1410));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1371 (.A(\mem[123][4] ),
    .X(net1411));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1372 (.A(\mem[66][5] ),
    .X(net1412));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1373 (.A(\mem[117][8] ),
    .X(net1413));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1374 (.A(\mem[118][4] ),
    .X(net1414));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1375 (.A(\mem[106][8] ),
    .X(net1415));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1376 (.A(\mem[75][8] ),
    .X(net1416));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1377 (.A(\mem[30][9] ),
    .X(net1417));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1378 (.A(\mem[68][3] ),
    .X(net1418));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1379 (.A(\mem[85][12] ),
    .X(net1419));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1380 (.A(\mem[62][8] ),
    .X(net1420));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1381 (.A(\mem[58][6] ),
    .X(net1421));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1382 (.A(\mem[25][8] ),
    .X(net1422));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1383 (.A(\mem[99][0] ),
    .X(net1423));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1384 (.A(\mem[59][14] ),
    .X(net1424));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1385 (.A(\mem[123][2] ),
    .X(net1425));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1386 (.A(\mem[117][13] ),
    .X(net1426));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1387 (.A(\mem[85][0] ),
    .X(net1427));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1388 (.A(\mem[77][5] ),
    .X(net1428));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1389 (.A(\mem[0][11] ),
    .X(net1429));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1390 (.A(\mem[58][0] ),
    .X(net1430));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1391 (.A(\mem[120][1] ),
    .X(net1431));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1392 (.A(\mem[73][4] ),
    .X(net1432));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1393 (.A(\mem[95][11] ),
    .X(net1433));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1394 (.A(\mem[29][3] ),
    .X(net1434));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1395 (.A(\mem[69][13] ),
    .X(net1435));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1396 (.A(\mem[28][8] ),
    .X(net1436));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1397 (.A(\mem[34][15] ),
    .X(net1437));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1398 (.A(\mem[16][15] ),
    .X(net1438));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1399 (.A(\mem[44][3] ),
    .X(net1439));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1400 (.A(\mem[120][0] ),
    .X(net1440));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1401 (.A(\mem[95][14] ),
    .X(net1441));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1402 (.A(\mem[110][7] ),
    .X(net1442));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1403 (.A(\mem[120][9] ),
    .X(net1443));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1404 (.A(\mem[15][3] ),
    .X(net1444));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1405 (.A(\mem[66][14] ),
    .X(net1445));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1406 (.A(\mem[43][5] ),
    .X(net1446));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1407 (.A(\mem[80][9] ),
    .X(net1447));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1408 (.A(\mem[64][1] ),
    .X(net1448));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1409 (.A(\mem[31][1] ),
    .X(net1449));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1410 (.A(\mem[5][1] ),
    .X(net1450));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1411 (.A(\mem[109][13] ),
    .X(net1451));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1412 (.A(\mem[19][11] ),
    .X(net1452));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1413 (.A(\mem[63][2] ),
    .X(net1453));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1414 (.A(\mem[70][12] ),
    .X(net1454));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1415 (.A(\mem[66][3] ),
    .X(net1455));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1416 (.A(\mem[98][5] ),
    .X(net1456));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1417 (.A(\mem[34][2] ),
    .X(net1457));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1418 (.A(\mem[75][7] ),
    .X(net1458));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1419 (.A(\mem[27][9] ),
    .X(net1459));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1420 (.A(\mem[82][9] ),
    .X(net1460));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1421 (.A(\mem[63][10] ),
    .X(net1461));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1422 (.A(\mem[86][0] ),
    .X(net1462));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1423 (.A(\mem[102][3] ),
    .X(net1463));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1424 (.A(\mem[71][6] ),
    .X(net1464));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1425 (.A(\mem[53][14] ),
    .X(net1465));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1426 (.A(\mem[2][10] ),
    .X(net1466));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1427 (.A(\mem[58][10] ),
    .X(net1467));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1428 (.A(\mem[125][7] ),
    .X(net1468));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1429 (.A(\mem[89][8] ),
    .X(net1469));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1430 (.A(\mem[22][2] ),
    .X(net1470));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1431 (.A(\mem[46][9] ),
    .X(net1471));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1432 (.A(\mem[25][13] ),
    .X(net1472));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1433 (.A(\mem[87][7] ),
    .X(net1473));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1434 (.A(\mem[93][15] ),
    .X(net1474));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1435 (.A(\mem[90][11] ),
    .X(net1475));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1436 (.A(\mem[58][9] ),
    .X(net1476));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1437 (.A(\mem[87][12] ),
    .X(net1477));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1438 (.A(\mem[127][5] ),
    .X(net1478));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1439 (.A(\mem[95][7] ),
    .X(net1479));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1440 (.A(\mem[65][14] ),
    .X(net1480));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1441 (.A(\mem[24][0] ),
    .X(net1481));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1442 (.A(\mem[53][10] ),
    .X(net1482));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1443 (.A(\mem[23][4] ),
    .X(net1483));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1444 (.A(\mem[81][3] ),
    .X(net1484));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1445 (.A(\mem[55][4] ),
    .X(net1485));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1446 (.A(\mem[58][14] ),
    .X(net1486));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1447 (.A(\mem[13][2] ),
    .X(net1487));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1448 (.A(\mem[89][11] ),
    .X(net1488));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1449 (.A(\mem[60][13] ),
    .X(net1489));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1450 (.A(\mem[78][11] ),
    .X(net1490));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1451 (.A(\mem[9][12] ),
    .X(net1491));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1452 (.A(\mem[46][14] ),
    .X(net1492));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1453 (.A(\mem[27][6] ),
    .X(net1493));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1454 (.A(\mem[78][5] ),
    .X(net1494));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1455 (.A(\mem[89][12] ),
    .X(net1495));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1456 (.A(\mem[45][10] ),
    .X(net1496));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1457 (.A(\mem[25][6] ),
    .X(net1497));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1458 (.A(\mem[17][5] ),
    .X(net1498));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1459 (.A(\mem[61][2] ),
    .X(net1499));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1460 (.A(\mem[58][3] ),
    .X(net1500));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1461 (.A(\mem[8][11] ),
    .X(net1501));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1462 (.A(\mem[93][5] ),
    .X(net1502));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1463 (.A(\mem[105][3] ),
    .X(net1503));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1464 (.A(\mem[90][0] ),
    .X(net1504));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1465 (.A(\mem[75][10] ),
    .X(net1505));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1466 (.A(\mem[90][3] ),
    .X(net1506));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1467 (.A(\mem[7][6] ),
    .X(net1507));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1468 (.A(\mem[65][15] ),
    .X(net1508));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1469 (.A(\mem[30][0] ),
    .X(net1509));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1470 (.A(\mem[29][4] ),
    .X(net1510));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1471 (.A(\mem[39][0] ),
    .X(net1511));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1472 (.A(\mem[39][12] ),
    .X(net1512));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1473 (.A(\mem[99][12] ),
    .X(net1513));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1474 (.A(\mem[51][6] ),
    .X(net1514));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1475 (.A(\mem[58][13] ),
    .X(net1515));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1476 (.A(\mem[50][2] ),
    .X(net1516));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1477 (.A(\mem[125][12] ),
    .X(net1517));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1478 (.A(\mem[13][8] ),
    .X(net1518));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1479 (.A(\mem[11][11] ),
    .X(net1519));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1480 (.A(\mem[11][14] ),
    .X(net1520));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1481 (.A(\mem[126][1] ),
    .X(net1521));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1482 (.A(\mem[123][9] ),
    .X(net1522));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1483 (.A(\mem[117][7] ),
    .X(net1523));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1484 (.A(\mem[87][14] ),
    .X(net1524));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1485 (.A(\mem[24][2] ),
    .X(net1525));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1486 (.A(\mem[11][8] ),
    .X(net1526));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1487 (.A(\mem[88][9] ),
    .X(net1527));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1488 (.A(\mem[117][5] ),
    .X(net1528));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1489 (.A(\mem[106][13] ),
    .X(net1529));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1490 (.A(\mem[30][4] ),
    .X(net1530));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1491 (.A(\mem[79][15] ),
    .X(net1531));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1492 (.A(\mem[41][5] ),
    .X(net1532));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1493 (.A(\mem[93][8] ),
    .X(net1533));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1494 (.A(\mem[79][10] ),
    .X(net1534));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1495 (.A(\mem[65][13] ),
    .X(net1535));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1496 (.A(\mem[77][3] ),
    .X(net1536));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1497 (.A(\mem[79][2] ),
    .X(net1537));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1498 (.A(\mem[47][2] ),
    .X(net1538));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1499 (.A(\mem[127][11] ),
    .X(net1539));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1500 (.A(\mem[108][0] ),
    .X(net1540));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1501 (.A(\mem[99][7] ),
    .X(net1541));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1502 (.A(\mem[62][2] ),
    .X(net1542));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1503 (.A(\mem[89][9] ),
    .X(net1543));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1504 (.A(\mem[85][11] ),
    .X(net1544));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1505 (.A(\mem[30][3] ),
    .X(net1545));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1506 (.A(\mem[91][13] ),
    .X(net1546));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1507 (.A(\mem[51][12] ),
    .X(net1547));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1508 (.A(\mem[89][4] ),
    .X(net1548));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1509 (.A(\mem[104][6] ),
    .X(net1549));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1510 (.A(\mem[92][0] ),
    .X(net1550));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1511 (.A(\mem[81][5] ),
    .X(net1551));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1512 (.A(\mem[111][13] ),
    .X(net1552));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1513 (.A(\mem[69][2] ),
    .X(net1553));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1514 (.A(\mem[85][9] ),
    .X(net1554));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1515 (.A(\mem[85][14] ),
    .X(net1555));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1516 (.A(\mem[93][3] ),
    .X(net1556));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1517 (.A(\mem[45][13] ),
    .X(net1557));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1518 (.A(\mem[22][14] ),
    .X(net1558));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1519 (.A(\mem[54][1] ),
    .X(net1559));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1520 (.A(\mem[47][11] ),
    .X(net1560));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1521 (.A(\mem[101][0] ),
    .X(net1561));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1522 (.A(\mem[91][4] ),
    .X(net1562));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1523 (.A(\mem[105][4] ),
    .X(net1563));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1524 (.A(\mem[14][12] ),
    .X(net1564));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1525 (.A(\mem[7][2] ),
    .X(net1565));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1526 (.A(\mem[102][9] ),
    .X(net1566));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1527 (.A(\mem[2][14] ),
    .X(net1567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1528 (.A(\mem[101][1] ),
    .X(net1568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1529 (.A(\mem[18][4] ),
    .X(net1569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1530 (.A(\mem[122][6] ),
    .X(net1570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1531 (.A(\mem[29][8] ),
    .X(net1571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1532 (.A(\mem[27][4] ),
    .X(net1572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1533 (.A(\mem[1][12] ),
    .X(net1573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1534 (.A(\mem[102][14] ),
    .X(net1574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1535 (.A(\mem[125][4] ),
    .X(net1575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1536 (.A(\mem[23][10] ),
    .X(net1576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1537 (.A(\mem[66][7] ),
    .X(net1577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1538 (.A(\mem[23][11] ),
    .X(net1578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1539 (.A(\mem[85][15] ),
    .X(net1579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1540 (.A(\mem[80][4] ),
    .X(net1580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1541 (.A(\mem[61][10] ),
    .X(net1581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1542 (.A(\mem[23][15] ),
    .X(net1582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1543 (.A(\mem[124][0] ),
    .X(net1583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1544 (.A(\mem[68][2] ),
    .X(net1584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1545 (.A(\mem[67][3] ),
    .X(net1585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1546 (.A(\mem[60][6] ),
    .X(net1586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1547 (.A(\mem[39][14] ),
    .X(net1587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1548 (.A(\mem[14][0] ),
    .X(net1588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1549 (.A(\mem[99][11] ),
    .X(net1589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1550 (.A(\mem[62][14] ),
    .X(net1590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1551 (.A(\mem[67][0] ),
    .X(net1591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1552 (.A(\mem[115][15] ),
    .X(net1592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1553 (.A(\mem[13][15] ),
    .X(net1593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1554 (.A(\mem[3][4] ),
    .X(net1594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1555 (.A(\mem[99][14] ),
    .X(net1595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1556 (.A(\mem[24][6] ),
    .X(net1596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1557 (.A(\mem[86][13] ),
    .X(net1597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1558 (.A(\mem[26][11] ),
    .X(net1598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1559 (.A(\mem[78][1] ),
    .X(net1599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1560 (.A(\mem[102][6] ),
    .X(net1600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1561 (.A(\mem[1][4] ),
    .X(net1601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1562 (.A(\mem[126][2] ),
    .X(net1602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1563 (.A(\mem[86][12] ),
    .X(net1603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1564 (.A(\mem[86][11] ),
    .X(net1604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1565 (.A(\mem[119][6] ),
    .X(net1605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1566 (.A(\mem[80][7] ),
    .X(net1606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1567 (.A(\mem[79][1] ),
    .X(net1607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1568 (.A(\mem[72][6] ),
    .X(net1608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1569 (.A(\mem[95][4] ),
    .X(net1609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1570 (.A(\mem[47][5] ),
    .X(net1610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1571 (.A(\mem[29][0] ),
    .X(net1611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1572 (.A(\mem[79][9] ),
    .X(net1612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1573 (.A(\mem[42][14] ),
    .X(net1613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1574 (.A(\mem[83][15] ),
    .X(net1614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1575 (.A(\mem[21][0] ),
    .X(net1615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1576 (.A(\mem[14][7] ),
    .X(net1616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1577 (.A(\mem[47][1] ),
    .X(net1617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1578 (.A(\mem[77][14] ),
    .X(net1618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1579 (.A(\mem[77][11] ),
    .X(net1619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1580 (.A(\mem[0][8] ),
    .X(net1620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1581 (.A(\mem[29][13] ),
    .X(net1621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1582 (.A(\mem[78][6] ),
    .X(net1622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1583 (.A(\mem[1][7] ),
    .X(net1623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1584 (.A(\mem[46][11] ),
    .X(net1624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1585 (.A(\mem[26][2] ),
    .X(net1625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1586 (.A(\mem[6][10] ),
    .X(net1626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1587 (.A(\mem[55][1] ),
    .X(net1627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1588 (.A(\mem[19][3] ),
    .X(net1628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1589 (.A(\mem[14][9] ),
    .X(net1629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1590 (.A(\mem[123][10] ),
    .X(net1630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1591 (.A(\mem[102][1] ),
    .X(net1631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1592 (.A(\mem[75][15] ),
    .X(net1632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1593 (.A(\mem[83][3] ),
    .X(net1633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1594 (.A(\mem[27][10] ),
    .X(net1634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1595 (.A(\mem[101][2] ),
    .X(net1635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1596 (.A(\mem[90][8] ),
    .X(net1636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1597 (.A(\mem[14][8] ),
    .X(net1637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1598 (.A(\mem[106][0] ),
    .X(net1638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1599 (.A(\mem[6][4] ),
    .X(net1639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1600 (.A(\mem[7][12] ),
    .X(net1640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1601 (.A(\mem[7][15] ),
    .X(net1641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1602 (.A(\mem[98][13] ),
    .X(net1642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1603 (.A(\mem[115][9] ),
    .X(net1643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1604 (.A(\mem[13][4] ),
    .X(net1644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1605 (.A(\mem[17][4] ),
    .X(net1645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1606 (.A(\mem[56][15] ),
    .X(net1646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1607 (.A(\mem[23][5] ),
    .X(net1647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1608 (.A(\mem[94][6] ),
    .X(net1648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1609 (.A(\mem[17][9] ),
    .X(net1649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1610 (.A(\mem[80][13] ),
    .X(net1650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1611 (.A(\mem[55][14] ),
    .X(net1651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1612 (.A(\mem[63][15] ),
    .X(net1652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1613 (.A(\mem[19][0] ),
    .X(net1653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1614 (.A(\mem[92][11] ),
    .X(net1654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1615 (.A(\mem[24][10] ),
    .X(net1655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1616 (.A(\mem[60][9] ),
    .X(net1656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1617 (.A(\mem[75][0] ),
    .X(net1657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1618 (.A(\mem[30][15] ),
    .X(net1658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1619 (.A(\mem[94][7] ),
    .X(net1659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1620 (.A(\mem[61][12] ),
    .X(net1660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1621 (.A(\mem[27][14] ),
    .X(net1661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1622 (.A(\mem[69][10] ),
    .X(net1662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1623 (.A(\mem[62][15] ),
    .X(net1663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1624 (.A(\mem[122][9] ),
    .X(net1664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1625 (.A(\mem[90][5] ),
    .X(net1665));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1626 (.A(\mem[30][10] ),
    .X(net1666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1627 (.A(\mem[21][6] ),
    .X(net1667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1628 (.A(\mem[31][0] ),
    .X(net1668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1629 (.A(\mem[65][5] ),
    .X(net1669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1630 (.A(\mem[126][12] ),
    .X(net1670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1631 (.A(\mem[59][2] ),
    .X(net1671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1632 (.A(\mem[54][15] ),
    .X(net1672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1633 (.A(\mem[11][15] ),
    .X(net1673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1634 (.A(\mem[94][3] ),
    .X(net1674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1635 (.A(\mem[30][11] ),
    .X(net1675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1636 (.A(\mem[109][12] ),
    .X(net1676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1637 (.A(\mem[123][7] ),
    .X(net1677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1638 (.A(\mem[69][4] ),
    .X(net1678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1639 (.A(\mem[94][1] ),
    .X(net1679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1640 (.A(\mem[111][8] ),
    .X(net1680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1641 (.A(\mem[45][14] ),
    .X(net1681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1642 (.A(\mem[13][7] ),
    .X(net1682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1643 (.A(\mem[95][8] ),
    .X(net1683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1644 (.A(\mem[119][12] ),
    .X(net1684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1645 (.A(\mem[23][14] ),
    .X(net1685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1646 (.A(\mem[77][1] ),
    .X(net1686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1647 (.A(\mem[59][10] ),
    .X(net1687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1648 (.A(\mem[27][12] ),
    .X(net1688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1649 (.A(\mem[27][11] ),
    .X(net1689));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1650 (.A(\mem[93][9] ),
    .X(net1690));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1651 (.A(\mem[81][6] ),
    .X(net1691));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1652 (.A(\mem[70][5] ),
    .X(net1692));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1653 (.A(\mem[23][6] ),
    .X(net1693));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1654 (.A(\mem[102][5] ),
    .X(net1694));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1655 (.A(\mem[91][11] ),
    .X(net1695));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1656 (.A(\mem[95][9] ),
    .X(net1696));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1657 (.A(\mem[23][2] ),
    .X(net1697));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1658 (.A(\mem[110][6] ),
    .X(net1698));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1659 (.A(\mem[56][3] ),
    .X(net1699));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1660 (.A(\mem[31][8] ),
    .X(net1700));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1661 (.A(\mem[111][5] ),
    .X(net1701));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1662 (.A(\mem[9][2] ),
    .X(net1702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1663 (.A(\mem[66][4] ),
    .X(net1703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1664 (.A(\mem[90][13] ),
    .X(net1704));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1665 (.A(\mem[9][10] ),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1666 (.A(\mem[59][7] ),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1667 (.A(\mem[124][9] ),
    .X(net1707));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1668 (.A(\mem[55][15] ),
    .X(net1708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1669 (.A(\mem[53][15] ),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1670 (.A(\mem[22][5] ),
    .X(net1710));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1671 (.A(\mem[31][3] ),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1672 (.A(\mem[27][15] ),
    .X(net1712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1673 (.A(\mem[95][12] ),
    .X(net1713));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1674 (.A(\mem[86][9] ),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1675 (.A(\mem[6][5] ),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1676 (.A(\mem[62][6] ),
    .X(net1716));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1677 (.A(\mem[33][7] ),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1678 (.A(\mem[81][13] ),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1679 (.A(\mem[20][5] ),
    .X(net1719));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1680 (.A(\mem[93][4] ),
    .X(net1720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1681 (.A(\mem[91][7] ),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1682 (.A(\mem[68][0] ),
    .X(net1722));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1683 (.A(\mem[11][5] ),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1684 (.A(\mem[104][14] ),
    .X(net1724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1685 (.A(\mem[121][10] ),
    .X(net1725));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1686 (.A(\mem[67][8] ),
    .X(net1726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1687 (.A(\mem[31][14] ),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1688 (.A(\mem[77][8] ),
    .X(net1728));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1689 (.A(\mem[8][3] ),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1690 (.A(\mem[6][2] ),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1691 (.A(\mem[23][12] ),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1692 (.A(\mem[29][2] ),
    .X(net1732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1693 (.A(\mem[101][5] ),
    .X(net1733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1694 (.A(\mem[95][2] ),
    .X(net1734));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1695 (.A(\mem[17][13] ),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1696 (.A(\mem[75][14] ),
    .X(net1736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1697 (.A(\mem[111][0] ),
    .X(net1737));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1698 (.A(\mem[110][15] ),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1699 (.A(\mem[55][3] ),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1700 (.A(\mem[14][14] ),
    .X(net1740));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1701 (.A(\mem[62][0] ),
    .X(net1741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1702 (.A(\mem[31][10] ),
    .X(net1742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1703 (.A(\mem[77][0] ),
    .X(net1743));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1704 (.A(\mem[25][12] ),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1705 (.A(\mem[91][0] ),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1706 (.A(\mem[62][1] ),
    .X(net1746));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1707 (.A(\mem[22][9] ),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1708 (.A(\mem[55][6] ),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1709 (.A(\mem[89][15] ),
    .X(net1749));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1710 (.A(\mem[89][6] ),
    .X(net1750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1711 (.A(\mem[11][10] ),
    .X(net1751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1712 (.A(\mem[94][4] ),
    .X(net1752));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1713 (.A(\mem[63][6] ),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1714 (.A(\mem[75][4] ),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1715 (.A(\mem[6][0] ),
    .X(net1755));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1716 (.A(\mem[35][12] ),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1717 (.A(\mem[73][8] ),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1718 (.A(\mem[34][12] ),
    .X(net1758));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1719 (.A(\mem[79][13] ),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1720 (.A(\mem[90][15] ),
    .X(net1760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1721 (.A(\mem[63][11] ),
    .X(net1761));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1722 (.A(\mem[25][14] ),
    .X(net1762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1723 (.A(\mem[30][2] ),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1724 (.A(\mem[51][0] ),
    .X(net1764));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1725 (.A(\mem[52][10] ),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1726 (.A(\mem[83][10] ),
    .X(net1766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1727 (.A(\mem[94][10] ),
    .X(net1767));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1728 (.A(\mem[85][2] ),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1729 (.A(\mem[27][8] ),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1730 (.A(\mem[54][4] ),
    .X(net1770));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1731 (.A(\mem[15][8] ),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1732 (.A(\mem[78][13] ),
    .X(net1772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1733 (.A(\mem[26][8] ),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1734 (.A(\mem[121][1] ),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1735 (.A(\mem[31][9] ),
    .X(net1775));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1736 (.A(\mem[14][2] ),
    .X(net1776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1737 (.A(\mem[25][15] ),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1738 (.A(\mem[26][12] ),
    .X(net1778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1739 (.A(\mem[79][0] ),
    .X(net1779));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1740 (.A(\mem[18][8] ),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1741 (.A(\mem[95][3] ),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1742 (.A(\mem[24][11] ),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1743 (.A(\mem[79][14] ),
    .X(net1783));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1744 (.A(\mem[86][7] ),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1745 (.A(\mem[87][0] ),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1746 (.A(\mem[83][13] ),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1747 (.A(\mem[93][14] ),
    .X(net1787));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1748 (.A(\mem[118][14] ),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1749 (.A(\mem[54][9] ),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1750 (.A(\mem[13][13] ),
    .X(net1790));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1751 (.A(\mem[89][5] ),
    .X(net1791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1752 (.A(\mem[55][2] ),
    .X(net1792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1753 (.A(\mem[27][3] ),
    .X(net1793));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1754 (.A(\mem[109][10] ),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1755 (.A(\mem[99][13] ),
    .X(net1795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1756 (.A(\mem[83][4] ),
    .X(net1796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1757 (.A(\mem[89][2] ),
    .X(net1797));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1758 (.A(\mem[47][14] ),
    .X(net1798));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1759 (.A(\mem[90][2] ),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1760 (.A(\mem[95][6] ),
    .X(net1800));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1761 (.A(\mem[85][10] ),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1762 (.A(\mem[66][6] ),
    .X(net1802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1763 (.A(\mem[7][1] ),
    .X(net1803));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1764 (.A(\mem[85][3] ),
    .X(net1804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1765 (.A(\mem[24][14] ),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1766 (.A(\mem[72][3] ),
    .X(net1806));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1767 (.A(\mem[63][4] ),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1768 (.A(\mem[75][11] ),
    .X(net1808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1769 (.A(\mem[43][1] ),
    .X(net1809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1770 (.A(\mem[54][7] ),
    .X(net1810));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1771 (.A(\mem[78][14] ),
    .X(net1811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1772 (.A(\mem[87][13] ),
    .X(net1812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1773 (.A(\mem[46][2] ),
    .X(net1813));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1774 (.A(\mem[94][8] ),
    .X(net1814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1775 (.A(\mem[77][10] ),
    .X(net1815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1776 (.A(\mem[111][2] ),
    .X(net1816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1777 (.A(\mem[83][11] ),
    .X(net1817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1778 (.A(\mem[11][12] ),
    .X(net1818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1779 (.A(\mem[12][0] ),
    .X(net1819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1780 (.A(\mem[75][2] ),
    .X(net1820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1781 (.A(\mem[65][3] ),
    .X(net1821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1782 (.A(\mem[89][3] ),
    .X(net1822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1783 (.A(\mem[27][5] ),
    .X(net1823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1784 (.A(\mem[89][14] ),
    .X(net1824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1785 (.A(\mem[54][8] ),
    .X(net1825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1786 (.A(\mem[19][4] ),
    .X(net1826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1787 (.A(\mem[14][11] ),
    .X(net1827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1788 (.A(\mem[122][4] ),
    .X(net1828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1789 (.A(\mem[78][8] ),
    .X(net1829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1790 (.A(\mem[85][4] ),
    .X(net1830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1791 (.A(\mem[6][6] ),
    .X(net1831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1792 (.A(\mem[30][6] ),
    .X(net1832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1793 (.A(\mem[23][13] ),
    .X(net1833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1794 (.A(\mem[14][3] ),
    .X(net1834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1795 (.A(\mem[91][2] ),
    .X(net1835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1796 (.A(\mem[19][12] ),
    .X(net1836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1797 (.A(\mem[78][9] ),
    .X(net1837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1798 (.A(\mem[7][11] ),
    .X(net1838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1799 (.A(\mem[65][12] ),
    .X(net1839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1800 (.A(\mem[3][8] ),
    .X(net1840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1801 (.A(\mem[119][4] ),
    .X(net1841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1802 (.A(\mem[86][4] ),
    .X(net1842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1803 (.A(\mem[29][10] ),
    .X(net1843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1804 (.A(\mem[2][3] ),
    .X(net1844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1805 (.A(\mem[95][5] ),
    .X(net1845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1806 (.A(\mem[108][11] ),
    .X(net1846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1807 (.A(\mem[25][10] ),
    .X(net1847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1808 (.A(\mem[55][12] ),
    .X(net1848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1809 (.A(\mem[94][11] ),
    .X(net1849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1810 (.A(\mem[21][7] ),
    .X(net1850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1811 (.A(\mem[31][4] ),
    .X(net1851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1812 (.A(\mem[27][1] ),
    .X(net1852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1813 (.A(\mem[109][9] ),
    .X(net1853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1814 (.A(\mem[95][10] ),
    .X(net1854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1815 (.A(\mem[79][8] ),
    .X(net1855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1816 (.A(\mem[19][8] ),
    .X(net1856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1817 (.A(\mem[93][11] ),
    .X(net1857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1818 (.A(\mem[63][13] ),
    .X(net1858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1819 (.A(\mem[75][12] ),
    .X(net1859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1820 (.A(\mem[31][5] ),
    .X(net1860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1821 (.A(\mem[27][0] ),
    .X(net1861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1822 (.A(\mem[90][14] ),
    .X(net1862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1823 (.A(\mem[87][3] ),
    .X(net1863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1824 (.A(\mem[27][7] ),
    .X(net1864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1825 (.A(\mem[118][5] ),
    .X(net1865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1826 (.A(\mem[104][7] ),
    .X(net1866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1827 (.A(\mem[3][7] ),
    .X(net1867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1828 (.A(\mem[38][15] ),
    .X(net1868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1829 (.A(\mem[43][3] ),
    .X(net1869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1830 (.A(\mem[77][4] ),
    .X(net1870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1831 (.A(\mem[13][14] ),
    .X(net1871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1832 (.A(\mem[83][14] ),
    .X(net1872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1833 (.A(\mem[30][1] ),
    .X(net1873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1834 (.A(\mem[69][8] ),
    .X(net1874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1835 (.A(\mem[75][13] ),
    .X(net1875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1836 (.A(\mem[78][10] ),
    .X(net1876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1837 (.A(\mem[94][13] ),
    .X(net1877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1838 (.A(\mem[65][11] ),
    .X(net1878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1839 (.A(\mem[121][12] ),
    .X(net1879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1840 (.A(\mem[13][10] ),
    .X(net1880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1841 (.A(\mem[94][2] ),
    .X(net1881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1842 (.A(\mem[91][14] ),
    .X(net1882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1843 (.A(\mem[54][13] ),
    .X(net1883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1844 (.A(\mem[58][5] ),
    .X(net1884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1845 (.A(\mem[93][0] ),
    .X(net1885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1846 (.A(\mem[7][7] ),
    .X(net1886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1847 (.A(\mem[70][9] ),
    .X(net1887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1848 (.A(\mem[30][12] ),
    .X(net1888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1849 (.A(\mem[85][13] ),
    .X(net1889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1850 (.A(\mem[31][13] ),
    .X(net1890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1851 (.A(\mem[89][1] ),
    .X(net1891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1852 (.A(\mem[94][15] ),
    .X(net1892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1853 (.A(\mem[31][15] ),
    .X(net1893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1854 (.A(\mem[3][5] ),
    .X(net1894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1855 (.A(\mem[87][15] ),
    .X(net1895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1856 (.A(\mem[83][7] ),
    .X(net1896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1857 (.A(\mem[71][15] ),
    .X(net1897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1858 (.A(\mem[39][7] ),
    .X(net1898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1859 (.A(\mem[44][8] ),
    .X(net1899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1860 (.A(\mem[58][2] ),
    .X(net1900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1861 (.A(\mem[86][3] ),
    .X(net1901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1862 (.A(\mem[39][8] ),
    .X(net1902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1863 (.A(\mem[75][3] ),
    .X(net1903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1864 (.A(\mem[7][9] ),
    .X(net1904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1865 (.A(\mem[30][13] ),
    .X(net1905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1866 (.A(\mem[97][5] ),
    .X(net1906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1867 (.A(\mem[55][11] ),
    .X(net1907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1868 (.A(\mem[80][2] ),
    .X(net1908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1869 (.A(\mem[93][12] ),
    .X(net1909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1870 (.A(\mem[43][10] ),
    .X(net1910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1871 (.A(\mem[94][12] ),
    .X(net1911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1872 (.A(\mem[106][4] ),
    .X(net1912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1873 (.A(\mem[6][3] ),
    .X(net1913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1874 (.A(\mem[79][3] ),
    .X(net1914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1875 (.A(\mem[91][9] ),
    .X(net1915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1876 (.A(\mem[28][6] ),
    .X(net1916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1877 (.A(\mem[3][6] ),
    .X(net1917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1878 (.A(\mem[72][2] ),
    .X(net1918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1879 (.A(\mem[49][15] ),
    .X(net1919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1880 (.A(\mem[71][4] ),
    .X(net1920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1881 (.A(\mem[104][8] ),
    .X(net1921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1882 (.A(\mem[78][4] ),
    .X(net1922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1883 (.A(\mem[51][8] ),
    .X(net1923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1884 (.A(\mem[72][0] ),
    .X(net1924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1885 (.A(\mem[86][15] ),
    .X(net1925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1886 (.A(\mem[23][9] ),
    .X(net1926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1887 (.A(\mem[30][7] ),
    .X(net1927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1888 (.A(\mem[7][10] ),
    .X(net1928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1889 (.A(\mem[86][2] ),
    .X(net1929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1890 (.A(\mem[73][1] ),
    .X(net1930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1891 (.A(\mem[47][13] ),
    .X(net1931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1892 (.A(\mem[58][4] ),
    .X(net1932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1893 (.A(\mem[67][4] ),
    .X(net1933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1894 (.A(\mem[30][8] ),
    .X(net1934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1895 (.A(\mem[87][10] ),
    .X(net1935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1896 (.A(\mem[104][13] ),
    .X(net1936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1897 (.A(\mem[69][7] ),
    .X(net1937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1898 (.A(\mem[120][15] ),
    .X(net1938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1899 (.A(\mem[91][5] ),
    .X(net1939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1900 (.A(\mem[19][2] ),
    .X(net1940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1901 (.A(\mem[75][9] ),
    .X(net1941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1902 (.A(\mem[111][6] ),
    .X(net1942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1903 (.A(\mem[83][2] ),
    .X(net1943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1904 (.A(\mem[69][9] ),
    .X(net1944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1905 (.A(\mem[62][13] ),
    .X(net1945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1906 (.A(\mem[23][3] ),
    .X(net1946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1907 (.A(\mem[58][8] ),
    .X(net1947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1908 (.A(\mem[14][15] ),
    .X(net1948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1909 (.A(\mem[11][6] ),
    .X(net1949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1910 (.A(\mem[94][9] ),
    .X(net1950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1911 (.A(\mem[14][4] ),
    .X(net1951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1912 (.A(\mem[80][1] ),
    .X(net1952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1913 (.A(\mem[71][1] ),
    .X(net1953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1914 (.A(\mem[90][1] ),
    .X(net1954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1915 (.A(\mem[108][10] ),
    .X(net1955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1916 (.A(\mem[91][10] ),
    .X(net1956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1917 (.A(\mem[24][12] ),
    .X(net1957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1918 (.A(\mem[23][0] ),
    .X(net1958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1919 (.A(\mem[83][0] ),
    .X(net1959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1920 (.A(\mem[13][11] ),
    .X(net1960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1921 (.A(\mem[80][8] ),
    .X(net1961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1922 (.A(\mem[40][15] ),
    .X(net1962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1923 (.A(\mem[86][14] ),
    .X(net1963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1924 (.A(\mem[101][6] ),
    .X(net1964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1925 (.A(\mem[78][7] ),
    .X(net1965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1926 (.A(\mem[91][12] ),
    .X(net1966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1927 (.A(\mem[11][13] ),
    .X(net1967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1928 (.A(\mem[8][13] ),
    .X(net1968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1929 (.A(\mem[83][9] ),
    .X(net1969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1930 (.A(\mem[51][14] ),
    .X(net1970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1931 (.A(\mem[71][9] ),
    .X(net1971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1932 (.A(\mem[71][5] ),
    .X(net1972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1933 (.A(\mem[87][2] ),
    .X(net1973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1934 (.A(\mem[85][5] ),
    .X(net1974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1935 (.A(\mem[79][11] ),
    .X(net1975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1936 (.A(\mem[88][1] ),
    .X(net1976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1937 (.A(\mem[77][7] ),
    .X(net1977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1938 (.A(\mem[126][0] ),
    .X(net1978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1939 (.A(\mem[71][0] ),
    .X(net1979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1940 (.A(\mem[91][8] ),
    .X(net1980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1941 (.A(\mem[83][5] ),
    .X(net1981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1942 (.A(\mem[90][6] ),
    .X(net1982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1943 (.A(\mem[71][2] ),
    .X(net1983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1944 (.A(\mem[110][0] ),
    .X(net1984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1945 (.A(\mem[66][2] ),
    .X(net1985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1946 (.A(\mem[94][0] ),
    .X(net1986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1947 (.A(\mem[67][7] ),
    .X(net1987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1948 (.A(\mem[85][1] ),
    .X(net1988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1949 (.A(\mem[7][0] ),
    .X(net1989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1950 (.A(\mem[29][14] ),
    .X(net1990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1951 (.A(\mem[3][1] ),
    .X(net1991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1952 (.A(\mem[86][8] ),
    .X(net1992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1953 (.A(\mem[75][6] ),
    .X(net1993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1954 (.A(\mem[30][5] ),
    .X(net1994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1955 (.A(\mem[79][12] ),
    .X(net1995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1956 (.A(\mem[91][1] ),
    .X(net1996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1957 (.A(\mem[95][1] ),
    .X(net1997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1958 (.A(\mem[69][0] ),
    .X(net1998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1959 (.A(\mem[115][4] ),
    .X(net1999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1960 (.A(\mem[39][10] ),
    .X(net2000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1961 (.A(\mem[15][0] ),
    .X(net2001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1962 (.A(\mem[29][7] ),
    .X(net2002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1963 (.A(\mem[71][14] ),
    .X(net2003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1964 (.A(\mem[78][2] ),
    .X(net2004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1965 (.A(\mem[23][8] ),
    .X(net2005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1966 (.A(\mem[93][1] ),
    .X(net2006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1967 (.A(\mem[87][8] ),
    .X(net2007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1968 (.A(\mem[87][9] ),
    .X(net2008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1969 (.A(\mem[117][14] ),
    .X(net2009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1970 (.A(\mem[83][8] ),
    .X(net2010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1971 (.A(\mem[17][14] ),
    .X(net2011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1972 (.A(\mem[11][3] ),
    .X(net2012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1973 (.A(\mem[108][6] ),
    .X(net2013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1974 (.A(\mem[95][15] ),
    .X(net2014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1975 (.A(\mem[3][13] ),
    .X(net2015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1976 (.A(\mem[83][6] ),
    .X(net2016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1977 (.A(\mem[83][12] ),
    .X(net2017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1978 (.A(\mem[71][12] ),
    .X(net2018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1979 (.A(\mem[75][1] ),
    .X(net2019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1980 (.A(\mem[3][9] ),
    .X(net2020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1981 (.A(\mem[11][0] ),
    .X(net2021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1982 (.A(\mem[18][6] ),
    .X(net2022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1983 (.A(\mem[87][1] ),
    .X(net2023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1984 (.A(\mem[11][7] ),
    .X(net2024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1985 (.A(\mem[7][8] ),
    .X(net2025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1986 (.A(\mem[71][10] ),
    .X(net2026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1987 (.A(\mem[11][4] ),
    .X(net2027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1988 (.A(\mem[3][3] ),
    .X(net2028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1989 (.A(\mem[71][8] ),
    .X(net2029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1990 (.A(\mem[29][11] ),
    .X(net2030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1991 (.A(\mem[104][0] ),
    .X(net2031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1992 (.A(\mem[10][0] ),
    .X(net2032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1993 (.A(\mem[78][0] ),
    .X(net2033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1994 (.A(\mem[9][0] ),
    .X(net2034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1995 (.A(\mem[49][13] ),
    .X(net2035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1996 (.A(\mem[78][3] ),
    .X(net2036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1997 (.A(\mem[93][10] ),
    .X(net2037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1998 (.A(\mem[71][7] ),
    .X(net2038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1999 (.A(\mem[80][11] ),
    .X(net2039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2000 (.A(\mem[69][3] ),
    .X(net2040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2001 (.A(\mem[104][15] ),
    .X(net2041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2002 (.A(\mem[75][5] ),
    .X(net2042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2003 (.A(\mem[29][15] ),
    .X(net2043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2004 (.A(\mem[104][2] ),
    .X(net2044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2005 (.A(\mem[86][1] ),
    .X(net2045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2006 (.A(\mem[71][3] ),
    .X(net2046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2007 (.A(\mem[51][5] ),
    .X(net2047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2008 (.A(\mem[39][2] ),
    .X(net2048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2009 (.A(\mem[7][5] ),
    .X(net2049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2010 (.A(\mem[87][5] ),
    .X(net2050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2011 (.A(\mem[88][5] ),
    .X(net2051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2012 (.A(\mem[91][6] ),
    .X(net2052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2013 (.A(\mem[83][1] ),
    .X(net2053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2014 (.A(\mem[49][12] ),
    .X(net2054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2015 (.A(\mem[67][2] ),
    .X(net2055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2016 (.A(\mem[11][2] ),
    .X(net2056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2017 (.A(\mem[80][6] ),
    .X(net2057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2018 (.A(\mem[71][11] ),
    .X(net2058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2019 (.A(\mem[29][12] ),
    .X(net2059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2020 (.A(\mem[49][14] ),
    .X(net2060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2021 (.A(\mem[86][5] ),
    .X(net2061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2022 (.A(\mem[3][11] ),
    .X(net2062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2023 (.A(\mem[49][9] ),
    .X(net2063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2024 (.A(\mem[49][1] ),
    .X(net2064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2025 (.A(\mem[8][15] ),
    .X(net2065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2026 (.A(\mem[3][2] ),
    .X(net2066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2027 (.A(\mem[80][10] ),
    .X(net2067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2028 (.A(\mem[80][14] ),
    .X(net2068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2029 (.A(\mem[3][0] ),
    .X(net2069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2030 (.A(\mem[49][5] ),
    .X(net2070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2031 (.A(\mem[87][6] ),
    .X(net2071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2032 (.A(\mem[69][1] ),
    .X(net2072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2033 (.A(\mem[5][0] ),
    .X(net2073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2034 (.A(\mem[3][10] ),
    .X(net2074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2035 (.A(\mem[80][12] ),
    .X(net2075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2036 (.A(\mem[71][13] ),
    .X(net2076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2037 (.A(\mem[49][6] ),
    .X(net2077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2038 (.A(\mem[86][6] ),
    .X(net2078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2039 (.A(\mem[3][15] ),
    .X(net2079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2040 (.A(\mem[3][12] ),
    .X(net2080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2041 (.A(\mem[49][8] ),
    .X(net2081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2042 (.A(\mem[49][0] ),
    .X(net2082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2043 (.A(\mem[85][6] ),
    .X(net2083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2044 (.A(\mem[49][2] ),
    .X(net2084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2045 (.A(\mem[49][3] ),
    .X(net2085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2046 (.A(\mem[49][7] ),
    .X(net2086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2047 (.A(\mem[3][14] ),
    .X(net2087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2048 (.A(\mem[49][4] ),
    .X(net2088));
 sky130_fd_sc_hd__diode_2 ANTENNA__12325__S (.DIODE(_02076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12323__S (.DIODE(_02076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12321__S (.DIODE(_02076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12319__S (.DIODE(_02076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12317__S (.DIODE(_02076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12315__S (.DIODE(_02076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12294__A (.DIODE(_02076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12313__S (.DIODE(_02077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12311__S (.DIODE(_02077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__S (.DIODE(_02077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12307__S (.DIODE(_02077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12305__S (.DIODE(_02077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12303__S (.DIODE(_02077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12301__S (.DIODE(_02077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__S (.DIODE(_02077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12297__S (.DIODE(_02077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12295__S (.DIODE(_02077_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12359__S (.DIODE(_02094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12357__S (.DIODE(_02094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12355__S (.DIODE(_02094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12353__S (.DIODE(_02094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12351__S (.DIODE(_02094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12349__S (.DIODE(_02094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12328__A (.DIODE(_02094_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12347__S (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12345__S (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12343__S (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__S (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12339__S (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12337__S (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12335__S (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12333__S (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12331__S (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12329__S (.DIODE(_02095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12394__S (.DIODE(_02113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12392__S (.DIODE(_02113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12390__S (.DIODE(_02113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12388__S (.DIODE(_02113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12386__S (.DIODE(_02113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12384__S (.DIODE(_02113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12363__A (.DIODE(_02113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12382__S (.DIODE(_02114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12380__S (.DIODE(_02114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12378__S (.DIODE(_02114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12376__S (.DIODE(_02114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12374__S (.DIODE(_02114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12372__S (.DIODE(_02114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12370__S (.DIODE(_02114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12368__S (.DIODE(_02114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12366__S (.DIODE(_02114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12364__S (.DIODE(_02114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12428__S (.DIODE(_02131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12426__S (.DIODE(_02131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12424__S (.DIODE(_02131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12422__S (.DIODE(_02131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__S (.DIODE(_02131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12418__S (.DIODE(_02131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12397__A (.DIODE(_02131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12416__S (.DIODE(_02132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12414__S (.DIODE(_02132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12412__S (.DIODE(_02132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12410__S (.DIODE(_02132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12408__S (.DIODE(_02132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12406__S (.DIODE(_02132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12404__S (.DIODE(_02132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12402__S (.DIODE(_02132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12400__S (.DIODE(_02132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12398__S (.DIODE(_02132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12463__S (.DIODE(_02150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12461__S (.DIODE(_02150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12459__S (.DIODE(_02150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12457__S (.DIODE(_02150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12455__S (.DIODE(_02150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12453__S (.DIODE(_02150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12432__A (.DIODE(_02150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12451__S (.DIODE(_02151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12449__S (.DIODE(_02151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12447__S (.DIODE(_02151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12445__S (.DIODE(_02151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12443__S (.DIODE(_02151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12441__S (.DIODE(_02151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__S (.DIODE(_02151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12437__S (.DIODE(_02151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12435__S (.DIODE(_02151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12433__S (.DIODE(_02151_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12498__S (.DIODE(_02169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12496__S (.DIODE(_02169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12494__S (.DIODE(_02169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12492__S (.DIODE(_02169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12490__S (.DIODE(_02169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12488__S (.DIODE(_02169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12467__A (.DIODE(_02169_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12486__S (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12484__S (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12482__S (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12480__S (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12478__S (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12476__S (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12474__S (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12472__S (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12470__S (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12468__S (.DIODE(_02170_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12533__S (.DIODE(_02188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12531__S (.DIODE(_02188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12529__S (.DIODE(_02188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12527__S (.DIODE(_02188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12525__S (.DIODE(_02188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12523__S (.DIODE(_02188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12502__A (.DIODE(_02188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12521__S (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12519__S (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12517__S (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12515__S (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__S (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12511__S (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12509__S (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12507__S (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12505__S (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12503__S (.DIODE(_02189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12567__S (.DIODE(_02206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12565__S (.DIODE(_02206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12563__S (.DIODE(_02206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12561__S (.DIODE(_02206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12559__S (.DIODE(_02206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12557__S (.DIODE(_02206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12536__A (.DIODE(_02206_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12555__S (.DIODE(_02207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12553__S (.DIODE(_02207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12551__S (.DIODE(_02207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12549__S (.DIODE(_02207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12547__S (.DIODE(_02207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12545__S (.DIODE(_02207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12543__S (.DIODE(_02207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12541__S (.DIODE(_02207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12539__S (.DIODE(_02207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12537__S (.DIODE(_02207_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__S (.DIODE(_02225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12600__S (.DIODE(_02225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12598__S (.DIODE(_02225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12596__S (.DIODE(_02225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12594__S (.DIODE(_02225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12592__S (.DIODE(_02225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12571__A (.DIODE(_02225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12590__S (.DIODE(_02226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12588__S (.DIODE(_02226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12586__S (.DIODE(_02226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12584__S (.DIODE(_02226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12582__S (.DIODE(_02226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12580__S (.DIODE(_02226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12578__S (.DIODE(_02226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12576__S (.DIODE(_02226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12574__S (.DIODE(_02226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12572__S (.DIODE(_02226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12637__S (.DIODE(_02244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12635__S (.DIODE(_02244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12633__S (.DIODE(_02244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12631__S (.DIODE(_02244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12629__S (.DIODE(_02244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12627__S (.DIODE(_02244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12606__A (.DIODE(_02244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12625__S (.DIODE(_02245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12623__S (.DIODE(_02245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12621__S (.DIODE(_02245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12619__S (.DIODE(_02245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12617__S (.DIODE(_02245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12615__S (.DIODE(_02245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12613__S (.DIODE(_02245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12611__S (.DIODE(_02245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__S (.DIODE(_02245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12607__S (.DIODE(_02245_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12672__S (.DIODE(_02263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12670__S (.DIODE(_02263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__S (.DIODE(_02263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12666__S (.DIODE(_02263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12664__S (.DIODE(_02263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12662__S (.DIODE(_02263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12641__A (.DIODE(_02263_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12660__S (.DIODE(_02264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12658__S (.DIODE(_02264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12656__S (.DIODE(_02264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12654__S (.DIODE(_02264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12652__S (.DIODE(_02264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12650__S (.DIODE(_02264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12648__S (.DIODE(_02264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12646__S (.DIODE(_02264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12644__S (.DIODE(_02264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12642__S (.DIODE(_02264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12707__S (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12705__S (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12703__S (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12701__S (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12699__S (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12697__S (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12676__A (.DIODE(_02282_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12695__S (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12693__S (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12691__S (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12689__S (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12687__S (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12685__S (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12683__S (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12681__S (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12679__S (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12677__S (.DIODE(_02283_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12742__S (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12740__S (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12738__S (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12736__S (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12734__S (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12732__S (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12711__A (.DIODE(_02301_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12730__S (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12728__S (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12726__S (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12724__S (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12722__S (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__S (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12718__S (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12716__S (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12714__S (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12712__S (.DIODE(_02302_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12776__S (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12774__S (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12772__S (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12770__S (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12768__S (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12766__S (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12745__A (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12764__S (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12762__S (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12760__S (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12758__S (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12756__S (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12754__S (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12752__S (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12750__S (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12748__S (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12746__S (.DIODE(_02320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12810__S (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12808__S (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12806__S (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12804__S (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12802__S (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12800__S (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12779__A (.DIODE(_02337_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12798__S (.DIODE(_02338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12796__S (.DIODE(_02338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12794__S (.DIODE(_02338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12792__S (.DIODE(_02338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12790__S (.DIODE(_02338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12788__S (.DIODE(_02338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12786__S (.DIODE(_02338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12784__S (.DIODE(_02338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12782__S (.DIODE(_02338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12780__S (.DIODE(_02338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08480__B (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08409__B (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08133__A1 (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08042__A1 (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07864__A1 (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__A1 (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07593__A1 (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07503__A1 (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06564__A (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06407__A (.DIODE(_02355_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07774__A1 (.DIODE(_02356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07549__A1 (.DIODE(_02356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07459__A1 (.DIODE(_02356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07369__A1 (.DIODE(_02356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07323__A1 (.DIODE(_02356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07276__A1 (.DIODE(_02356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07096__A1 (.DIODE(_02356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06998__A1 (.DIODE(_02356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06896__A1 (.DIODE(_02356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06563__A1 (.DIODE(_02356_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__A (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08212__A (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08102__A (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07772__B1 (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07321__B1 (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07048__A (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06662__A (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06565__A (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06533__A (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06409__A (.DIODE(_02357_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08132__A1 (.DIODE(_02358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08041__A1 (.DIODE(_02358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__A1 (.DIODE(_02358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07743__A (.DIODE(_02358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07682__A1 (.DIODE(_02358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07592__A1 (.DIODE(_02358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07292__A (.DIODE(_02358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__A (.DIODE(_02358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06850__A (.DIODE(_02358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06470__A (.DIODE(_02358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06836__A (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06581__A (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06572__A (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06510__A (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06480__A (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06429__B (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06426__A (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06422__B (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06419__B (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06412__A_N (.DIODE(_02359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06655__A (.DIODE(_02360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06571__A (.DIODE(_02360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06552__A (.DIODE(_02360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06508__A (.DIODE(_02360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06483__A (.DIODE(_02360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06461__A (.DIODE(_02360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06429__A (.DIODE(_02360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06424__A (.DIODE(_02360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06422__A (.DIODE(_02360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06412__B (.DIODE(_02360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07097__A (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06953__A (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06843__A (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06788__A (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06623__A (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06589__A (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06566__A (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06450__A (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06436__A (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06414__A (.DIODE(_02362_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__A2 (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08007__A2 (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07829__A2 (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07648__A2 (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07326__A2 (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07233__A2 (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07049__A2 (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06949__A2 (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06831__A2 (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06418__A2 (.DIODE(_02363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08089__B1 (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__B1 (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07821__B1 (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07640__B1 (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07550__B1 (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06567__A (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06473__A (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06417__A (.DIODE(_02365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07730__B1 (.DIODE(_02366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07596__B1 (.DIODE(_02366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07506__B1 (.DIODE(_02366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07416__B1 (.DIODE(_02366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07326__B1 (.DIODE(_02366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07233__B1 (.DIODE(_02366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07049__B1 (.DIODE(_02366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06949__B1 (.DIODE(_02366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06831__B1 (.DIODE(_02366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06418__B1 (.DIODE(_02366_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__A2 (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07010__A (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06853__A (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06632__A (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06605__A (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06594__A (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06496__A (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06458__A (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06444__A (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06421__A (.DIODE(_02369_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08104__A2 (.DIODE(_02370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08014__A2 (.DIODE(_02370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07836__A2 (.DIODE(_02370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07732__A2 (.DIODE(_02370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07655__A2 (.DIODE(_02370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__A2 (.DIODE(_02370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06951__A2 (.DIODE(_02370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06834__A2 (.DIODE(_02370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06477__A2 (.DIODE(_02370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06428__A2 (.DIODE(_02370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07688__B1 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07598__B1 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07508__B1 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07418__B1 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07328__B1 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__B1 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07052__B1 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06951__B1 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06834__B1 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06428__B1 (.DIODE(_02372_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06868__A (.DIODE(_02373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06855__A (.DIODE(_02373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06722__A (.DIODE(_02373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06625__A (.DIODE(_02373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06607__A (.DIODE(_02373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06580__A (.DIODE(_02373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06537__A (.DIODE(_02373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06517__A (.DIODE(_02373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06438__A (.DIODE(_02373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06425__A (.DIODE(_02373_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__S0 (.DIODE(_02374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07309__S0 (.DIODE(_02374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07234__A (.DIODE(_02374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07051__A (.DIODE(_02374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06982__A (.DIODE(_02374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06950__A (.DIODE(_02374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06833__A (.DIODE(_02374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06644__A (.DIODE(_02374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06476__A (.DIODE(_02374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06427__A (.DIODE(_02374_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08093__C_N (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08003__C_N (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07825__C_N (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06890__A (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06725__A (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06677__A (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06554__A (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06550__A (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06476__B (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06427__B (.DIODE(_02375_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06971__A (.DIODE(_02378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06865__A (.DIODE(_02378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06621__A (.DIODE(_02378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06430__A (.DIODE(_02378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08109__B (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08019__B (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06841__A (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06701__A (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06613__A (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06586__A (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06575__A (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06489__A (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06446__A (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06431__A (.DIODE(_02379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08096__A2 (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08006__A2 (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__A2 (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07419__A2 (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07329__A2 (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07236__A2 (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__A2 (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06952__A2 (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06835__A2 (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06435__A2 (.DIODE(_02380_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06654__A (.DIODE(_02381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06556__A_N (.DIODE(_02381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06548__B (.DIODE(_02381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06545__A (.DIODE(_02381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06534__A (.DIODE(_02381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06525__A (.DIODE(_02381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06522__A (.DIODE(_02381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06466__B (.DIODE(_02381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06447__A (.DIODE(_02381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06433__A (.DIODE(_02381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08106__B1 (.DIODE(_02383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__B1 (.DIODE(_02383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07419__B1 (.DIODE(_02383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07329__B1 (.DIODE(_02383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07236__B1 (.DIODE(_02383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__B1 (.DIODE(_02383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06952__B1 (.DIODE(_02383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06835__B1 (.DIODE(_02383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06482__B1 (.DIODE(_02383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06435__B1 (.DIODE(_02383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08111__A2 (.DIODE(_02385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08021__A2 (.DIODE(_02385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07843__A2 (.DIODE(_02385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07662__A2 (.DIODE(_02385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07572__A2 (.DIODE(_02385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07482__A2 (.DIODE(_02385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06838__A2 (.DIODE(_02385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06486__A2 (.DIODE(_02385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06474__B (.DIODE(_02385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06442__A2 (.DIODE(_02385_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08104__B1 (.DIODE(_02386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07732__B1 (.DIODE(_02386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__B1 (.DIODE(_02386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07238__B1 (.DIODE(_02386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07055__B1 (.DIODE(_02386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06955__B1 (.DIODE(_02386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06838__B1 (.DIODE(_02386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06696__A (.DIODE(_02386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06486__B1 (.DIODE(_02386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06442__B1 (.DIODE(_02386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08103__A (.DIODE(_02387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07731__A (.DIODE(_02387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07420__A (.DIODE(_02387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07330__A (.DIODE(_02387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07278__A (.DIODE(_02387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07237__A (.DIODE(_02387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07054__A (.DIODE(_02387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06954__A (.DIODE(_02387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06837__A (.DIODE(_02387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06441__A (.DIODE(_02387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07281__A (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06921__A (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06869__A (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06856__A (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06832__A (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06626__A (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06597__A (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06484__A (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06463__A (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06440__A (.DIODE(_02388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08103__B (.DIODE(_02389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08013__B (.DIODE(_02389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07835__B (.DIODE(_02389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07731__B (.DIODE(_02389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07654__B (.DIODE(_02389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07564__B (.DIODE(_02389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07474__B (.DIODE(_02389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07384__B (.DIODE(_02389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07278__B (.DIODE(_02389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06441__C_N (.DIODE(_02389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07755__A2 (.DIODE(_02393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07741__A2 (.DIODE(_02393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07304__A2 (.DIODE(_02393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07290__A2 (.DIODE(_02393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06840__A (.DIODE(_02393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06695__A (.DIODE(_02393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06612__A (.DIODE(_02393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06585__A (.DIODE(_02393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06488__A (.DIODE(_02393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06445__A (.DIODE(_02393_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08108__A2 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08018__A2 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07840__A2 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07659__A2 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07569__A2 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__A2 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07389__A2 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07117__A2 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07020__A2 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06454__A2 (.DIODE(_02394_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08106__A2 (.DIODE(_02395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__A2 (.DIODE(_02395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07838__A2 (.DIODE(_02395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07657__A2 (.DIODE(_02395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07567__A2 (.DIODE(_02395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07477__A2 (.DIODE(_02395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07387__A2 (.DIODE(_02395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07115__A2 (.DIODE(_02395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07018__A2 (.DIODE(_02395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06449__A2 (.DIODE(_02395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08096__B1 (.DIODE(_02396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08006__B1 (.DIODE(_02396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07828__B1 (.DIODE(_02396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07647__B1 (.DIODE(_02396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06587__A (.DIODE(_02396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06490__A (.DIODE(_02396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06448__A (.DIODE(_02396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07693__B1 (.DIODE(_02397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__B1 (.DIODE(_02397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__B1 (.DIODE(_02397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07423__B1 (.DIODE(_02397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__B1 (.DIODE(_02397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07240__B1 (.DIODE(_02397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07057__B1 (.DIODE(_02397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06957__B1 (.DIODE(_02397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06842__B1 (.DIODE(_02397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06449__B1 (.DIODE(_02397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__A2 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08017__A2 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__A2 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07658__A2 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__A2 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07478__A2 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07388__A2 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07116__A2 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06852__A (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06453__A2 (.DIODE(_02399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08371__B (.DIODE(_02400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__B1 (.DIODE(_02400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08001__B1 (.DIODE(_02400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__B1 (.DIODE(_02400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07642__B1 (.DIODE(_02400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06968__A (.DIODE(_02400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06617__A (.DIODE(_02400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06590__A (.DIODE(_02400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06493__A (.DIODE(_02400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06452__A (.DIODE(_02400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__B1 (.DIODE(_02401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08017__B1 (.DIODE(_02401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07514__B1 (.DIODE(_02401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07424__B1 (.DIODE(_02401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07334__B1 (.DIODE(_02401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07241__B1 (.DIODE(_02401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07058__B1 (.DIODE(_02401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06958__B1 (.DIODE(_02401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06844__B1 (.DIODE(_02401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06453__B1 (.DIODE(_02401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08298__B (.DIODE(_02404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08209__B (.DIODE(_02404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08094__A2 (.DIODE(_02404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__A2 (.DIODE(_02404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06872__A (.DIODE(_02404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06691__A (.DIODE(_02404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06629__A (.DIODE(_02404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06616__A (.DIODE(_02404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06492__A (.DIODE(_02404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06456__A (.DIODE(_02404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__A2 (.DIODE(_02405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08022__A2 (.DIODE(_02405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07844__A2 (.DIODE(_02405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07738__A2 (.DIODE(_02405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07663__A2 (.DIODE(_02405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07573__A2 (.DIODE(_02405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07297__A2 (.DIODE(_02405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__A2 (.DIODE(_02405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06593__A (.DIODE(_02405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06457__A (.DIODE(_02405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07915__A2 (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07245__A2 (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07193__A2 (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07062__A2 (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06962__A2 (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06849__A2 (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06783__A2 (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06721__A (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06502__A2 (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06469__A2 (.DIODE(_02406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08114__A2 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08024__A2 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07846__A2 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07665__A2 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07575__A2 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__A2 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07061__A2 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__A2 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06848__A2 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06465__A2 (.DIODE(_02407_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__A (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07064__A (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06867__A (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06854__A (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06716__A (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06633__A (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06624__A (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06595__A (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06497__A (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06460__A (.DIODE(_02408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08114__B1 (.DIODE(_02409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08024__B1 (.DIODE(_02409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07846__B1 (.DIODE(_02409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07665__B1 (.DIODE(_02409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07337__B1 (.DIODE(_02409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__B1 (.DIODE(_02409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07061__B1 (.DIODE(_02409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__B1 (.DIODE(_02409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06848__B1 (.DIODE(_02409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06465__B1 (.DIODE(_02409_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07039__A (.DIODE(_02410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06940__A (.DIODE(_02410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06846__A (.DIODE(_02410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06676__A (.DIODE(_02410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06673__A (.DIODE(_02410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06634__A (.DIODE(_02410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06596__A (.DIODE(_02410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06498__A (.DIODE(_02410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06478__A (.DIODE(_02410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06462__A (.DIODE(_02410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__A (.DIODE(_02411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08023__A (.DIODE(_02411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07845__A (.DIODE(_02411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__S0 (.DIODE(_02411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07664__A (.DIODE(_02411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07574__A (.DIODE(_02411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07484__A (.DIODE(_02411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07312__S0 (.DIODE(_02411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06778__A (.DIODE(_02411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06464__A (.DIODE(_02411_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07696__B (.DIODE(_02412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07606__B (.DIODE(_02412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07516__B (.DIODE(_02412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07426__B (.DIODE(_02412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07336__B (.DIODE(_02412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07243__B (.DIODE(_02412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07060__B (.DIODE(_02412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06960__B (.DIODE(_02412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06847__B (.DIODE(_02412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06464__B (.DIODE(_02412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07753__B1 (.DIODE(_02416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07302__B1 (.DIODE(_02416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__B1 (.DIODE(_02416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07075__B1 (.DIODE(_02416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06975__B1 (.DIODE(_02416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06878__A (.DIODE(_02416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06873__B1 (.DIODE(_02416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06600__A (.DIODE(_02416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06501__A (.DIODE(_02416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06468__A (.DIODE(_02416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__B1 (.DIODE(_02417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07428__C1 (.DIODE(_02417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07338__C1 (.DIODE(_02417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07245__C1 (.DIODE(_02417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07198__B1 (.DIODE(_02417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07062__C1 (.DIODE(_02417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06962__C1 (.DIODE(_02417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06849__C1 (.DIODE(_02417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06729__A (.DIODE(_02417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06469__C1 (.DIODE(_02417_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06563__A2 (.DIODE(_02419_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08409__A (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08300__A (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__A (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08026__A (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07848__A (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06851__A (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06640__A (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06603__A (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06504__A (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06472__A (.DIODE(_02420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__A (.DIODE(_02421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08034__A (.DIODE(_02421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07856__A (.DIODE(_02421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__A (.DIODE(_02421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__A (.DIODE(_02421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07585__A (.DIODE(_02421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07495__A (.DIODE(_02421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07405__A (.DIODE(_02421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__A (.DIODE(_02421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06503__A (.DIODE(_02421_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08698__C (.DIODE(_02422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08105__C1 (.DIODE(_02422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08015__C1 (.DIODE(_02422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07837__C1 (.DIODE(_02422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07656__C1 (.DIODE(_02422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07277__B1 (.DIODE(_02422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06859__A (.DIODE(_02422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06693__A (.DIODE(_02422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06610__A (.DIODE(_02422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06487__A1 (.DIODE(_02422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08094__B1 (.DIODE(_02424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__B1 (.DIODE(_02424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__B1 (.DIODE(_02424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07645__B1 (.DIODE(_02424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07555__B1 (.DIODE(_02424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07465__B1 (.DIODE(_02424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07375__B1 (.DIODE(_02424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07103__B1 (.DIODE(_02424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07004__B1 (.DIODE(_02424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06477__B1 (.DIODE(_02424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07769__S0 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07740__A (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07318__S0 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__A (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07271__S0 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07091__S0 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06993__S0 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06891__S0 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06551__S0 (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06479__A (.DIODE(_02427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07932__S (.DIODE(_02428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__S (.DIODE(_02428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07906__S0 (.DIODE(_02428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07210__S (.DIODE(_02428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07206__S (.DIODE(_02428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07184__S0 (.DIODE(_02428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06807__S (.DIODE(_02428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06803__S (.DIODE(_02428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06801__A (.DIODE(_02428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06482__A2 (.DIODE(_02428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07754__B (.DIODE(_02429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07740__B (.DIODE(_02429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07303__B (.DIODE(_02429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__B (.DIODE(_02429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07076__B (.DIODE(_02429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06976__B (.DIODE(_02429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06874__B (.DIODE(_02429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06543__A (.DIODE(_02429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06499__B (.DIODE(_02429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06481__A (.DIODE(_02429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08117__S1 (.DIODE(_02430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08027__S1 (.DIODE(_02430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07949__S1 (.DIODE(_02430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07921__B (.DIODE(_02430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07227__S1 (.DIODE(_02430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07199__B (.DIODE(_02430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06825__S1 (.DIODE(_02430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06791__B (.DIODE(_02430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06779__B (.DIODE(_02430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06482__A3 (.DIODE(_02430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__A (.DIODE(_02432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07969__A (.DIODE(_02432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__A (.DIODE(_02432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__S0 (.DIODE(_02432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07700__A (.DIODE(_02432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07610__A (.DIODE(_02432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07520__A (.DIODE(_02432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__A (.DIODE(_02432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07311__S0 (.DIODE(_02432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06485__A (.DIODE(_02432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__B (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07969__B (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07791__B (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07700__B (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07610__B (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07112__B (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07015__B (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06911__B (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06608__B (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06485__C_N (.DIODE(_02433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07869__A2 (.DIODE(_02437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07749__A2 (.DIODE(_02437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07739__A2 (.DIODE(_02437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07298__A2 (.DIODE(_02437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07287__A2 (.DIODE(_02437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07252__A2 (.DIODE(_02437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07071__A2 (.DIODE(_02437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06970__A2 (.DIODE(_02437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06863__A2 (.DIODE(_02437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06495__A2 (.DIODE(_02437_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07747__A2 (.DIODE(_02438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07737__A2 (.DIODE(_02438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07733__A2 (.DIODE(_02438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07296__A2 (.DIODE(_02438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07280__A2 (.DIODE(_02438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07250__A2 (.DIODE(_02438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07069__A2 (.DIODE(_02438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06967__A2 (.DIODE(_02438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06861__A2 (.DIODE(_02438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06491__A2 (.DIODE(_02438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08115__A1 (.DIODE(_02439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08025__A1 (.DIODE(_02439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07847__A1 (.DIODE(_02439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07737__B1 (.DIODE(_02439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07666__A1 (.DIODE(_02439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__B1 (.DIODE(_02439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06864__A (.DIODE(_02439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06714__A (.DIODE(_02439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06620__A (.DIODE(_02439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06491__B1 (.DIODE(_02439_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07748__A2 (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07524__A2 (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07434__A2 (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07344__A2 (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07251__A2 (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07070__A2 (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07009__A (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06969__A2 (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06862__A2 (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06494__A2 (.DIODE(_02441_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09781__A (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07919__B1 (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07748__B1 (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07738__B1 (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07297__B1 (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__B1 (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07148__A (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06862__B1 (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06707__A (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06494__B1 (.DIODE(_02442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__A2 (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07531__A2 (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07441__A2 (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07351__A2 (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07258__A2 (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07077__A2 (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06977__A2 (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06875__A2 (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06712__A (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06500__A2 (.DIODE(_02445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07711__B1 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__B1 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07531__B1 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07441__B1 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07351__B1 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07258__B1 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07077__B1 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06977__B1 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06875__B1 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06500__B1 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07754__A (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07530__A (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07440__A (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07350__A (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07257__A (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07076__A (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06976__A (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06874__A (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06542__A (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06499__A (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06502__B1 (.DIODE(_02449_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__A1 (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07807__A1 (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07742__C1 (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07626__A1 (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07291__C1 (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07263__A1 (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07128__A1 (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06790__B1 (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06648__A1 (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06502__C1 (.DIODE(_02450_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__A1 (.DIODE(_02453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07451__A (.DIODE(_02453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07361__A (.DIODE(_02453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07322__A1 (.DIODE(_02453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07268__A (.DIODE(_02453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07087__A (.DIODE(_02453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06990__A (.DIODE(_02453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06887__A (.DIODE(_02453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06732__A (.DIODE(_02453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06532__A (.DIODE(_02453_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08092__B1 (.DIODE(_02454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__B1 (.DIODE(_02454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07824__B1 (.DIODE(_02454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07643__B1 (.DIODE(_02454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07553__B1 (.DIODE(_02454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07463__B1 (.DIODE(_02454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07068__A (.DIODE(_02454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06703__A (.DIODE(_02454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06614__A (.DIODE(_02454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06506__A (.DIODE(_02454_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__A1 (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07747__B1 (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07733__B1 (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07313__B2 (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07296__B1 (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07280__B1 (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06967__B1 (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06861__B1 (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06647__A (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06507__A (.DIODE(_02455_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__B2 (.DIODE(_02456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__A1 (.DIODE(_02456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07985__A1 (.DIODE(_02456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07716__A1 (.DIODE(_02456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07536__A1 (.DIODE(_02456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07446__A1 (.DIODE(_02456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07356__A1 (.DIODE(_02456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07031__A1 (.DIODE(_02456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06928__A1 (.DIODE(_02456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06521__A1 (.DIODE(_02456_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07358__S0 (.DIODE(_02457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07265__S0 (.DIODE(_02457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07084__S0 (.DIODE(_02457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06987__S0 (.DIODE(_02457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06884__S0 (.DIODE(_02457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06879__A (.DIODE(_02457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06651__A (.DIODE(_02457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06641__A (.DIODE(_02457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06527__S0 (.DIODE(_02457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06509__A (.DIODE(_02457_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08120__S0 (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08030__S0 (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07852__S0 (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07671__S0 (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__S0 (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07491__S0 (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07401__S0 (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07129__S0 (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07032__S0 (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06513__S0 (.DIODE(_02458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08090__B (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08000__B (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07822__B (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07641__B (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06930__A (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06668__A (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06656__A (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06635__A (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06539__A (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06511__A (.DIODE(_02459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07760__S1 (.DIODE(_02460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07084__S1 (.DIODE(_02460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06987__S1 (.DIODE(_02460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06980__A (.DIODE(_02460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06884__S1 (.DIODE(_02460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06652__A (.DIODE(_02460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06642__A (.DIODE(_02460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06527__S1 (.DIODE(_02460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06519__A (.DIODE(_02460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06512__A (.DIODE(_02460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08120__S1 (.DIODE(_02461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08030__S1 (.DIODE(_02461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07852__S1 (.DIODE(_02461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07671__S1 (.DIODE(_02461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__S1 (.DIODE(_02461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07491__S1 (.DIODE(_02461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07401__S1 (.DIODE(_02461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07129__S1 (.DIODE(_02461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06880__S1 (.DIODE(_02461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06513__S1 (.DIODE(_02461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__B1 (.DIODE(_02463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08022__B1 (.DIODE(_02463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07844__B1 (.DIODE(_02463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07663__B1 (.DIODE(_02463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07573__B1 (.DIODE(_02463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07483__B1 (.DIODE(_02463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07393__B1 (.DIODE(_02463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07121__B1 (.DIODE(_02463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07024__B1 (.DIODE(_02463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06515__A (.DIODE(_02463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__C1 (.DIODE(_02464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08011__C1 (.DIODE(_02464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07833__C1 (.DIODE(_02464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__B2 (.DIODE(_02464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07652__C1 (.DIODE(_02464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07562__C1 (.DIODE(_02464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07472__C1 (.DIODE(_02464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__C1 (.DIODE(_02464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07313__A1 (.DIODE(_02464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06516__A (.DIODE(_02464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__B2 (.DIODE(_02465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07985__B2 (.DIODE(_02465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__B1 (.DIODE(_02465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07716__B2 (.DIODE(_02465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07536__B2 (.DIODE(_02465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07446__B2 (.DIODE(_02465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07356__B2 (.DIODE(_02465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07168__B1 (.DIODE(_02465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06928__B2 (.DIODE(_02465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06521__B1 (.DIODE(_02465_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08090__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08000__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07822__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07641__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07551__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07371__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07099__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07000__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06518__A (.DIODE(_02466_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08118__S0 (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08028__S0 (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07264__S0 (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07083__S0 (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06986__S0 (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06883__S0 (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06733__A (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06708__A (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06524__S0 (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06520__S0 (.DIODE(_02467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08118__S1 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08028__S1 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07447__S1 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07357__S1 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07264__S1 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07083__S1 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06986__S1 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06883__S1 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06524__S1 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06520__S1 (.DIODE(_02468_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07951__A1 (.DIODE(_02472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07450__A1 (.DIODE(_02472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07360__A1 (.DIODE(_02472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07267__A1 (.DIODE(_02472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07229__A1 (.DIODE(_02472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07086__A1 (.DIODE(_02472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06989__A1 (.DIODE(_02472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06886__A1 (.DIODE(_02472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06768__A (.DIODE(_02472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06531__A1 (.DIODE(_02472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__A (.DIODE(_02475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07759__A (.DIODE(_02475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07308__A (.DIODE(_02475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07266__A (.DIODE(_02475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07228__A (.DIODE(_02475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07085__A (.DIODE(_02475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06988__A (.DIODE(_02475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06885__A (.DIODE(_02475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06770__A (.DIODE(_02475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06528__A (.DIODE(_02475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07936__B1_N (.DIODE(_02479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__A1 (.DIODE(_02479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07360__C1 (.DIODE(_02479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__A1 (.DIODE(_02479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07267__C1 (.DIODE(_02479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07214__B1_N (.DIODE(_02479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07086__C1 (.DIODE(_02479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06989__C1 (.DIODE(_02479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06886__C1 (.DIODE(_02479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06531__C1 (.DIODE(_02479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06563__B1 (.DIODE(_02481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07638__A1 (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07548__A1 (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07458__A1 (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07368__A1 (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__A1 (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07095__A1 (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06997__A1 (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06895__A1 (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06690__A (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06562__A1 (.DIODE(_02482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08623__C (.DIODE(_02483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08125__A (.DIODE(_02483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06663__A (.DIODE(_02483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06535__A (.DIODE(_02483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12709__A (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12223__A (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11655__A (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11586__A (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11000__A (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10489__A (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__A1 (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07320__A1 (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07088__A (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06536__A (.DIODE(_02484_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08749__A (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__A1 (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07900__A1 (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07222__A1 (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07178__A1 (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06996__A1 (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06894__A1 (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06820__A1 (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06761__A1 (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06559__A1 (.DIODE(_02485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__A (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08009__A (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__A (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07751__A (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07744__A (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07650__A (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07300__A (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07293__A (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06664__A (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06538__A (.DIODE(_02486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07632__S0 (.DIODE(_02487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07542__S0 (.DIODE(_02487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07452__S0 (.DIODE(_02487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07362__S0 (.DIODE(_02487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07269__S0 (.DIODE(_02487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07089__S0 (.DIODE(_02487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06991__S0 (.DIODE(_02487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06888__S0 (.DIODE(_02487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06745__A (.DIODE(_02487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06541__S0 (.DIODE(_02487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__S1 (.DIODE(_02488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07758__S1 (.DIODE(_02488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07311__S1 (.DIODE(_02488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07309__S1 (.DIODE(_02488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07307__S1 (.DIODE(_02488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06983__A (.DIODE(_02488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06755__A (.DIODE(_02488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06665__A (.DIODE(_02488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06645__A (.DIODE(_02488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06540__A (.DIODE(_02488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__S1 (.DIODE(_02489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07868__B (.DIODE(_02489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07362__S1 (.DIODE(_02489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07269__S1 (.DIODE(_02489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07145__B (.DIODE(_02489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07089__S1 (.DIODE(_02489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06991__S1 (.DIODE(_02489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06888__S1 (.DIODE(_02489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06699__B (.DIODE(_02489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06541__S1 (.DIODE(_02489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07921__A (.DIODE(_02491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07453__S0 (.DIODE(_02491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__S0 (.DIODE(_02491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07270__S0 (.DIODE(_02491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07199__A (.DIODE(_02491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07090__S0 (.DIODE(_02491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06992__S0 (.DIODE(_02491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06889__S0 (.DIODE(_02491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06791__A (.DIODE(_02491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06544__S0 (.DIODE(_02491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09096__B (.DIODE(_02492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08955__B (.DIODE(_02492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08783__B (.DIODE(_02492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07871__C_N (.DIODE(_02492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__C_N (.DIODE(_02492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07090__S1 (.DIODE(_02492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06992__S1 (.DIODE(_02492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06889__S1 (.DIODE(_02492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06709__C_N (.DIODE(_02492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06544__S1 (.DIODE(_02492_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08855__A (.DIODE(_02495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08783__C (.DIODE(_02495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08371__A (.DIODE(_02495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__A (.DIODE(_02495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__B2 (.DIODE(_02495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07320__B2 (.DIODE(_02495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06937__A (.DIODE(_02495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06671__A (.DIODE(_02495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06547__A (.DIODE(_02495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__B2 (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07900__B2 (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07222__B2 (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07178__B2 (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07094__B2 (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06996__B2 (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06894__B2 (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06820__B2 (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06761__B2 (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06559__B2 (.DIODE(_02496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09025__A (.DIODE(_02497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08955__C (.DIODE(_02497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08298__A (.DIODE(_02497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06938__A (.DIODE(_02497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06754__A (.DIODE(_02497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06672__A (.DIODE(_02497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06549__A (.DIODE(_02497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11930__A (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11362__A (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11069__A (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10778__A (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07768__A1 (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07317__A1 (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07093__A1 (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06995__A1 (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06893__A1 (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06558__A1 (.DIODE(_02498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08129__S1 (.DIODE(_02499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08038__S1 (.DIODE(_02499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07860__S1 (.DIODE(_02499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07769__S1 (.DIODE(_02499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07679__S1 (.DIODE(_02499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07589__S1 (.DIODE(_02499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07499__S1 (.DIODE(_02499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07318__S1 (.DIODE(_02499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06734__A (.DIODE(_02499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06551__S1 (.DIODE(_02499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08121__S0 (.DIODE(_02501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08031__S0 (.DIODE(_02501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07853__S0 (.DIODE(_02501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07672__S0 (.DIODE(_02501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__S0 (.DIODE(_02501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07492__S0 (.DIODE(_02501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07402__S0 (.DIODE(_02501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07130__S0 (.DIODE(_02501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06697__A (.DIODE(_02501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06553__A (.DIODE(_02501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07770__S0 (.DIODE(_02502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07767__S0 (.DIODE(_02502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07766__S0 (.DIODE(_02502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__S0 (.DIODE(_02502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07316__S0 (.DIODE(_02502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07315__S0 (.DIODE(_02502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07092__S0 (.DIODE(_02502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06994__S0 (.DIODE(_02502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06892__S0 (.DIODE(_02502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06555__S0 (.DIODE(_02502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07766__S1 (.DIODE(_02503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07545__S1 (.DIODE(_02503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__S1 (.DIODE(_02503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07365__S1 (.DIODE(_02503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07315__S1 (.DIODE(_02503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07272__S1 (.DIODE(_02503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07092__S1 (.DIODE(_02503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06994__S1 (.DIODE(_02503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06892__S1 (.DIODE(_02503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06555__S1 (.DIODE(_02503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09166__A (.DIODE(_02505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09096__C (.DIODE(_02505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08209__A (.DIODE(_02505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06942__A (.DIODE(_02505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06759__A (.DIODE(_02505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06679__A (.DIODE(_02505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06557__A (.DIODE(_02505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12639__A (.DIODE(_02506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12500__A (.DIODE(_02506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12069__A (.DIODE(_02506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11500__A (.DIODE(_02506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07768__B2 (.DIODE(_02506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07317__B2 (.DIODE(_02506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07093__B2 (.DIODE(_02506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06995__B2 (.DIODE(_02506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06893__B2 (.DIODE(_02506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06558__B2 (.DIODE(_02506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06559__C1 (.DIODE(_02507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06562__A2 (.DIODE(_02508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08132__B1 (.DIODE(_02509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08041__B1 (.DIODE(_02509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__B1 (.DIODE(_02509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__C1 (.DIODE(_02509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07682__B1 (.DIODE(_02509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07592__B1 (.DIODE(_02509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07502__B1 (.DIODE(_02509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07322__C1 (.DIODE(_02509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06682__A (.DIODE(_02509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06561__A (.DIODE(_02509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07548__B1 (.DIODE(_02510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07458__B1 (.DIODE(_02510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07368__B1 (.DIODE(_02510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__B1 (.DIODE(_02510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07095__B1 (.DIODE(_02510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06997__B1 (.DIODE(_02510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06895__B1 (.DIODE(_02510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06813__B (.DIODE(_02510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06689__A (.DIODE(_02510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06562__B1 (.DIODE(_02510_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06563__B2 (.DIODE(_02511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08088__A1 (.DIODE(_02513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07998__A1 (.DIODE(_02513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07820__A1 (.DIODE(_02513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__A1 (.DIODE(_02513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07639__A1 (.DIODE(_02513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07413__A1 (.DIODE(_02513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07141__A1 (.DIODE(_02513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07045__A1 (.DIODE(_02513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06946__A1 (.DIODE(_02513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06684__A1 (.DIODE(_02513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08012__A (.DIODE(_02514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07834__A (.DIODE(_02514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07653__A (.DIODE(_02514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07563__A (.DIODE(_02514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07473__A (.DIODE(_02514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07383__A (.DIODE(_02514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07111__A (.DIODE(_02514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07014__A (.DIODE(_02514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06910__A (.DIODE(_02514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06602__A (.DIODE(_02514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08045__A2 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07955__A2 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07777__A2 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07686__A2 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07596__A2 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07506__A2 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07416__A2 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06999__A2 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06897__A2 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06568__A2 (.DIODE(_02515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08045__B1 (.DIODE(_02516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07955__B1 (.DIODE(_02516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07777__B1 (.DIODE(_02516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07686__B1 (.DIODE(_02516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07460__B1 (.DIODE(_02516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07370__B1 (.DIODE(_02516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07098__B1 (.DIODE(_02516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06999__B1 (.DIODE(_02516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06897__B1 (.DIODE(_02516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06568__B1 (.DIODE(_02516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08001__A2 (.DIODE(_02518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__A2 (.DIODE(_02518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07642__A2 (.DIODE(_02518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07552__A2 (.DIODE(_02518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07462__A2 (.DIODE(_02518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07372__A2 (.DIODE(_02518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07100__A2 (.DIODE(_02518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07001__A2 (.DIODE(_02518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06899__A2 (.DIODE(_02518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06574__A2 (.DIODE(_02518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__B1 (.DIODE(_02519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07957__B1 (.DIODE(_02519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07779__B1 (.DIODE(_02519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07552__B1 (.DIODE(_02519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07462__B1 (.DIODE(_02519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07372__B1 (.DIODE(_02519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07100__B1 (.DIODE(_02519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07001__B1 (.DIODE(_02519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06899__B1 (.DIODE(_02519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06574__B1 (.DIODE(_02519_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__A (.DIODE(_02520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07956__A (.DIODE(_02520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07778__A (.DIODE(_02520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07687__A (.DIODE(_02520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07597__A (.DIODE(_02520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07507__A (.DIODE(_02520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07417__A (.DIODE(_02520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07327__A (.DIODE(_02520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06898__A (.DIODE(_02520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06573__A (.DIODE(_02520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__A2 (.DIODE(_02524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07958__A2 (.DIODE(_02524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07780__A2 (.DIODE(_02524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07689__A2 (.DIODE(_02524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07599__A2 (.DIODE(_02524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__A2 (.DIODE(_02524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07101__A2 (.DIODE(_02524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07002__A2 (.DIODE(_02524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06900__A2 (.DIODE(_02524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06577__A2 (.DIODE(_02524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__B1 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07958__B1 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07780__B1 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07689__B1 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07599__B1 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07373__B1 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07101__B1 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07002__B1 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06900__B1 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06577__B1 (.DIODE(_02525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08050__A2 (.DIODE(_02527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07826__A2 (.DIODE(_02527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07645__A2 (.DIODE(_02527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07555__A2 (.DIODE(_02527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07465__A2 (.DIODE(_02527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07375__A2 (.DIODE(_02527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07103__A2 (.DIODE(_02527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07004__A2 (.DIODE(_02527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06902__A2 (.DIODE(_02527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06583__A2 (.DIODE(_02527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08050__B1 (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07960__B1 (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07782__B1 (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07691__B1 (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07601__B1 (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07511__B1 (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07421__B1 (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__B1 (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06902__B1 (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06583__B1 (.DIODE(_02528_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08049__A (.DIODE(_02529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07959__A (.DIODE(_02529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07781__A (.DIODE(_02529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07690__A (.DIODE(_02529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__A (.DIODE(_02529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07510__A (.DIODE(_02529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07102__A (.DIODE(_02529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07003__A (.DIODE(_02529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06901__A (.DIODE(_02529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06582__A (.DIODE(_02529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08049__C_N (.DIODE(_02530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07959__C_N (.DIODE(_02530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07644__C_N (.DIODE(_02530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__C_N (.DIODE(_02530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07464__C_N (.DIODE(_02530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07374__C_N (.DIODE(_02530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07102__C_N (.DIODE(_02530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07003__C_N (.DIODE(_02530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06901__C_N (.DIODE(_02530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06582__C_N (.DIODE(_02530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08054__A2 (.DIODE(_02534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07964__A2 (.DIODE(_02534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07649__A2 (.DIODE(_02534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07559__A2 (.DIODE(_02534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07469__A2 (.DIODE(_02534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07379__A2 (.DIODE(_02534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07107__A2 (.DIODE(_02534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07008__A2 (.DIODE(_02534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06906__A2 (.DIODE(_02534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06592__A2 (.DIODE(_02534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__A2 (.DIODE(_02535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07962__A2 (.DIODE(_02535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07647__A2 (.DIODE(_02535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07557__A2 (.DIODE(_02535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07467__A2 (.DIODE(_02535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07377__A2 (.DIODE(_02535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07105__A2 (.DIODE(_02535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07006__A2 (.DIODE(_02535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06904__A2 (.DIODE(_02535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06588__A2 (.DIODE(_02535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__B1 (.DIODE(_02536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07962__B1 (.DIODE(_02536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07784__B1 (.DIODE(_02536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07557__B1 (.DIODE(_02536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07467__B1 (.DIODE(_02536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07377__B1 (.DIODE(_02536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07105__B1 (.DIODE(_02536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07006__B1 (.DIODE(_02536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06904__B1 (.DIODE(_02536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06588__B1 (.DIODE(_02536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08053__A2 (.DIODE(_02538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07963__A2 (.DIODE(_02538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07558__A2 (.DIODE(_02538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07468__A2 (.DIODE(_02538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07378__A2 (.DIODE(_02538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07106__A2 (.DIODE(_02538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07007__A2 (.DIODE(_02538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06905__A2 (.DIODE(_02538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06604__A (.DIODE(_02538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06591__A2 (.DIODE(_02538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08053__B1 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07963__B1 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07785__B1 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07694__B1 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__B1 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07378__B1 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07106__B1 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07007__B1 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06905__B1 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06591__B1 (.DIODE(_02539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08057__A2 (.DIODE(_02542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07967__A2 (.DIODE(_02542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07789__A2 (.DIODE(_02542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07698__A2 (.DIODE(_02542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07608__A2 (.DIODE(_02542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07518__A2 (.DIODE(_02542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07428__A2 (.DIODE(_02542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07338__A2 (.DIODE(_02542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06909__A2 (.DIODE(_02542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06601__A2 (.DIODE(_02542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08056__A2 (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07966__A2 (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07788__A2 (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07697__A2 (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__A2 (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07517__A2 (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07427__A2 (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07337__A2 (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06908__A2 (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06599__A2 (.DIODE(_02543_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08056__B1 (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07966__B1 (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07788__B1 (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07697__B1 (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__B1 (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07517__B1 (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07427__B1 (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07012__B1 (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06908__B1 (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06599__B1 (.DIODE(_02544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08055__A (.DIODE(_02545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07965__A (.DIODE(_02545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07560__A (.DIODE(_02545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07470__A (.DIODE(_02545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07380__A (.DIODE(_02545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07108__A (.DIODE(_02545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07011__A (.DIODE(_02545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06907__A (.DIODE(_02545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06667__A (.DIODE(_02545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06598__A (.DIODE(_02545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08055__B (.DIODE(_02546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07965__B (.DIODE(_02546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__B (.DIODE(_02546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07560__B (.DIODE(_02546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07470__B (.DIODE(_02546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07380__B (.DIODE(_02546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07108__B (.DIODE(_02546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07011__B (.DIODE(_02546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06907__B (.DIODE(_02546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06598__B (.DIODE(_02546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08057__C1 (.DIODE(_02549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07967__C1 (.DIODE(_02549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07789__C1 (.DIODE(_02549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07698__C1 (.DIODE(_02549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07608__C1 (.DIODE(_02549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07518__C1 (.DIODE(_02549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__C1 (.DIODE(_02549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07013__C1 (.DIODE(_02549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06909__C1 (.DIODE(_02549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06601__C1 (.DIODE(_02549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06684__A2 (.DIODE(_02551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__A (.DIODE(_02552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07982__A (.DIODE(_02552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07667__A (.DIODE(_02552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07577__A (.DIODE(_02552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07487__A (.DIODE(_02552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07397__A (.DIODE(_02552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07125__A (.DIODE(_02552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07028__A (.DIODE(_02552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06925__A (.DIODE(_02552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06639__A (.DIODE(_02552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08061__A2 (.DIODE(_02553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07971__A2 (.DIODE(_02553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07793__A2 (.DIODE(_02553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07566__A2 (.DIODE(_02553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07476__A2 (.DIODE(_02553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07386__A2 (.DIODE(_02553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07114__A2 (.DIODE(_02553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07017__A2 (.DIODE(_02553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06913__A2 (.DIODE(_02553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06611__A2 (.DIODE(_02553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08060__A2 (.DIODE(_02554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07970__A2 (.DIODE(_02554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07792__A2 (.DIODE(_02554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07565__A2 (.DIODE(_02554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07475__A2 (.DIODE(_02554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07385__A2 (.DIODE(_02554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07113__A2 (.DIODE(_02554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07016__A2 (.DIODE(_02554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06912__A2 (.DIODE(_02554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06609__A2 (.DIODE(_02554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08014__B1 (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07836__B1 (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07655__B1 (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07565__B1 (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07475__B1 (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07385__B1 (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07113__B1 (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07016__B1 (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06912__B1 (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06609__B1 (.DIODE(_02555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08013__A (.DIODE(_02556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07835__A (.DIODE(_02556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07654__A (.DIODE(_02556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07564__A (.DIODE(_02556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07474__A (.DIODE(_02556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07384__A (.DIODE(_02556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07112__A (.DIODE(_02556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07015__A (.DIODE(_02556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06911__A (.DIODE(_02556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06608__A (.DIODE(_02556_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08061__C1 (.DIODE(_02559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07971__C1 (.DIODE(_02559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07793__C1 (.DIODE(_02559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07566__C1 (.DIODE(_02559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07476__C1 (.DIODE(_02559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07386__C1 (.DIODE(_02559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07114__C1 (.DIODE(_02559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07017__C1 (.DIODE(_02559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06913__C1 (.DIODE(_02559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06611__C1 (.DIODE(_02559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08064__A2 (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07974__A2 (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07796__A2 (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07705__A2 (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07615__A2 (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07525__A2 (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07435__A2 (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__A2 (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06916__A2 (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06619__A2 (.DIODE(_02561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08062__A2 (.DIODE(_02562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07972__A2 (.DIODE(_02562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__A2 (.DIODE(_02562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07703__A2 (.DIODE(_02562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07613__A2 (.DIODE(_02562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07523__A2 (.DIODE(_02562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07433__A2 (.DIODE(_02562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07343__A2 (.DIODE(_02562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06914__A2 (.DIODE(_02562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06615__A2 (.DIODE(_02562_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__B1 (.DIODE(_02563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07838__B1 (.DIODE(_02563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07657__B1 (.DIODE(_02563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07567__B1 (.DIODE(_02563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07477__B1 (.DIODE(_02563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07387__B1 (.DIODE(_02563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07115__B1 (.DIODE(_02563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07018__B1 (.DIODE(_02563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06914__B1 (.DIODE(_02563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06615__B1 (.DIODE(_02563_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08063__A2 (.DIODE(_02565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07973__A2 (.DIODE(_02565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__A2 (.DIODE(_02565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07730__A2 (.DIODE(_02565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07704__A2 (.DIODE(_02565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07614__A2 (.DIODE(_02565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07277__A2 (.DIODE(_02565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__A2 (.DIODE(_02565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06915__A2 (.DIODE(_02565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06618__A2 (.DIODE(_02565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08063__B1 (.DIODE(_02566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__B1 (.DIODE(_02566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07658__B1 (.DIODE(_02566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__B1 (.DIODE(_02566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07478__B1 (.DIODE(_02566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07388__B1 (.DIODE(_02566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07116__B1 (.DIODE(_02566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__B1 (.DIODE(_02566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06915__B1 (.DIODE(_02566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06618__B1 (.DIODE(_02566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08071__A1 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07981__A1 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07803__A1 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07576__A1 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07486__A1 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07396__A1 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__A1 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07027__A1 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06924__A1 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06638__A1 (.DIODE(_02569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08065__B (.DIODE(_02570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07841__B (.DIODE(_02570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07660__B (.DIODE(_02570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07570__B (.DIODE(_02570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07480__B (.DIODE(_02570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07390__B (.DIODE(_02570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07118__B (.DIODE(_02570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07021__B (.DIODE(_02570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06917__B (.DIODE(_02570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06622__B (.DIODE(_02570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08067__A2 (.DIODE(_02572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07977__A2 (.DIODE(_02572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__A2 (.DIODE(_02572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07708__A2 (.DIODE(_02572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07618__A2 (.DIODE(_02572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07392__A2 (.DIODE(_02572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07120__A2 (.DIODE(_02572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07023__A2 (.DIODE(_02572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06919__A2 (.DIODE(_02572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06628__A2 (.DIODE(_02572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08067__B1 (.DIODE(_02573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07977__B1 (.DIODE(_02573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__B1 (.DIODE(_02573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07708__B1 (.DIODE(_02573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07618__B1 (.DIODE(_02573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__B1 (.DIODE(_02573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07438__B1 (.DIODE(_02573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07023__B1 (.DIODE(_02573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06919__B1 (.DIODE(_02573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06628__B1 (.DIODE(_02573_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08066__A (.DIODE(_02574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07976__A (.DIODE(_02574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07798__A (.DIODE(_02574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07707__A (.DIODE(_02574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07481__A (.DIODE(_02574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__A (.DIODE(_02574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07119__A (.DIODE(_02574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07022__A (.DIODE(_02574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06918__A (.DIODE(_02574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06627__A (.DIODE(_02574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08066__C_N (.DIODE(_02575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07976__C_N (.DIODE(_02575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07661__C_N (.DIODE(_02575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07571__C_N (.DIODE(_02575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07481__C_N (.DIODE(_02575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07391__C_N (.DIODE(_02575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07119__C_N (.DIODE(_02575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07022__C_N (.DIODE(_02575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06918__C_N (.DIODE(_02575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06627__C_N (.DIODE(_02575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08068__B1 (.DIODE(_02579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07978__B1 (.DIODE(_02579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07800__B1 (.DIODE(_02579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07709__B1 (.DIODE(_02579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07619__B1 (.DIODE(_02579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07529__B1 (.DIODE(_02579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07439__B1 (.DIODE(_02579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07349__B1 (.DIODE(_02579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06920__B1 (.DIODE(_02579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06631__B1 (.DIODE(_02579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06638__B1 (.DIODE(_02580_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08070__A2 (.DIODE(_02581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07980__A2 (.DIODE(_02581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07802__A2 (.DIODE(_02581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07711__A2 (.DIODE(_02581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07485__A2 (.DIODE(_02581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07395__A2 (.DIODE(_02581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07123__A2 (.DIODE(_02581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07026__A2 (.DIODE(_02581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06923__A2 (.DIODE(_02581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06637__A2 (.DIODE(_02581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08070__B1 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07980__B1 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07802__B1 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07575__B1 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07485__B1 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07395__B1 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07123__B1 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07026__B1 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06923__B1 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06637__B1 (.DIODE(_02582_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08069__A (.DIODE(_02583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07979__A (.DIODE(_02583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07801__A (.DIODE(_02583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07710__A (.DIODE(_02583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07620__A (.DIODE(_02583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07394__A (.DIODE(_02583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07122__A (.DIODE(_02583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07025__A (.DIODE(_02583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06922__A (.DIODE(_02583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06636__A (.DIODE(_02583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08069__B (.DIODE(_02584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07979__B (.DIODE(_02584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07801__B (.DIODE(_02584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07710__B (.DIODE(_02584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07620__B (.DIODE(_02584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07530__B (.DIODE(_02584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07440__B (.DIODE(_02584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07350__B (.DIODE(_02584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07257__B (.DIODE(_02584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06636__B (.DIODE(_02584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06639__D (.DIODE(_02587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06684__A3 (.DIODE(_02588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08080__A (.DIODE(_02589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07990__A (.DIODE(_02589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07812__A (.DIODE(_02589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07721__A (.DIODE(_02589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07631__A (.DIODE(_02589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07541__A (.DIODE(_02589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07133__A (.DIODE(_02589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07036__A (.DIODE(_02589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06934__A (.DIODE(_02589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06661__A (.DIODE(_02589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08073__S0 (.DIODE(_02590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07983__S0 (.DIODE(_02590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07668__S0 (.DIODE(_02590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__S0 (.DIODE(_02590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07488__S0 (.DIODE(_02590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07398__S0 (.DIODE(_02590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07126__S0 (.DIODE(_02590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07029__S0 (.DIODE(_02590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06926__S0 (.DIODE(_02590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06643__S0 (.DIODE(_02590_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08073__S1 (.DIODE(_02591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07849__S1 (.DIODE(_02591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07668__S1 (.DIODE(_02591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__S1 (.DIODE(_02591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07488__S1 (.DIODE(_02591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07398__S1 (.DIODE(_02591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07126__S1 (.DIODE(_02591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07029__S1 (.DIODE(_02591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06926__S1 (.DIODE(_02591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06643__S1 (.DIODE(_02591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08074__S0 (.DIODE(_02593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07850__S0 (.DIODE(_02593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07669__S0 (.DIODE(_02593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07579__S0 (.DIODE(_02593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07489__S0 (.DIODE(_02593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07399__S0 (.DIODE(_02593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07127__S0 (.DIODE(_02593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07030__S0 (.DIODE(_02593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06927__S0 (.DIODE(_02593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06646__S0 (.DIODE(_02593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08074__S1 (.DIODE(_02594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07850__S1 (.DIODE(_02594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07669__S1 (.DIODE(_02594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07579__S1 (.DIODE(_02594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07489__S1 (.DIODE(_02594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07399__S1 (.DIODE(_02594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07127__S1 (.DIODE(_02594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07030__S1 (.DIODE(_02594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06927__S1 (.DIODE(_02594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06646__S1 (.DIODE(_02594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07870__B1 (.DIODE(_02596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07807__B2 (.DIODE(_02596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07626__B2 (.DIODE(_02596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07263__B2 (.DIODE(_02596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__B1 (.DIODE(_02596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07128__B2 (.DIODE(_02596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07082__B2 (.DIODE(_02596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06985__B2 (.DIODE(_02596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06882__B2 (.DIODE(_02596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06648__B2 (.DIODE(_02596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06661__B (.DIODE(_02597_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08079__A1 (.DIODE(_02599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07989__A1 (.DIODE(_02599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07811__A1 (.DIODE(_02599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07720__A1 (.DIODE(_02599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07630__A1 (.DIODE(_02599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07540__A1 (.DIODE(_02599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07132__A1 (.DIODE(_02599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07035__A1 (.DIODE(_02599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06933__A1 (.DIODE(_02599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06660__A1 (.DIODE(_02599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__S0 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__S0 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07808__S0 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07717__S0 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__S0 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07537__S0 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07447__S0 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07357__S0 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06929__S0 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06653__S0 (.DIODE(_02600_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__S1 (.DIODE(_02601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__S1 (.DIODE(_02601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07808__S1 (.DIODE(_02601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07717__S1 (.DIODE(_02601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__S1 (.DIODE(_02601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07537__S1 (.DIODE(_02601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07032__S1 (.DIODE(_02601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06929__S1 (.DIODE(_02601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06795__A (.DIODE(_02601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06653__S1 (.DIODE(_02601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06660__A2 (.DIODE(_02602_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08078__A (.DIODE(_02603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07988__A (.DIODE(_02603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07810__A (.DIODE(_02603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07719__A (.DIODE(_02603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__A (.DIODE(_02603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07539__A (.DIODE(_02603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07449__A (.DIODE(_02603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07359__A (.DIODE(_02603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06932__A (.DIODE(_02603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06658__A (.DIODE(_02603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08077__S0 (.DIODE(_02604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07987__S0 (.DIODE(_02604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07809__S0 (.DIODE(_02604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07718__S0 (.DIODE(_02604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07628__S0 (.DIODE(_02604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07538__S0 (.DIODE(_02604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07448__S0 (.DIODE(_02604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07033__S0 (.DIODE(_02604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06931__S0 (.DIODE(_02604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06657__S0 (.DIODE(_02604_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08077__S1 (.DIODE(_02605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07987__S1 (.DIODE(_02605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07809__S1 (.DIODE(_02605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07718__S1 (.DIODE(_02605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07628__S1 (.DIODE(_02605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07538__S1 (.DIODE(_02605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07448__S1 (.DIODE(_02605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07358__S1 (.DIODE(_02605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07265__S1 (.DIODE(_02605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06657__S1 (.DIODE(_02605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08079__C1 (.DIODE(_02608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07989__C1 (.DIODE(_02608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07811__C1 (.DIODE(_02608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07720__C1 (.DIODE(_02608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07630__C1 (.DIODE(_02608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07540__C1 (.DIODE(_02608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07450__C1 (.DIODE(_02608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07035__C1 (.DIODE(_02608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06933__C1 (.DIODE(_02608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06660__C1 (.DIODE(_02608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06684__B1 (.DIODE(_02610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08040__A1 (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07862__A1 (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07681__A1 (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07591__A1 (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07501__A1 (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07411__A1 (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07139__A1 (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07043__A1 (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06944__A1 (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06681__A1 (.DIODE(_02612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08081__S0 (.DIODE(_02613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07991__S0 (.DIODE(_02613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07813__S0 (.DIODE(_02613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07722__S0 (.DIODE(_02613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07496__S0 (.DIODE(_02613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__S0 (.DIODE(_02613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07134__S0 (.DIODE(_02613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07037__S0 (.DIODE(_02613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06935__S0 (.DIODE(_02613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06666__S0 (.DIODE(_02613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08081__S1 (.DIODE(_02614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07991__S1 (.DIODE(_02614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07813__S1 (.DIODE(_02614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07722__S1 (.DIODE(_02614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07632__S1 (.DIODE(_02614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07542__S1 (.DIODE(_02614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07452__S1 (.DIODE(_02614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07037__S1 (.DIODE(_02614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06935__S1 (.DIODE(_02614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06666__S1 (.DIODE(_02614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08082__S0 (.DIODE(_02616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07992__S0 (.DIODE(_02616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07814__S0 (.DIODE(_02616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__S0 (.DIODE(_02616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07633__S0 (.DIODE(_02616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07543__S0 (.DIODE(_02616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__S0 (.DIODE(_02616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07038__S0 (.DIODE(_02616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06936__S0 (.DIODE(_02616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06670__S0 (.DIODE(_02616_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09166__C_N (.DIODE(_02617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09025__C_N (.DIODE(_02617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08623__B (.DIODE(_02617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08128__S1 (.DIODE(_02617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08037__S1 (.DIODE(_02617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07859__S1 (.DIODE(_02617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__S1 (.DIODE(_02617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07312__S1 (.DIODE(_02617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06798__A (.DIODE(_02617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06669__A (.DIODE(_02617_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__S1 (.DIODE(_02618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07858__S1 (.DIODE(_02618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07677__S1 (.DIODE(_02618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07587__S1 (.DIODE(_02618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07497__S1 (.DIODE(_02618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07407__S1 (.DIODE(_02618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__S1 (.DIODE(_02618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07038__S1 (.DIODE(_02618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06936__S1 (.DIODE(_02618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06670__S1 (.DIODE(_02618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06681__B1 (.DIODE(_02619_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08086__B2 (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07996__B2 (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07818__B2 (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07727__B2 (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07637__B2 (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__B2 (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__B2 (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07367__B2 (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07274__B2 (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06681__B2 (.DIODE(_02620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__A1 (.DIODE(_02621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07995__A1 (.DIODE(_02621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07817__A1 (.DIODE(_02621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07726__A1 (.DIODE(_02621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07636__A1 (.DIODE(_02621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07546__A1 (.DIODE(_02621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07456__A1 (.DIODE(_02621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07366__A1 (.DIODE(_02621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07273__A1 (.DIODE(_02621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06680__A1 (.DIODE(_02621_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08083__S0 (.DIODE(_02622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07993__S0 (.DIODE(_02622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07815__S0 (.DIODE(_02622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07724__S0 (.DIODE(_02622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07634__S0 (.DIODE(_02622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07544__S0 (.DIODE(_02622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07454__S0 (.DIODE(_02622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07364__S0 (.DIODE(_02622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06939__S0 (.DIODE(_02622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06675__S0 (.DIODE(_02622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08083__S1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07993__S1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__S1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07588__S1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07498__S1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07408__S1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07136__S1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07040__S1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06939__S1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06675__S1 (.DIODE(_02623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08084__S0 (.DIODE(_02625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07994__S0 (.DIODE(_02625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07816__S0 (.DIODE(_02625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__S0 (.DIODE(_02625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07635__S0 (.DIODE(_02625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07545__S0 (.DIODE(_02625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__S0 (.DIODE(_02625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07365__S0 (.DIODE(_02625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07272__S0 (.DIODE(_02625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06678__S0 (.DIODE(_02625_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08084__S1 (.DIODE(_02626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07994__S1 (.DIODE(_02626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07816__S1 (.DIODE(_02626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__S1 (.DIODE(_02626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07635__S1 (.DIODE(_02626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07409__S1 (.DIODE(_02626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07137__S1 (.DIODE(_02626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07041__S1 (.DIODE(_02626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06941__S1 (.DIODE(_02626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06678__S1 (.DIODE(_02626_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__B2 (.DIODE(_02628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07995__B2 (.DIODE(_02628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07817__B2 (.DIODE(_02628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07726__B2 (.DIODE(_02628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07636__B2 (.DIODE(_02628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07546__B2 (.DIODE(_02628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07456__B2 (.DIODE(_02628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07366__B2 (.DIODE(_02628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07273__B2 (.DIODE(_02628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06680__B2 (.DIODE(_02628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06681__C1 (.DIODE(_02629_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06684__B2 (.DIODE(_02632_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__S (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08043__S (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07938__C1 (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07865__S (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07775__S (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07684__S (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07594__S (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07216__C1 (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06814__C1 (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06686__A (.DIODE(_02634_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07954__A1_N (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07504__S (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07414__S (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07324__S (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07232__A1_N (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07142__S (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07046__S (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06947__S (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06830__A1_N (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06687__S (.DIODE(_02635_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07953__C1 (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__A1 (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07909__B1 (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07231__C1 (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07188__A1 (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07187__B1 (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06829__C1 (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06777__B (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06776__A1 (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06775__B1 (.DIODE(_02637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07953__A1 (.DIODE(_02638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__A (.DIODE(_02638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07880__A (.DIODE(_02638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07231__A1 (.DIODE(_02638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07179__A (.DIODE(_02638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07158__A (.DIODE(_02638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06829__A1 (.DIODE(_02638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06777__A (.DIODE(_02638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06762__A (.DIODE(_02638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06731__A (.DIODE(_02638_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__B (.DIODE(_02639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08105__A2 (.DIODE(_02639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08015__A2 (.DIODE(_02639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07919__A2 (.DIODE(_02639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07837__A2 (.DIODE(_02639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07656__A2 (.DIODE(_02639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07197__A2 (.DIODE(_02639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06787__A2 (.DIODE(_02639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06706__A (.DIODE(_02639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06692__A (.DIODE(_02639_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__A2 (.DIODE(_02640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07885__A2 (.DIODE(_02640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07875__A2 (.DIODE(_02640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07191__A2 (.DIODE(_02640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07163__A2 (.DIODE(_02640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07153__A2 (.DIODE(_02640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__A2 (.DIODE(_02640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06739__A2 (.DIODE(_02640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06719__A2 (.DIODE(_02640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06694__A2 (.DIODE(_02640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07913__C1 (.DIODE(_02641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07883__C1 (.DIODE(_02641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07867__B1 (.DIODE(_02641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07295__C1 (.DIODE(_02641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07191__C1 (.DIODE(_02641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07161__C1 (.DIODE(_02641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07144__B1 (.DIODE(_02641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06781__C1 (.DIODE(_02641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06737__C1 (.DIODE(_02641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06694__B1 (.DIODE(_02641_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07892__A2 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__A2 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07878__A2 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07170__A2 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07160__A2 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07156__A2 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07146__A2 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06736__A2 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06728__A2 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06700__A2 (.DIODE(_02643_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12639__B (.DIODE(_02644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12500__B (.DIODE(_02644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12223__B (.DIODE(_02644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12069__B (.DIODE(_02644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11930__B (.DIODE(_02644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07869__B1 (.DIODE(_02644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07193__B1 (.DIODE(_02644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07146__B1 (.DIODE(_02644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06783__B1 (.DIODE(_02644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06700__B1 (.DIODE(_02644_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09166__B (.DIODE(_02645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09025__B (.DIODE(_02645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08623__A (.DIODE(_02645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08117__S0 (.DIODE(_02645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08027__S0 (.DIODE(_02645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07949__S0 (.DIODE(_02645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07849__S0 (.DIODE(_02645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07227__S0 (.DIODE(_02645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06825__S0 (.DIODE(_02645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06698__A (.DIODE(_02645_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__S0 (.DIODE(_02646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07871__A (.DIODE(_02646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07868__A (.DIODE(_02646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__S0 (.DIODE(_02646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07145__A (.DIODE(_02646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06796__S0 (.DIODE(_02646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06771__S0 (.DIODE(_02646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06763__A (.DIODE(_02646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06750__A (.DIODE(_02646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06699__A (.DIODE(_02646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07917__B (.DIODE(_02649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__A2 (.DIODE(_02649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07887__B (.DIODE(_02649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__A2 (.DIODE(_02649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__B (.DIODE(_02649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07192__A2 (.DIODE(_02649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07165__B (.DIODE(_02649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06785__B (.DIODE(_02649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06782__A2 (.DIODE(_02649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06702__A (.DIODE(_02649_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07884__A2 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__A2 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07870__A2 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07162__A2 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__A2 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__A2 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06741__B (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06738__A2 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06715__A2 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06705__A2 (.DIODE(_02650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08029__A1 (.DIODE(_02651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07914__B1 (.DIODE(_02651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07851__A1 (.DIODE(_02651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07670__A1 (.DIODE(_02651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07580__A1 (.DIODE(_02651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07490__A1 (.DIODE(_02651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07400__A1 (.DIODE(_02651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07192__B1 (.DIODE(_02651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06782__B1 (.DIODE(_02651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06704__A (.DIODE(_02651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07947__B2 (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__B2 (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07884__B1 (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07225__B2 (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07182__B2 (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07162__B1 (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06823__A1 (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06767__A1 (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06738__B1 (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06705__B1 (.DIODE(_02652_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08662__B (.DIODE(_02654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08517__B (.DIODE(_02654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__B (.DIODE(_02654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__A2 (.DIODE(_02654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07872__A2 (.DIODE(_02654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07867__A2 (.DIODE(_02654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07167__A2 (.DIODE(_02654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__A2 (.DIODE(_02654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06743__A2 (.DIODE(_02654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06710__A2 (.DIODE(_02654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__B1 (.DIODE(_02655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07882__B1 (.DIODE(_02655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07878__B1 (.DIODE(_02655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07167__B1 (.DIODE(_02655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07160__B1 (.DIODE(_02655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07156__B1 (.DIODE(_02655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06743__B1 (.DIODE(_02655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06736__B1 (.DIODE(_02655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06728__B1 (.DIODE(_02655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06710__B1 (.DIODE(_02655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09096__A (.DIODE(_02656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08955__A (.DIODE(_02656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08783__A (.DIODE(_02656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07948__S0 (.DIODE(_02656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07945__S0 (.DIODE(_02656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07226__S0 (.DIODE(_02656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07223__S0 (.DIODE(_02656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__A (.DIODE(_02656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06821__S0 (.DIODE(_02656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06709__A (.DIODE(_02656_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08098__A2 (.DIODE(_02660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08008__A2 (.DIODE(_02660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07922__A2 (.DIODE(_02660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07912__A2 (.DIODE(_02660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07830__A2 (.DIODE(_02660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07200__A2 (.DIODE(_02660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07190__A2 (.DIODE(_02660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06792__A2 (.DIODE(_02660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06780__A2 (.DIODE(_02660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06713__A (.DIODE(_02660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__A2 (.DIODE(_02661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07886__A2 (.DIODE(_02661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07876__A2 (.DIODE(_02661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07194__A2 (.DIODE(_02661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07164__A2 (.DIODE(_02661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07154__A2 (.DIODE(_02661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06784__A2 (.DIODE(_02661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06747__A2 (.DIODE(_02661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06740__A2 (.DIODE(_02661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06720__A2 (.DIODE(_02661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07923__A1 (.DIODE(_02662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__A1 (.DIODE(_02662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__B1 (.DIODE(_02662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07305__A1 (.DIODE(_02662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__A1 (.DIODE(_02662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__A1 (.DIODE(_02662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07152__B1 (.DIODE(_02662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06793__A1 (.DIODE(_02662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06748__A1 (.DIODE(_02662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06715__B1 (.DIODE(_02662_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08100__B1 (.DIODE(_02664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08010__B1 (.DIODE(_02664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07832__B1 (.DIODE(_02664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07651__B1 (.DIODE(_02664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07561__B1 (.DIODE(_02664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07471__B1 (.DIODE(_02664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07381__B1 (.DIODE(_02664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07301__B1 (.DIODE(_02664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07109__B1 (.DIODE(_02664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06717__A (.DIODE(_02664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07922__B1 (.DIODE(_02665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07915__B1 (.DIODE(_02665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07912__B1 (.DIODE(_02665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07200__B1 (.DIODE(_02665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07197__B1 (.DIODE(_02665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07190__B1 (.DIODE(_02665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06792__B1 (.DIODE(_02665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06787__B1 (.DIODE(_02665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06780__B1 (.DIODE(_02665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06718__A (.DIODE(_02665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08749__B (.DIODE(_02666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07892__B1 (.DIODE(_02666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07885__B1 (.DIODE(_02666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07875__B1 (.DIODE(_02666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07170__B1 (.DIODE(_02666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07163__B1 (.DIODE(_02666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07153__B1 (.DIODE(_02666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06747__B1 (.DIODE(_02666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06739__B1 (.DIODE(_02666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06719__B1 (.DIODE(_02666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__A2 (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07883__A2 (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07879__A2 (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07168__A2 (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07161__A2 (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__A2 (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06781__A2 (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06744__A2 (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06737__A2 (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06730__A2 (.DIODE(_02669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08093__A (.DIODE(_02670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08003__A (.DIODE(_02670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07825__A (.DIODE(_02670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07758__S0 (.DIODE(_02670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07644__A (.DIODE(_02670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07554__A (.DIODE(_02670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07464__A (.DIODE(_02670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07374__A (.DIODE(_02670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07307__S0 (.DIODE(_02670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06723__A (.DIODE(_02670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__S0 (.DIODE(_02671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08035__S0 (.DIODE(_02671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__A (.DIODE(_02671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__S0 (.DIODE(_02671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07676__S0 (.DIODE(_02671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07586__S0 (.DIODE(_02671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07196__A (.DIODE(_02671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06881__S0 (.DIODE(_02671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06786__A (.DIODE(_02671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06724__A (.DIODE(_02671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__S0 (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07888__A (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07877__A (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07176__S0 (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07166__A (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07155__A (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06822__S0 (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06758__S0 (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06742__A (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06727__A (.DIODE(_02672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07918__C_N (.DIODE(_02673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__B (.DIODE(_02673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07770__S1 (.DIODE(_02673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07767__S1 (.DIODE(_02673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__S1 (.DIODE(_02673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07316__S1 (.DIODE(_02673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07196__C_N (.DIODE(_02673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07189__B (.DIODE(_02673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06786__C_N (.DIODE(_02673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06726__A (.DIODE(_02673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08698__B (.DIODE(_02674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__S1 (.DIODE(_02674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07906__S1 (.DIODE(_02674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__B (.DIODE(_02674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07184__S1 (.DIODE(_02674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07169__B (.DIODE(_02674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06771__S1 (.DIODE(_02674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06751__A (.DIODE(_02674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06746__B (.DIODE(_02674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06727__B (.DIODE(_02674_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07947__A1 (.DIODE(_02677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__A1 (.DIODE(_02677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07879__C1 (.DIODE(_02677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07225__A1 (.DIODE(_02677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07182__A1 (.DIODE(_02677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__C1 (.DIODE(_02677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06823__B2 (.DIODE(_02677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06767__B2 (.DIODE(_02677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06744__B1 (.DIODE(_02677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06730__C1 (.DIODE(_02677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06776__A2 (.DIODE(_02679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07952__A (.DIODE(_02680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07909__A1 (.DIODE(_02680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07894__A (.DIODE(_02680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07230__A (.DIODE(_02680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07187__A1 (.DIODE(_02680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07172__A (.DIODE(_02680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06828__A (.DIODE(_02680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06813__A (.DIODE(_02680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06775__A1 (.DIODE(_02680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06749__A (.DIODE(_02680_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08855__B (.DIODE(_02681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07946__S0 (.DIODE(_02681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07897__S0 (.DIODE(_02681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07881__A (.DIODE(_02681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07224__S0 (.DIODE(_02681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07175__S0 (.DIODE(_02681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07159__A (.DIODE(_02681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06824__S0 (.DIODE(_02681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06757__S0 (.DIODE(_02681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06735__A (.DIODE(_02681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08855__C_N (.DIODE(_02682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07888__C_N (.DIODE(_02682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07881__B (.DIODE(_02682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07877__B (.DIODE(_02682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07166__C_N (.DIODE(_02682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07159__B (.DIODE(_02682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07155__B (.DIODE(_02682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06764__A (.DIODE(_02682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06742__C_N (.DIODE(_02682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06735__B (.DIODE(_02682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07942__S0 (.DIODE(_02693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07941__S0 (.DIODE(_02693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07935__S0 (.DIODE(_02693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__A (.DIODE(_02693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07219__S0 (.DIODE(_02693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07213__S0 (.DIODE(_02693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07169__A (.DIODE(_02693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06817__S0 (.DIODE(_02693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06810__S0 (.DIODE(_02693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06746__A (.DIODE(_02693_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06776__A3 (.DIODE(_02697_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07940__S0 (.DIODE(_02698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07939__S0 (.DIODE(_02698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__S0 (.DIODE(_02698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__S0 (.DIODE(_02698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07217__S0 (.DIODE(_02698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07174__S0 (.DIODE(_02698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06816__S0 (.DIODE(_02698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06815__S0 (.DIODE(_02698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06753__S0 (.DIODE(_02698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06752__S0 (.DIODE(_02698_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07939__S1 (.DIODE(_02699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__S1 (.DIODE(_02699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07895__S1 (.DIODE(_02699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07217__S1 (.DIODE(_02699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07181__S1 (.DIODE(_02699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07174__S1 (.DIODE(_02699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07173__S1 (.DIODE(_02699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06766__S1 (.DIODE(_02699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06753__S1 (.DIODE(_02699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06752__S1 (.DIODE(_02699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10212__A (.DIODE(_02702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09061__A (.DIODE(_02702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08553__A (.DIODE(_02702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08410__A (.DIODE(_02702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07943__A1 (.DIODE(_02702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__A1 (.DIODE(_02702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07221__A1 (.DIODE(_02702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07177__A1 (.DIODE(_02702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06819__A1 (.DIODE(_02702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06760__A1 (.DIODE(_02702_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__S1 (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08035__S1 (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__S1 (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07676__S1 (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07586__S1 (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07496__S1 (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07406__S1 (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07134__S1 (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06881__S1 (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06756__A (.DIODE(_02703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07946__S1 (.DIODE(_02704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07935__S1 (.DIODE(_02704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__S1 (.DIODE(_02704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07224__S1 (.DIODE(_02704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07213__S1 (.DIODE(_02704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07176__S1 (.DIODE(_02704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06822__S1 (.DIODE(_02704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06810__S1 (.DIODE(_02704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06758__S1 (.DIODE(_02704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06757__S1 (.DIODE(_02704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10916__A (.DIODE(_02707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09782__A (.DIODE(_02707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09202__A (.DIODE(_02707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08263__A (.DIODE(_02707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07943__B2 (.DIODE(_02707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__B2 (.DIODE(_02707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07221__B2 (.DIODE(_02707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07177__B2 (.DIODE(_02707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06819__B2 (.DIODE(_02707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06760__B2 (.DIODE(_02707_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06762__B (.DIODE(_02709_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07905__S0 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07903__S0 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07895__S0 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07183__S0 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07181__S0 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__S0 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07173__S0 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06769__S0 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06766__S0 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06765__S0 (.DIODE(_02711_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07933__A_N (.DIODE(_02712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07905__S1 (.DIODE(_02712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07903__S1 (.DIODE(_02712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07902__S1 (.DIODE(_02712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07211__A_N (.DIODE(_02712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07183__S1 (.DIODE(_02712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__S1 (.DIODE(_02712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06808__A_N (.DIODE(_02712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06769__S1 (.DIODE(_02712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06765__S1 (.DIODE(_02712_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06775__A2 (.DIODE(_02715_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07934__C1 (.DIODE(_02716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07930__C1 (.DIODE(_02716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07908__A1 (.DIODE(_02716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07212__C1 (.DIODE(_02716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07208__C1 (.DIODE(_02716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07186__A1 (.DIODE(_02716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06827__A1 (.DIODE(_02716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06809__C1 (.DIODE(_02716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06805__C1 (.DIODE(_02716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06774__A1 (.DIODE(_02716_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07936__A1 (.DIODE(_02718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07926__A (.DIODE(_02718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07907__A (.DIODE(_02718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07214__A1 (.DIODE(_02718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07204__A (.DIODE(_02718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07185__A (.DIODE(_02718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06826__A (.DIODE(_02718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06811__A1 (.DIODE(_02718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06797__A (.DIODE(_02718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06772__A (.DIODE(_02718_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07951__C1 (.DIODE(_02721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07937__A1 (.DIODE(_02721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07908__C1 (.DIODE(_02721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07229__C1 (.DIODE(_02721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07215__A1 (.DIODE(_02721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07186__C1 (.DIODE(_02721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06827__C1 (.DIODE(_02721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06812__A1 (.DIODE(_02721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06811__B1_N (.DIODE(_02721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06774__C1 (.DIODE(_02721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__S0 (.DIODE(_02726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__S0 (.DIODE(_02726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07911__A (.DIODE(_02726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07858__S0 (.DIODE(_02726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07677__S0 (.DIODE(_02726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07587__S0 (.DIODE(_02726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07497__S0 (.DIODE(_02726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07407__S0 (.DIODE(_02726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07189__A (.DIODE(_02726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06779__A (.DIODE(_02726_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07735__A2 (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__A2 (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07438__A2 (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07348__A2 (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07283__A2 (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07255__A2 (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07074__A2 (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06974__A2 (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06871__A2 (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06789__A (.DIODE(_02736_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12709__B (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11586__B (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11000__B (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10420__B (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09851__B (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07920__A2 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07742__A2 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07291__A2 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07198__A2 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06790__A2 (.DIODE(_02737_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06814__A2 (.DIODE(_02742_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07948__S1 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07945__S1 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07897__S1 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07226__S1 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07223__S1 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__S1 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07175__S1 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06824__S1 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06821__S1 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06796__S1 (.DIODE(_02743_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08082__S1 (.DIODE(_02746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07992__S1 (.DIODE(_02746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07814__S1 (.DIODE(_02746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__S1 (.DIODE(_02746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07633__S1 (.DIODE(_02746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07543__S1 (.DIODE(_02746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07453__S1 (.DIODE(_02746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__S1 (.DIODE(_02746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07270__S1 (.DIODE(_02746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06799__A (.DIODE(_02746_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07942__S1 (.DIODE(_02747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07941__S1 (.DIODE(_02747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07929__A_N (.DIODE(_02747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__S1 (.DIODE(_02747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07219__S1 (.DIODE(_02747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07207__A_N (.DIODE(_02747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06818__S1 (.DIODE(_02747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06817__S1 (.DIODE(_02747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06804__A_N (.DIODE(_02747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06800__A (.DIODE(_02747_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07940__S1 (.DIODE(_02748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07934__A1 (.DIODE(_02748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07930__A1 (.DIODE(_02748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__S1 (.DIODE(_02748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07212__A1 (.DIODE(_02748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07208__A1 (.DIODE(_02748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06816__S1 (.DIODE(_02748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06815__S1 (.DIODE(_02748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06809__A1 (.DIODE(_02748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06805__A1 (.DIODE(_02748_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08698__A_N (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07931__S (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07927__S (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07902__S0 (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__S0 (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07209__S (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07205__S (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06818__S0 (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06806__S (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06802__S (.DIODE(_02749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06809__A2 (.DIODE(_02754_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06830__B2 (.DIODE(_02777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07778__B (.DIODE(_02779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07687__B (.DIODE(_02779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07597__B (.DIODE(_02779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07507__B (.DIODE(_02779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07417__B (.DIODE(_02779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07327__B (.DIODE(_02779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07234__B (.DIODE(_02779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07051__B (.DIODE(_02779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06950__B (.DIODE(_02779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06833__B (.DIODE(_02779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07781__C_N (.DIODE(_02783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07690__C_N (.DIODE(_02783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__C_N (.DIODE(_02783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07510__C_N (.DIODE(_02783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07420__C_N (.DIODE(_02783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07330__C_N (.DIODE(_02783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07237__C_N (.DIODE(_02783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07054__C_N (.DIODE(_02783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06954__C_N (.DIODE(_02783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06837__C_N (.DIODE(_02783_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07786__A2 (.DIODE(_02787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07695__A2 (.DIODE(_02787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07605__A2 (.DIODE(_02787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07515__A2 (.DIODE(_02787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07425__A2 (.DIODE(_02787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07335__A2 (.DIODE(_02787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07242__A2 (.DIODE(_02787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07059__A2 (.DIODE(_02787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06959__A2 (.DIODE(_02787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06845__A2 (.DIODE(_02787_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07784__A2 (.DIODE(_02788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07693__A2 (.DIODE(_02788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__A2 (.DIODE(_02788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07513__A2 (.DIODE(_02788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07423__A2 (.DIODE(_02788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__A2 (.DIODE(_02788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07240__A2 (.DIODE(_02788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07057__A2 (.DIODE(_02788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06957__A2 (.DIODE(_02788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06842__A2 (.DIODE(_02788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07785__A2 (.DIODE(_02790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07694__A2 (.DIODE(_02790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__A2 (.DIODE(_02790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07514__A2 (.DIODE(_02790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07424__A2 (.DIODE(_02790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07334__A2 (.DIODE(_02790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07241__A2 (.DIODE(_02790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07058__A2 (.DIODE(_02790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06958__A2 (.DIODE(_02790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06844__A2 (.DIODE(_02790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07787__A (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07696__A (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07606__A (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07516__A (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07426__A (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07336__A (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07243__A (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07060__A (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06960__A (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06847__A (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06896__A2 (.DIODE(_02797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07804__A (.DIODE(_02798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07713__A (.DIODE(_02798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07623__A (.DIODE(_02798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07533__A (.DIODE(_02798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07443__A (.DIODE(_02798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07353__A (.DIODE(_02798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07260__A (.DIODE(_02798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07079__A (.DIODE(_02798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06979__A (.DIODE(_02798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06877__A (.DIODE(_02798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07746__A2 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__A2 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07612__A2 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07522__A2 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07432__A2 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07342__A2 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07249__A2 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07067__A2 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06966__A2 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06860__A2 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07745__A2 (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07701__A2 (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__A2 (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07521__A2 (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07431__A2 (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07341__A2 (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07248__A2 (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07066__A2 (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__A2 (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06858__A2 (.DIODE(_02800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08111__B1 (.DIODE(_02801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08021__B1 (.DIODE(_02801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07843__B1 (.DIODE(_02801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07662__B1 (.DIODE(_02801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07572__B1 (.DIODE(_02801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07482__B1 (.DIODE(_02801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07392__B1 (.DIODE(_02801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07120__B1 (.DIODE(_02801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__B1 (.DIODE(_02801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06858__B1 (.DIODE(_02801_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08110__A (.DIODE(_02802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08020__A (.DIODE(_02802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07842__A (.DIODE(_02802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07661__A (.DIODE(_02802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07571__A (.DIODE(_02802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07340__A (.DIODE(_02802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07247__A (.DIODE(_02802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07065__A (.DIODE(_02802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06964__A (.DIODE(_02802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06857__A (.DIODE(_02802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08110__C_N (.DIODE(_02803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08020__C_N (.DIODE(_02803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07842__C_N (.DIODE(_02803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07520__B (.DIODE(_02803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__B (.DIODE(_02803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07340__B (.DIODE(_02803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07247__B (.DIODE(_02803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07065__B (.DIODE(_02803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06964__B (.DIODE(_02803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06857__B (.DIODE(_02803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06860__B1 (.DIODE(_02805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07746__C1 (.DIODE(_02806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__C1 (.DIODE(_02806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07612__C1 (.DIODE(_02806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07522__C1 (.DIODE(_02806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07432__C1 (.DIODE(_02806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07342__C1 (.DIODE(_02806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07249__C1 (.DIODE(_02806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07067__C1 (.DIODE(_02806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06966__C1 (.DIODE(_02806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06860__C1 (.DIODE(_02806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07756__A1 (.DIODE(_02811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__A1 (.DIODE(_02811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07622__A1 (.DIODE(_02811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07532__A1 (.DIODE(_02811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__A1 (.DIODE(_02811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07352__A1 (.DIODE(_02811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07259__A1 (.DIODE(_02811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07078__A1 (.DIODE(_02811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06978__A1 (.DIODE(_02811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06876__A1 (.DIODE(_02811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08092__A2 (.DIODE(_02812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__A2 (.DIODE(_02812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07824__A2 (.DIODE(_02812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07750__B (.DIODE(_02812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07643__A2 (.DIODE(_02812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07553__A2 (.DIODE(_02812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07463__A2 (.DIODE(_02812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07373__A2 (.DIODE(_02812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07299__B (.DIODE(_02812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06866__B (.DIODE(_02812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07752__B1 (.DIODE(_02814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07745__B1 (.DIODE(_02814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07735__B1 (.DIODE(_02814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07348__B1 (.DIODE(_02814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07294__B1 (.DIODE(_02814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07283__B1 (.DIODE(_02814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07255__B1 (.DIODE(_02814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07074__B1 (.DIODE(_02814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06974__B1 (.DIODE(_02814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06871__B1 (.DIODE(_02814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07734__A (.DIODE(_02815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07617__A (.DIODE(_02815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07527__A (.DIODE(_02815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07437__A (.DIODE(_02815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07347__A (.DIODE(_02815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07282__A (.DIODE(_02815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07254__A (.DIODE(_02815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07073__A (.DIODE(_02815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06973__A (.DIODE(_02815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06870__A (.DIODE(_02815_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07798__C_N (.DIODE(_02816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07707__C_N (.DIODE(_02816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07617__C_N (.DIODE(_02816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07527__C_N (.DIODE(_02816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07437__C_N (.DIODE(_02816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07347__C_N (.DIODE(_02816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07254__C_N (.DIODE(_02816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07073__C_N (.DIODE(_02816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06973__C_N (.DIODE(_02816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06870__C_N (.DIODE(_02816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07753__A2 (.DIODE(_02819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07619__A2 (.DIODE(_02819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07529__A2 (.DIODE(_02819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07439__A2 (.DIODE(_02819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07349__A2 (.DIODE(_02819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07302__A2 (.DIODE(_02819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__A2 (.DIODE(_02819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07075__A2 (.DIODE(_02819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06975__A2 (.DIODE(_02819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06873__A2 (.DIODE(_02819_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06876__B2 (.DIODE(_02822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06877__D (.DIODE(_02823_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08029__B2 (.DIODE(_02825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07851__B2 (.DIODE(_02825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07670__B2 (.DIODE(_02825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07580__B2 (.DIODE(_02825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07490__B2 (.DIODE(_02825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07400__B2 (.DIODE(_02825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07082__A1 (.DIODE(_02825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07031__B2 (.DIODE(_02825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06985__A1 (.DIODE(_02825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06882__A1 (.DIODE(_02825_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07805__S0 (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07714__S0 (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07624__S0 (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07534__S0 (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__S0 (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07354__S0 (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07261__S0 (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07080__S0 (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06981__S0 (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06880__S0 (.DIODE(_02826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06896__B1 (.DIODE(_02834_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07815__S1 (.DIODE(_02837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07724__S1 (.DIODE(_02837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07634__S1 (.DIODE(_02837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07544__S1 (.DIODE(_02837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07454__S1 (.DIODE(_02837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07364__S1 (.DIODE(_02837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07271__S1 (.DIODE(_02837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07091__S1 (.DIODE(_02837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06993__S1 (.DIODE(_02837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06891__S1 (.DIODE(_02837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06895__A2 (.DIODE(_02841_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06896__B2 (.DIODE(_02842_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06946__A2 (.DIODE(_02857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06924__B1 (.DIODE(_02867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__B (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08023__B (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07845__B (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07664__B (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07574__B (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07484__B (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07394__B (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07122__B (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07025__B (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06922__B (.DIODE(_02868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06925__D (.DIODE(_02871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06946__A3 (.DIODE(_02872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06934__B (.DIODE(_02875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06933__A2 (.DIODE(_02876_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08121__S1 (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08031__S1 (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07853__S1 (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07672__S1 (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__S1 (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07492__S1 (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07402__S1 (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07130__S1 (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07033__S1 (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06931__S1 (.DIODE(_02877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06946__B1 (.DIODE(_02881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06944__B1 (.DIODE(_02883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08131__B2 (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08040__B2 (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07862__B2 (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07681__B2 (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07591__B2 (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07501__B2 (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07411__B2 (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07139__B2 (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07043__B2 (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06944__B2 (.DIODE(_02884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08130__A1 (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08039__A1 (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07861__A1 (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07680__A1 (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07590__A1 (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07500__A1 (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__A1 (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07138__A1 (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07042__A1 (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06943__A1 (.DIODE(_02885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08129__S0 (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08038__S0 (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07860__S0 (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07679__S0 (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07589__S0 (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07499__S0 (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07409__S0 (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07137__S0 (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07041__S0 (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06941__S0 (.DIODE(_02887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08130__B2 (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08039__B2 (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07861__B2 (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07680__B2 (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07590__B2 (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07500__B2 (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__B2 (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07138__B2 (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07042__B2 (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06943__B2 (.DIODE(_02889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06944__C1 (.DIODE(_02890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06946__B2 (.DIODE(_02892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07960__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07782__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07691__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07601__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07511__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07421__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07238__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07055__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06955__A2 (.DIODE(_02899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06998__A2 (.DIODE(_02909_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06966__B1 (.DIODE(_02911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07973__B1 (.DIODE(_02914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__B1 (.DIODE(_02914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07704__B1 (.DIODE(_02914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07614__B1 (.DIODE(_02914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07524__B1 (.DIODE(_02914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07434__B1 (.DIODE(_02914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07344__B1 (.DIODE(_02914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07251__B1 (.DIODE(_02914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07070__B1 (.DIODE(_02914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06969__B1 (.DIODE(_02914_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07975__B (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07797__B (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07706__B (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07616__B (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07526__B (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07436__B (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07346__B (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07253__B (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07072__B (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06972__B (.DIODE(_02917_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06978__B2 (.DIODE(_02923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06979__D (.DIODE(_02924_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07983__S1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07805__S1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07714__S1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07624__S1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07534__S1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__S1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07354__S1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07261__S1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07080__S1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06981__S1 (.DIODE(_02926_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07984__S0 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07806__S0 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07715__S0 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07625__S0 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07535__S0 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07445__S0 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07355__S0 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07262__S0 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07081__S0 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06984__S0 (.DIODE(_02928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07984__S1 (.DIODE(_02929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07806__S1 (.DIODE(_02929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07715__S1 (.DIODE(_02929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07625__S1 (.DIODE(_02929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07535__S1 (.DIODE(_02929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07445__S1 (.DIODE(_02929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07355__S1 (.DIODE(_02929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07262__S1 (.DIODE(_02929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07081__S1 (.DIODE(_02929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06984__S1 (.DIODE(_02929_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06998__B1 (.DIODE(_02936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06997__A2 (.DIODE(_02942_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06998__B2 (.DIODE(_02943_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__A2 (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08011__A2 (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07833__A2 (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07652__A2 (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07562__A2 (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07472__A2 (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__A2 (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07295__A2 (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__A2 (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07013__A2 (.DIODE(_02955_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08100__A2 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08010__A2 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07832__A2 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07651__A2 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07561__A2 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07471__A2 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07381__A2 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07294__A2 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07109__A2 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07012__A2 (.DIODE(_02956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07045__A2 (.DIODE(_02960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07027__B1 (.DIODE(_02970_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07028__D (.DIODE(_02973_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07045__A3 (.DIODE(_02974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07036__B (.DIODE(_02977_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07035__A2 (.DIODE(_02978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07045__B1 (.DIODE(_02982_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08128__S0 (.DIODE(_02985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08037__S0 (.DIODE(_02985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07859__S0 (.DIODE(_02985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__S0 (.DIODE(_02985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07588__S0 (.DIODE(_02985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07498__S0 (.DIODE(_02985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07408__S0 (.DIODE(_02985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07303__A (.DIODE(_02985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07136__S0 (.DIODE(_02985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07040__S0 (.DIODE(_02985_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07045__B2 (.DIODE(_02990_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08058__A (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07968__A (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07790__A (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07699__A (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07609__A (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07519__A (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07429__A (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07339__A (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07246__A (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07063__A (.DIODE(_02993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08047__A2 (.DIODE(_02995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07957__A2 (.DIODE(_02995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07779__A2 (.DIODE(_02995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07688__A2 (.DIODE(_02995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07598__A2 (.DIODE(_02995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07508__A2 (.DIODE(_02995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07418__A2 (.DIODE(_02995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07328__A2 (.DIODE(_02995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__A2 (.DIODE(_02995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07052__A2 (.DIODE(_02995_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07096__A2 (.DIODE(_03008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08060__B1 (.DIODE(_03009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07970__B1 (.DIODE(_03009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07792__B1 (.DIODE(_03009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07701__B1 (.DIODE(_03009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__B1 (.DIODE(_03009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07521__B1 (.DIODE(_03009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07431__B1 (.DIODE(_03009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07341__B1 (.DIODE(_03009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07248__B1 (.DIODE(_03009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07066__B1 (.DIODE(_03009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07067__B1 (.DIODE(_03011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08062__B1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07972__B1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07794__B1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07703__B1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07613__B1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07523__B1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07433__B1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07343__B1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07250__B1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07069__B1 (.DIODE(_03013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07078__B2 (.DIODE(_03022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07079__D (.DIODE(_03023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07096__B1 (.DIODE(_03032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08086__A1 (.DIODE(_03033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07996__A1 (.DIODE(_03033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07818__A1 (.DIODE(_03033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07727__A1 (.DIODE(_03033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07637__A1 (.DIODE(_03033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__A1 (.DIODE(_03033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__A1 (.DIODE(_03033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07367__A1 (.DIODE(_03033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07274__A1 (.DIODE(_03033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07094__A1 (.DIODE(_03033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07095__A2 (.DIODE(_03039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07096__B2 (.DIODE(_03040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08089__A2 (.DIODE(_03042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__A2 (.DIODE(_03042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07821__A2 (.DIODE(_03042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07752__A2 (.DIODE(_03042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07640__A2 (.DIODE(_03042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07550__A2 (.DIODE(_03042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07460__A2 (.DIODE(_03042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07370__A2 (.DIODE(_03042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07301__A2 (.DIODE(_03042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07098__A2 (.DIODE(_03042_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07141__A2 (.DIODE(_03056_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__B1 (.DIODE(_03066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07125__D (.DIODE(_03069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07141__A3 (.DIODE(_03070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07133__B (.DIODE(_03073_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07141__B1 (.DIODE(_03078_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07141__B2 (.DIODE(_03085_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__B (.DIODE(_03092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09202__B (.DIODE(_03092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09061__B (.DIODE(_03092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08588__B (.DIODE(_03092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08553__B (.DIODE(_03092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08410__B (.DIODE(_03092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08336__B (.DIODE(_03092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08263__B (.DIODE(_03092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07872__B1 (.DIODE(_03092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__B1 (.DIODE(_03092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07188__A2 (.DIODE(_03102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__B1 (.DIODE(_03112_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07188__A3 (.DIODE(_03116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07179__B (.DIODE(_03122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07187__A2 (.DIODE(_03126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07216__A2 (.DIODE(_03146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07212__A2 (.DIODE(_03153_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07231__A2 (.DIODE(_03166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07232__B2 (.DIODE(_03175_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07276__A2 (.DIODE(_03189_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07259__B2 (.DIODE(_03201_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07260__D (.DIODE(_03202_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07276__B1 (.DIODE(_03211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07274__C1 (.DIODE(_03216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__A2 (.DIODE(_03217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07276__B2 (.DIODE(_03218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__B (.DIODE(_03224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08009__B (.DIODE(_03224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__B (.DIODE(_03224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07751__C_N (.DIODE(_03224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07744__B (.DIODE(_03224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07734__C_N (.DIODE(_03224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07650__B (.DIODE(_03224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07300__C_N (.DIODE(_03224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07293__B (.DIODE(_03224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07282__C_N (.DIODE(_03224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__B1 (.DIODE(_03231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08007__B1 (.DIODE(_03231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07829__B1 (.DIODE(_03231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07755__B1 (.DIODE(_03231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07741__B1 (.DIODE(_03231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07648__B1 (.DIODE(_03231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07558__B1 (.DIODE(_03231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07468__B1 (.DIODE(_03231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07304__B1 (.DIODE(_03231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07290__B1 (.DIODE(_03231_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07323__A2 (.DIODE(_03235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07323__A3 (.DIODE(_03249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07310__B (.DIODE(_03252_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__B1 (.DIODE(_03256_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07322__A2 (.DIODE(_03257_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07322__B1 (.DIODE(_03264_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07369__A2 (.DIODE(_03281_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07352__B2 (.DIODE(_03293_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07353__D (.DIODE(_03294_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07361__B (.DIODE(_03298_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07369__B1 (.DIODE(_03303_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07367__C1 (.DIODE(_03308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07368__A2 (.DIODE(_03309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07369__B2 (.DIODE(_03310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07413__A2 (.DIODE(_03325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07396__B1 (.DIODE(_03335_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07397__D (.DIODE(_03338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07413__A3 (.DIODE(_03339_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07405__B (.DIODE(_03342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07413__B1 (.DIODE(_03347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07412__A2 (.DIODE(_03353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07413__B2 (.DIODE(_03354_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07459__A2 (.DIODE(_03370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__B2 (.DIODE(_03382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07443__D (.DIODE(_03383_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07451__B (.DIODE(_03387_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07459__B1 (.DIODE(_03392_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__C1 (.DIODE(_03397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07458__A2 (.DIODE(_03398_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07459__B2 (.DIODE(_03399_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07503__A2 (.DIODE(_03414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07486__B1 (.DIODE(_03424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07487__D (.DIODE(_03427_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07503__A3 (.DIODE(_03428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07495__B (.DIODE(_03431_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07503__B1 (.DIODE(_03436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07503__B2 (.DIODE(_03443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07549__A2 (.DIODE(_03459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07532__B2 (.DIODE(_03471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07533__D (.DIODE(_03472_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07541__B (.DIODE(_03476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07549__B1 (.DIODE(_03481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07547__C1 (.DIODE(_03486_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07548__A2 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07549__B2 (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07593__A2 (.DIODE(_03503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07576__B1 (.DIODE(_03513_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07577__D (.DIODE(_03516_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07593__A3 (.DIODE(_03517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07585__B (.DIODE(_03520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07584__A2 (.DIODE(_03521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07593__B1 (.DIODE(_03525_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07592__A2 (.DIODE(_03531_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07609__D (.DIODE(_03547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07639__A2 (.DIODE(_03548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07622__A3 (.DIODE(_03557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07622__B2 (.DIODE(_03560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07623__D (.DIODE(_03561_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07639__B1 (.DIODE(_03570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07637__C1 (.DIODE(_03575_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07638__A2 (.DIODE(_03576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07639__B2 (.DIODE(_03577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07684__A0 (.DIODE(_03578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07653__D (.DIODE(_03591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__A2 (.DIODE(_03592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07667__D (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07675__B (.DIODE(_03609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__B1 (.DIODE(_03614_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07682__A2 (.DIODE(_03620_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__A2 (.DIODE(_03637_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__A3 (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07713__D (.DIODE(_03650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07721__B (.DIODE(_03654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__B1 (.DIODE(_03659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07727__C1 (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__A2 (.DIODE(_03665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__B2 (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07774__A2 (.DIODE(_03681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__A2 (.DIODE(_03703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07768__B1 (.DIODE(_03705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__B1 (.DIODE(_03708_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__B1 (.DIODE(_03710_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07790__C (.DIODE(_03723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07820__A2 (.DIODE(_03727_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07804__D (.DIODE(_03740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07820__B1 (.DIODE(_03749_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__A2 (.DIODE(_03755_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07820__B2 (.DIODE(_03756_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07864__A2 (.DIODE(_03771_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07848__D (.DIODE(_03784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07856__B (.DIODE(_03788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07855__A2 (.DIODE(_03789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07864__B1 (.DIODE(_03793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__A2 (.DIODE(_03799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__A2 (.DIODE(_03816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__A3 (.DIODE(_03830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__B (.DIODE(_03836_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07909__A2 (.DIODE(_03840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07938__A2 (.DIODE(_03860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07926__B (.DIODE(_03861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07934__A2 (.DIODE(_03867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07953__A2 (.DIODE(_03880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07954__B2 (.DIODE(_03889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07968__C (.DIODE(_03899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07998__A2 (.DIODE(_03903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07982__D (.DIODE(_03916_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07990__B (.DIODE(_03920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07998__B1 (.DIODE(_03925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07996__C1 (.DIODE(_03930_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07997__A2 (.DIODE(_03931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07998__B2 (.DIODE(_03932_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08012__D (.DIODE(_03946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08042__A2 (.DIODE(_03947_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08026__D (.DIODE(_03960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08034__B (.DIODE(_03964_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08042__B1 (.DIODE(_03969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08041__A2 (.DIODE(_03975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08058__C (.DIODE(_03988_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08088__A2 (.DIODE(_03992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08071__A3 (.DIODE(_04001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__D (.DIODE(_04005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08080__B (.DIODE(_04009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08088__B1 (.DIODE(_04014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08087__A2 (.DIODE(_04020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08088__B2 (.DIODE(_04021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08102__D (.DIODE(_04035_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08133__A2 (.DIODE(_04036_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__D (.DIODE(_04049_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__B (.DIODE(_04053_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08133__B1 (.DIODE(_04058_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10420__A (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09920__A (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09851__A (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09339__A (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08662__A (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08588__A (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08517__A (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08445__A (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08336__A (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08131__A1 (.DIODE(_04059_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08131__C1 (.DIODE(_04064_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08132__A2 (.DIODE(_04065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12104__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11535__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11139__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10915__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10592__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10126__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09731__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08697__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08208__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08137__A (.DIODE(_04069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12746__A0 (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12712__A0 (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12677__A0 (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08821__A1 (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08787__A1 (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08751__A1 (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08630__A1 (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08377__A1 (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__A1 (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08146__A1 (.DIODE(_04070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12293__A (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11724__A (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11140__A (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10558__A (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09425__A (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08921__A (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08819__A (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__A (.DIODE(_04072_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10489__C (.DIODE(_04075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10420__C (.DIODE(_04075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10385__A (.DIODE(_04075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10316__A (.DIODE(_04075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10212__C (.DIODE(_04075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08263__C (.DIODE(_04075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08143__A (.DIODE(_04075_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10455__A_N (.DIODE(_04076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10281__A (.DIODE(_04076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10247__A (.DIODE(_04076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10177__A (.DIODE(_04076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__A (.DIODE(_04076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10092__A (.DIODE(_04076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__A (.DIODE(_04076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10023__A (.DIODE(_04076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__A (.DIODE(_04076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__B (.DIODE(_04076_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12110__A (.DIODE(_04080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11541__A (.DIODE(_04080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11144__A (.DIODE(_04080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10921__A (.DIODE(_04080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10597__A (.DIODE(_04080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10132__A (.DIODE(_04080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09736__A (.DIODE(_04080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08704__A (.DIODE(_04080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08218__A (.DIODE(_04080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08149__A (.DIODE(_04080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12748__A0 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12714__A0 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12679__A0 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__A1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08789__A1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08753__A1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__A1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08379__A1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08306__A1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08150__A1 (.DIODE(_04081_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12113__A (.DIODE(_04083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11544__A (.DIODE(_04083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11147__A (.DIODE(_04083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10924__A (.DIODE(_04083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10600__A (.DIODE(_04083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10135__A (.DIODE(_04083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09739__A (.DIODE(_04083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08707__A (.DIODE(_04083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__A (.DIODE(_04083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08153__A (.DIODE(_04083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12750__A0 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12716__A0 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12681__A0 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__A1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08791__A1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08755__A1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08634__A1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__A1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08308__A1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08154__A1 (.DIODE(_04084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12116__A (.DIODE(_04086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11547__A (.DIODE(_04086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11150__A (.DIODE(_04086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__A (.DIODE(_04086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10603__A (.DIODE(_04086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10138__A (.DIODE(_04086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09742__A (.DIODE(_04086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08710__A (.DIODE(_04086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08224__A (.DIODE(_04086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08157__A (.DIODE(_04086_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12752__A0 (.DIODE(_04087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12718__A0 (.DIODE(_04087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12683__A0 (.DIODE(_04087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08827__A1 (.DIODE(_04087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08793__A1 (.DIODE(_04087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__A1 (.DIODE(_04087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08636__A1 (.DIODE(_04087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08383__A1 (.DIODE(_04087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08310__A1 (.DIODE(_04087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08158__A1 (.DIODE(_04087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12119__A (.DIODE(_04089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11550__A (.DIODE(_04089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11153__A (.DIODE(_04089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10930__A (.DIODE(_04089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10606__A (.DIODE(_04089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10141__A (.DIODE(_04089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09745__A (.DIODE(_04089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08713__A (.DIODE(_04089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08227__A (.DIODE(_04089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08161__A (.DIODE(_04089_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12754__A0 (.DIODE(_04090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12720__A0 (.DIODE(_04090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12685__A0 (.DIODE(_04090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08829__A1 (.DIODE(_04090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08795__A1 (.DIODE(_04090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08759__A1 (.DIODE(_04090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08638__A1 (.DIODE(_04090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08385__A1 (.DIODE(_04090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08312__A1 (.DIODE(_04090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08162__A1 (.DIODE(_04090_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12122__A (.DIODE(_04092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11553__A (.DIODE(_04092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__A (.DIODE(_04092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10933__A (.DIODE(_04092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10609__A (.DIODE(_04092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__A (.DIODE(_04092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09748__A (.DIODE(_04092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08716__A (.DIODE(_04092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08230__A (.DIODE(_04092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08165__A (.DIODE(_04092_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12756__A0 (.DIODE(_04093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12722__A0 (.DIODE(_04093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12687__A0 (.DIODE(_04093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08831__A1 (.DIODE(_04093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08797__A1 (.DIODE(_04093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08761__A1 (.DIODE(_04093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08640__A1 (.DIODE(_04093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__A1 (.DIODE(_04093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08314__A1 (.DIODE(_04093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08166__A1 (.DIODE(_04093_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12125__A (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11556__A (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11159__A (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__A (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10612__A (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10147__A (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09751__A (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08719__A (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__A (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08169__A (.DIODE(_04095_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12758__A0 (.DIODE(_04096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12724__A0 (.DIODE(_04096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12689__A0 (.DIODE(_04096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08833__A1 (.DIODE(_04096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08799__A1 (.DIODE(_04096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08763__A1 (.DIODE(_04096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08642__A1 (.DIODE(_04096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__A1 (.DIODE(_04096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08316__A1 (.DIODE(_04096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08170__A1 (.DIODE(_04096_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12128__A (.DIODE(_04098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11559__A (.DIODE(_04098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11162__A (.DIODE(_04098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10939__A (.DIODE(_04098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10615__A (.DIODE(_04098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__A (.DIODE(_04098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09754__A (.DIODE(_04098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08722__A (.DIODE(_04098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__A (.DIODE(_04098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__A (.DIODE(_04098_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12760__A0 (.DIODE(_04099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12726__A0 (.DIODE(_04099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12691__A0 (.DIODE(_04099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08835__A1 (.DIODE(_04099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08801__A1 (.DIODE(_04099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08765__A1 (.DIODE(_04099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08644__A1 (.DIODE(_04099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08391__A1 (.DIODE(_04099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__A1 (.DIODE(_04099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08174__A1 (.DIODE(_04099_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12131__A (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11562__A (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11165__A (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10942__A (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10618__A (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10153__A (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09757__A (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08725__A (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08239__A (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08177__A (.DIODE(_04101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12762__A0 (.DIODE(_04102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12728__A0 (.DIODE(_04102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12693__A0 (.DIODE(_04102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08837__A1 (.DIODE(_04102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08803__A1 (.DIODE(_04102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__A1 (.DIODE(_04102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08646__A1 (.DIODE(_04102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__A1 (.DIODE(_04102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08320__A1 (.DIODE(_04102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08178__A1 (.DIODE(_04102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12134__A (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11565__A (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11168__A (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10945__A (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10621__A (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__A (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09760__A (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08728__A (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08242__A (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08181__A (.DIODE(_04104_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12764__A0 (.DIODE(_04105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12730__A0 (.DIODE(_04105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12695__A0 (.DIODE(_04105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08839__A1 (.DIODE(_04105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08805__A1 (.DIODE(_04105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08769__A1 (.DIODE(_04105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08648__A1 (.DIODE(_04105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08395__A1 (.DIODE(_04105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08322__A1 (.DIODE(_04105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__A1 (.DIODE(_04105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12137__A (.DIODE(_04107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11568__A (.DIODE(_04107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__A (.DIODE(_04107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10948__A (.DIODE(_04107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10624__A (.DIODE(_04107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10159__A (.DIODE(_04107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09763__A (.DIODE(_04107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08731__A (.DIODE(_04107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08245__A (.DIODE(_04107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08185__A (.DIODE(_04107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12766__A0 (.DIODE(_04108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12732__A0 (.DIODE(_04108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12697__A0 (.DIODE(_04108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__A1 (.DIODE(_04108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08807__A1 (.DIODE(_04108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08771__A1 (.DIODE(_04108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08650__A1 (.DIODE(_04108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08397__A1 (.DIODE(_04108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08324__A1 (.DIODE(_04108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08186__A1 (.DIODE(_04108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12140__A (.DIODE(_04110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11571__A (.DIODE(_04110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__A (.DIODE(_04110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__A (.DIODE(_04110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10627__A (.DIODE(_04110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10162__A (.DIODE(_04110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09766__A (.DIODE(_04110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08734__A (.DIODE(_04110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08248__A (.DIODE(_04110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08189__A (.DIODE(_04110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12768__A0 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12734__A0 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12699__A0 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08843__A1 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08809__A1 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08773__A1 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08652__A1 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__A1 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__A1 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08190__A1 (.DIODE(_04111_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__A (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11574__A (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11177__A (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10954__A (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10630__A (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10165__A (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__A (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08737__A (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08251__A (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08193__A (.DIODE(_04113_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12770__A0 (.DIODE(_04114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12736__A0 (.DIODE(_04114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12701__A0 (.DIODE(_04114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__A1 (.DIODE(_04114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08811__A1 (.DIODE(_04114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08775__A1 (.DIODE(_04114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08654__A1 (.DIODE(_04114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08401__A1 (.DIODE(_04114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08328__A1 (.DIODE(_04114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__A1 (.DIODE(_04114_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12146__A (.DIODE(_04116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11577__A (.DIODE(_04116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11180__A (.DIODE(_04116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10957__A (.DIODE(_04116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10633__A (.DIODE(_04116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10168__A (.DIODE(_04116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09772__A (.DIODE(_04116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08740__A (.DIODE(_04116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08254__A (.DIODE(_04116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08197__A (.DIODE(_04116_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12772__A0 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12738__A0 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12703__A0 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08847__A1 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08813__A1 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08777__A1 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08656__A1 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__A1 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08330__A1 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08198__A1 (.DIODE(_04117_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12149__A (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11580__A (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11183__A (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10960__A (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10636__A (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10171__A (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09775__A (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08743__A (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08257__A (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08201__A (.DIODE(_04119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12774__A0 (.DIODE(_04120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12740__A0 (.DIODE(_04120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12705__A0 (.DIODE(_04120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08849__A1 (.DIODE(_04120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08815__A1 (.DIODE(_04120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08779__A1 (.DIODE(_04120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08658__A1 (.DIODE(_04120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08405__A1 (.DIODE(_04120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08332__A1 (.DIODE(_04120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08202__A1 (.DIODE(_04120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12152__A (.DIODE(_04122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11583__A (.DIODE(_04122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__A (.DIODE(_04122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10963__A (.DIODE(_04122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10639__A (.DIODE(_04122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10174__A (.DIODE(_04122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09778__A (.DIODE(_04122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08746__A (.DIODE(_04122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08260__A (.DIODE(_04122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08205__A (.DIODE(_04122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12776__A0 (.DIODE(_04123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12742__A0 (.DIODE(_04123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12707__A0 (.DIODE(_04123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08851__A1 (.DIODE(_04123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08817__A1 (.DIODE(_04123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08781__A1 (.DIODE(_04123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08660__A1 (.DIODE(_04123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08407__A1 (.DIODE(_04123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08334__A1 (.DIODE(_04123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08206__A1 (.DIODE(_04123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08665__A0 (.DIODE(_04125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08591__A0 (.DIODE(_04125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08556__A0 (.DIODE(_04125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08520__A0 (.DIODE(_04125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08485__A0 (.DIODE(_04125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__A0 (.DIODE(_04125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08413__A0 (.DIODE(_04125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08339__A0 (.DIODE(_04125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08266__A0 (.DIODE(_04125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08216__A0 (.DIODE(_04125_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12778__A (.DIODE(_04127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12569__A (.DIODE(_04127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11999__A (.DIODE(_04127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10847__A (.DIODE(_04127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10281__B (.DIODE(_04127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09697__A (.DIODE(_04127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09132__A (.DIODE(_04127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08213__A (.DIODE(_04127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08261__S (.DIODE(_04131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08258__S (.DIODE(_04131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08255__S (.DIODE(_04131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08252__S (.DIODE(_04131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08249__S (.DIODE(_04131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08246__S (.DIODE(_04131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08215__A (.DIODE(_04131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08243__S (.DIODE(_04132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08240__S (.DIODE(_04132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08237__S (.DIODE(_04132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08234__S (.DIODE(_04132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__S (.DIODE(_04132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08228__S (.DIODE(_04132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08225__S (.DIODE(_04132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08222__S (.DIODE(_04132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08219__S (.DIODE(_04132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08216__S (.DIODE(_04132_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08667__A0 (.DIODE(_04134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__A0 (.DIODE(_04134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08558__A0 (.DIODE(_04134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__A0 (.DIODE(_04134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08487__A0 (.DIODE(_04134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08450__A0 (.DIODE(_04134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08415__A0 (.DIODE(_04134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__A0 (.DIODE(_04134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08268__A0 (.DIODE(_04134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08219__A0 (.DIODE(_04134_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08669__A0 (.DIODE(_04136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__A0 (.DIODE(_04136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08560__A0 (.DIODE(_04136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08524__A0 (.DIODE(_04136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08489__A0 (.DIODE(_04136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08452__A0 (.DIODE(_04136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08417__A0 (.DIODE(_04136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08343__A0 (.DIODE(_04136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08270__A0 (.DIODE(_04136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08222__A0 (.DIODE(_04136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08671__A0 (.DIODE(_04138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08597__A0 (.DIODE(_04138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08562__A0 (.DIODE(_04138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08526__A0 (.DIODE(_04138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08491__A0 (.DIODE(_04138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08454__A0 (.DIODE(_04138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08419__A0 (.DIODE(_04138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08345__A0 (.DIODE(_04138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08272__A0 (.DIODE(_04138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08225__A0 (.DIODE(_04138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08673__A0 (.DIODE(_04140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__A0 (.DIODE(_04140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08564__A0 (.DIODE(_04140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08528__A0 (.DIODE(_04140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08493__A0 (.DIODE(_04140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08456__A0 (.DIODE(_04140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08421__A0 (.DIODE(_04140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08347__A0 (.DIODE(_04140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08274__A0 (.DIODE(_04140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08228__A0 (.DIODE(_04140_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08675__A0 (.DIODE(_04142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08601__A0 (.DIODE(_04142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08566__A0 (.DIODE(_04142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__A0 (.DIODE(_04142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08495__A0 (.DIODE(_04142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08458__A0 (.DIODE(_04142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08423__A0 (.DIODE(_04142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08349__A0 (.DIODE(_04142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08276__A0 (.DIODE(_04142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__A0 (.DIODE(_04142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08677__A0 (.DIODE(_04144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08603__A0 (.DIODE(_04144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08568__A0 (.DIODE(_04144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__A0 (.DIODE(_04144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08497__A0 (.DIODE(_04144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08460__A0 (.DIODE(_04144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08425__A0 (.DIODE(_04144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08351__A0 (.DIODE(_04144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08278__A0 (.DIODE(_04144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08234__A0 (.DIODE(_04144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08679__A0 (.DIODE(_04146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08605__A0 (.DIODE(_04146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08570__A0 (.DIODE(_04146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08534__A0 (.DIODE(_04146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08499__A0 (.DIODE(_04146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08462__A0 (.DIODE(_04146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08427__A0 (.DIODE(_04146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08353__A0 (.DIODE(_04146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08280__A0 (.DIODE(_04146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08237__A0 (.DIODE(_04146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08681__A0 (.DIODE(_04148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08607__A0 (.DIODE(_04148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__A0 (.DIODE(_04148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08536__A0 (.DIODE(_04148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08501__A0 (.DIODE(_04148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08464__A0 (.DIODE(_04148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08429__A0 (.DIODE(_04148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08355__A0 (.DIODE(_04148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08282__A0 (.DIODE(_04148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08240__A0 (.DIODE(_04148_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08683__A0 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08609__A0 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08574__A0 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08538__A0 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08503__A0 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08466__A0 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08431__A0 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__A0 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08284__A0 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08243__A0 (.DIODE(_04150_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08685__A0 (.DIODE(_04152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08611__A0 (.DIODE(_04152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08576__A0 (.DIODE(_04152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__A0 (.DIODE(_04152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08505__A0 (.DIODE(_04152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08468__A0 (.DIODE(_04152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08433__A0 (.DIODE(_04152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08359__A0 (.DIODE(_04152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08286__A0 (.DIODE(_04152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08246__A0 (.DIODE(_04152_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08687__A0 (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08613__A0 (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__A0 (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08542__A0 (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08507__A0 (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08470__A0 (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08435__A0 (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08361__A0 (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08288__A0 (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08249__A0 (.DIODE(_04154_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08689__A0 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08615__A0 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08580__A0 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08544__A0 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08509__A0 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08472__A0 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08437__A0 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08363__A0 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08290__A0 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08252__A0 (.DIODE(_04156_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08691__A0 (.DIODE(_04158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08617__A0 (.DIODE(_04158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08582__A0 (.DIODE(_04158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08546__A0 (.DIODE(_04158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08511__A0 (.DIODE(_04158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08474__A0 (.DIODE(_04158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08439__A0 (.DIODE(_04158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08365__A0 (.DIODE(_04158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08292__A0 (.DIODE(_04158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08255__A0 (.DIODE(_04158_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08693__A0 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08619__A0 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08584__A0 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08548__A0 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08513__A0 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__A0 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08441__A0 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08367__A0 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08294__A0 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08258__A0 (.DIODE(_04160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08695__A0 (.DIODE(_04162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08621__A0 (.DIODE(_04162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__A0 (.DIODE(_04162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08550__A0 (.DIODE(_04162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08515__A0 (.DIODE(_04162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__A0 (.DIODE(_04162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08443__A0 (.DIODE(_04162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08369__A0 (.DIODE(_04162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08296__A0 (.DIODE(_04162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08261__A0 (.DIODE(_04162_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08284__S (.DIODE(_04166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08282__S (.DIODE(_04166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08280__S (.DIODE(_04166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08278__S (.DIODE(_04166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08276__S (.DIODE(_04166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08274__S (.DIODE(_04166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08272__S (.DIODE(_04166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08270__S (.DIODE(_04166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08268__S (.DIODE(_04166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08266__S (.DIODE(_04166_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12430__A (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11860__A (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11292__B (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10351__A (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__B (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09561__A (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08991__A (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__A (.DIODE(_04184_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11035__A_N (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11000__C (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10966__A (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10916__C (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10778__C (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08336__C (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08301__A (.DIODE(_04185_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08334__S (.DIODE(_04187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08332__S (.DIODE(_04187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08330__S (.DIODE(_04187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08328__S (.DIODE(_04187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__S (.DIODE(_04187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08324__S (.DIODE(_04187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08303__A (.DIODE(_04187_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08322__S (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08320__S (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__S (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08316__S (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08314__S (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08312__S (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08310__S (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08308__S (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08306__S (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__S (.DIODE(_04188_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12361__A (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11223__B (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10642__B (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10057__B (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09629__A (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09493__A (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08482__A (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__A (.DIODE(_04225_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08407__S (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08405__S (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__S (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08401__S (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__S (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08397__S (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08376__A (.DIODE(_04228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08395__S (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__S (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08391__S (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__S (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__S (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08385__S (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08383__S (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__S (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08379__S (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08377__S (.DIODE(_04229_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09920__C (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09886__A_N (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09851__C (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__A (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09782__C (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09375__A (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08410__C (.DIODE(_04246_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08443__S (.DIODE(_04248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08441__S (.DIODE(_04248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08439__S (.DIODE(_04248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08437__S (.DIODE(_04248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08435__S (.DIODE(_04248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08433__S (.DIODE(_04248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08412__A (.DIODE(_04248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08431__S (.DIODE(_04249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08429__S (.DIODE(_04249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08427__S (.DIODE(_04249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08425__S (.DIODE(_04249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08423__S (.DIODE(_04249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08421__S (.DIODE(_04249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08419__S (.DIODE(_04249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08417__S (.DIODE(_04249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08415__S (.DIODE(_04249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08413__S (.DIODE(_04249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__S (.DIODE(_04267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__S (.DIODE(_04267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08474__S (.DIODE(_04267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08472__S (.DIODE(_04267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08470__S (.DIODE(_04267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08468__S (.DIODE(_04267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08447__A (.DIODE(_04267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08466__S (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08464__S (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08462__S (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08460__S (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08458__S (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08456__S (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08454__S (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08452__S (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08450__S (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08448__S (.DIODE(_04268_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12223__C (.DIODE(_04285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12069__C (.DIODE(_04285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11999__B (.DIODE(_04285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11930__C (.DIODE(_04285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11860__B (.DIODE(_04285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08517__C (.DIODE(_04285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08481__A (.DIODE(_04285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12189__A_N (.DIODE(_04286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12105__A (.DIODE(_04286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12034__A (.DIODE(_04286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11965__A (.DIODE(_04286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11895__A (.DIODE(_04286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11826__A (.DIODE(_04286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11758__A (.DIODE(_04286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11724__B (.DIODE(_04286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11690__A (.DIODE(_04286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08482__B (.DIODE(_04286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08515__S (.DIODE(_04288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08513__S (.DIODE(_04288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08511__S (.DIODE(_04288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08509__S (.DIODE(_04288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08507__S (.DIODE(_04288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08505__S (.DIODE(_04288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08484__A (.DIODE(_04288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08503__S (.DIODE(_04289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08501__S (.DIODE(_04289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08499__S (.DIODE(_04289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08497__S (.DIODE(_04289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08495__S (.DIODE(_04289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08493__S (.DIODE(_04289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08491__S (.DIODE(_04289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08489__S (.DIODE(_04289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08487__S (.DIODE(_04289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08485__S (.DIODE(_04289_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08550__S (.DIODE(_04307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08548__S (.DIODE(_04307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08546__S (.DIODE(_04307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08544__S (.DIODE(_04307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08542__S (.DIODE(_04307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08540__S (.DIODE(_04307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08519__A (.DIODE(_04307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08538__S (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08536__S (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08534__S (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08532__S (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__S (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08528__S (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08526__S (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08524__S (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__S (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08520__S (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12709__C (.DIODE(_04325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12639__C (.DIODE(_04325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12569__B (.DIODE(_04325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12430__B (.DIODE(_04325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12258__A (.DIODE(_04325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08588__C (.DIODE(_04325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08553__C (.DIODE(_04325_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__S (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08584__S (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08582__S (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08580__S (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08578__S (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08576__S (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08555__A (.DIODE(_04327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08574__S (.DIODE(_04328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08572__S (.DIODE(_04328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08570__S (.DIODE(_04328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08568__S (.DIODE(_04328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08566__S (.DIODE(_04328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08564__S (.DIODE(_04328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08562__S (.DIODE(_04328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08560__S (.DIODE(_04328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08558__S (.DIODE(_04328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08556__S (.DIODE(_04328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08621__S (.DIODE(_04346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08619__S (.DIODE(_04346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08617__S (.DIODE(_04346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08615__S (.DIODE(_04346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08613__S (.DIODE(_04346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08611__S (.DIODE(_04346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08590__A (.DIODE(_04346_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08609__S (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08607__S (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08605__S (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08603__S (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08601__S (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08599__S (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08597__S (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__S (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__S (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08591__S (.DIODE(_04347_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12674__B (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12105__B (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11536__B (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10966__B (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10385__B (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__B (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09237__B (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08628__A (.DIODE(_04365_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12500__C (.DIODE(_04367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12155__A (.DIODE(_04367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11069__C (.DIODE(_04367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08749__C (.DIODE(_04367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08700__A_N (.DIODE(_04367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08662__C (.DIODE(_04367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08627__A (.DIODE(_04367_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12778__B (.DIODE(_04368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11792__A (.DIODE(_04368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11431__A (.DIODE(_04368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10710__A (.DIODE(_04368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10351__B (.DIODE(_04368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09989__A (.DIODE(_04368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09629__B (.DIODE(_04368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__A (.DIODE(_04368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08921__B (.DIODE(_04368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08628__B (.DIODE(_04368_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08648__S (.DIODE(_04370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08646__S (.DIODE(_04370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08644__S (.DIODE(_04370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08642__S (.DIODE(_04370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08640__S (.DIODE(_04370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08638__S (.DIODE(_04370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08636__S (.DIODE(_04370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08634__S (.DIODE(_04370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__S (.DIODE(_04370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08630__S (.DIODE(_04370_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08695__S (.DIODE(_04388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08693__S (.DIODE(_04388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08691__S (.DIODE(_04388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08689__S (.DIODE(_04388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08687__S (.DIODE(_04388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08685__S (.DIODE(_04388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08664__A (.DIODE(_04388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08683__S (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08681__S (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08679__S (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08677__S (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08675__S (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08673__S (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08671__S (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08669__S (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08667__S (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08665__S (.DIODE(_04389_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10060__A0 (.DIODE(_04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09923__A0 (.DIODE(_04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09888__A0 (.DIODE(_04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09854__A0 (.DIODE(_04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09785__A0 (.DIODE(_04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09342__A0 (.DIODE(_04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09307__A0 (.DIODE(_04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09205__A0 (.DIODE(_04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09064__A0 (.DIODE(_04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08702__A0 (.DIODE(_04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12744__B (.DIODE(_04408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12189__B (.DIODE(_04408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11621__B (.DIODE(_04408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11035__B (.DIODE(_04408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10455__B (.DIODE(_04408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09886__B (.DIODE(_04408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09305__B (.DIODE(_04408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08700__B (.DIODE(_04408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08729__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08726__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08723__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08720__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08717__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08714__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08711__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08708__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08705__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08702__S (.DIODE(_04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10062__A0 (.DIODE(_04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09925__A0 (.DIODE(_04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09890__A0 (.DIODE(_04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09856__A0 (.DIODE(_04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09787__A0 (.DIODE(_04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09344__A0 (.DIODE(_04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09309__A0 (.DIODE(_04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09207__A0 (.DIODE(_04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09066__A0 (.DIODE(_04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08705__A0 (.DIODE(_04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10064__A0 (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09927__A0 (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09892__A0 (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09858__A0 (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09789__A0 (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09346__A0 (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09311__A0 (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09209__A0 (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09068__A0 (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08708__A0 (.DIODE(_04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10066__A0 (.DIODE(_04416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09929__A0 (.DIODE(_04416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09894__A0 (.DIODE(_04416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09860__A0 (.DIODE(_04416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09791__A0 (.DIODE(_04416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09348__A0 (.DIODE(_04416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__A0 (.DIODE(_04416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09211__A0 (.DIODE(_04416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__A0 (.DIODE(_04416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08711__A0 (.DIODE(_04416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10068__A0 (.DIODE(_04418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09931__A0 (.DIODE(_04418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09896__A0 (.DIODE(_04418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09862__A0 (.DIODE(_04418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09793__A0 (.DIODE(_04418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09350__A0 (.DIODE(_04418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__A0 (.DIODE(_04418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09213__A0 (.DIODE(_04418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__A0 (.DIODE(_04418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08714__A0 (.DIODE(_04418_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10070__A0 (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09933__A0 (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09898__A0 (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09864__A0 (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__A0 (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09352__A0 (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09317__A0 (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09215__A0 (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09074__A0 (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08717__A0 (.DIODE(_04420_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10072__A0 (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__A0 (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__A0 (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09866__A0 (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09797__A0 (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09354__A0 (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09319__A0 (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09217__A0 (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09076__A0 (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08720__A0 (.DIODE(_04422_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10074__A0 (.DIODE(_04424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09937__A0 (.DIODE(_04424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09902__A0 (.DIODE(_04424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09868__A0 (.DIODE(_04424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09799__A0 (.DIODE(_04424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09356__A0 (.DIODE(_04424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09321__A0 (.DIODE(_04424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09219__A0 (.DIODE(_04424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09078__A0 (.DIODE(_04424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08723__A0 (.DIODE(_04424_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10076__A0 (.DIODE(_04426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__A0 (.DIODE(_04426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09904__A0 (.DIODE(_04426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09870__A0 (.DIODE(_04426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__A0 (.DIODE(_04426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09358__A0 (.DIODE(_04426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09323__A0 (.DIODE(_04426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__A0 (.DIODE(_04426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__A0 (.DIODE(_04426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08726__A0 (.DIODE(_04426_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10078__A0 (.DIODE(_04428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__A0 (.DIODE(_04428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09906__A0 (.DIODE(_04428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__A0 (.DIODE(_04428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09803__A0 (.DIODE(_04428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__A0 (.DIODE(_04428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__A0 (.DIODE(_04428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09223__A0 (.DIODE(_04428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09082__A0 (.DIODE(_04428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08729__A0 (.DIODE(_04428_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10080__A0 (.DIODE(_04430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09943__A0 (.DIODE(_04430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09908__A0 (.DIODE(_04430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09874__A0 (.DIODE(_04430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__A0 (.DIODE(_04430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09362__A0 (.DIODE(_04430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09327__A0 (.DIODE(_04430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09225__A0 (.DIODE(_04430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09084__A0 (.DIODE(_04430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08732__A0 (.DIODE(_04430_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10082__A0 (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09945__A0 (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__A0 (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09876__A0 (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09807__A0 (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09364__A0 (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09329__A0 (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__A0 (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__A0 (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08735__A0 (.DIODE(_04432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10084__A0 (.DIODE(_04434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09947__A0 (.DIODE(_04434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09912__A0 (.DIODE(_04434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09878__A0 (.DIODE(_04434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09809__A0 (.DIODE(_04434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09366__A0 (.DIODE(_04434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09331__A0 (.DIODE(_04434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__A0 (.DIODE(_04434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09088__A0 (.DIODE(_04434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08738__A0 (.DIODE(_04434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10086__A0 (.DIODE(_04436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__A0 (.DIODE(_04436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09914__A0 (.DIODE(_04436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09880__A0 (.DIODE(_04436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09811__A0 (.DIODE(_04436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09368__A0 (.DIODE(_04436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09333__A0 (.DIODE(_04436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__A0 (.DIODE(_04436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09090__A0 (.DIODE(_04436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08741__A0 (.DIODE(_04436_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10088__A0 (.DIODE(_04438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__A0 (.DIODE(_04438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09916__A0 (.DIODE(_04438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09882__A0 (.DIODE(_04438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09813__A0 (.DIODE(_04438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__A0 (.DIODE(_04438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09335__A0 (.DIODE(_04438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__A0 (.DIODE(_04438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09092__A0 (.DIODE(_04438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08744__A0 (.DIODE(_04438_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10090__A0 (.DIODE(_04440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09953__A0 (.DIODE(_04440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09918__A0 (.DIODE(_04440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09884__A0 (.DIODE(_04440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09815__A0 (.DIODE(_04440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09372__A0 (.DIODE(_04440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09337__A0 (.DIODE(_04440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09235__A0 (.DIODE(_04440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09094__A0 (.DIODE(_04440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08747__A0 (.DIODE(_04440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08781__S (.DIODE(_04442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08779__S (.DIODE(_04442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08777__S (.DIODE(_04442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08775__S (.DIODE(_04442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08773__S (.DIODE(_04442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08771__S (.DIODE(_04442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08750__A (.DIODE(_04442_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08769__S (.DIODE(_04443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08767__S (.DIODE(_04443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08765__S (.DIODE(_04443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08763__S (.DIODE(_04443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08761__S (.DIODE(_04443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08759__S (.DIODE(_04443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__S (.DIODE(_04443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08755__S (.DIODE(_04443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08753__S (.DIODE(_04443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08751__S (.DIODE(_04443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12259__B (.DIODE(_04461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11792__B (.DIODE(_04461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11690__B (.DIODE(_04461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11105__B (.DIODE(_04461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10524__B (.DIODE(_04461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__B (.DIODE(_04461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__B (.DIODE(_04461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08785__B (.DIODE(_04461_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08817__S (.DIODE(_04462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08815__S (.DIODE(_04462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08813__S (.DIODE(_04462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08811__S (.DIODE(_04462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08809__S (.DIODE(_04462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08807__S (.DIODE(_04462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08786__A (.DIODE(_04462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08805__S (.DIODE(_04463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08803__S (.DIODE(_04463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08801__S (.DIODE(_04463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08799__S (.DIODE(_04463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08797__S (.DIODE(_04463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08795__S (.DIODE(_04463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08793__S (.DIODE(_04463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08791__S (.DIODE(_04463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08789__S (.DIODE(_04463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08787__S (.DIODE(_04463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08851__S (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08849__S (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08847__S (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__S (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08843__S (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08841__S (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08820__A (.DIODE(_04480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08839__S (.DIODE(_04481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08837__S (.DIODE(_04481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08835__S (.DIODE(_04481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08833__S (.DIODE(_04481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08831__S (.DIODE(_04481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08829__S (.DIODE(_04481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08827__S (.DIODE(_04481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08825__S (.DIODE(_04481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08823__S (.DIODE(_04481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08821__S (.DIODE(_04481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12780__A1 (.DIODE(_04498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12537__A1 (.DIODE(_04498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12398__A1 (.DIODE(_04498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12329__A1 (.DIODE(_04498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12295__A1 (.DIODE(_04498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12261__A1 (.DIODE(_04498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12157__A1 (.DIODE(_04498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11967__A1 (.DIODE(_04498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09374__A (.DIODE(_04498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08854__A (.DIODE(_04498_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09273__A1 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09239__A1 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09170__A1 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09134__A1 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09100__A1 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09029__A1 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08993__A1 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08959__A1 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08923__A1 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08859__A1 (.DIODE(_04499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12327__B (.DIODE(_04501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11758__B (.DIODE(_04501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11189__B (.DIODE(_04501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10593__B (.DIODE(_04501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10023__B (.DIODE(_04501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09459__B (.DIODE(_04501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__B (.DIODE(_04501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08857__B (.DIODE(_04501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08919__S (.DIODE(_04502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08915__S (.DIODE(_04502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08911__S (.DIODE(_04502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__S (.DIODE(_04502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08903__S (.DIODE(_04502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08899__S (.DIODE(_04502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08858__A (.DIODE(_04502_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08895__S (.DIODE(_04503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08891__S (.DIODE(_04503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08887__S (.DIODE(_04503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08883__S (.DIODE(_04503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08879__S (.DIODE(_04503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08875__S (.DIODE(_04503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08871__S (.DIODE(_04503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08867__S (.DIODE(_04503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08863__S (.DIODE(_04503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08859__S (.DIODE(_04503_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12782__A1 (.DIODE(_04505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12539__A1 (.DIODE(_04505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12400__A1 (.DIODE(_04505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12331__A1 (.DIODE(_04505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12297__A1 (.DIODE(_04505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12263__A1 (.DIODE(_04505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12159__A1 (.DIODE(_04505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11969__A1 (.DIODE(_04505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__A (.DIODE(_04505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08862__A (.DIODE(_04505_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09275__A1 (.DIODE(_04506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09241__A1 (.DIODE(_04506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__A1 (.DIODE(_04506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09136__A1 (.DIODE(_04506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09102__A1 (.DIODE(_04506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09031__A1 (.DIODE(_04506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08995__A1 (.DIODE(_04506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08961__A1 (.DIODE(_04506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08925__A1 (.DIODE(_04506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08863__A1 (.DIODE(_04506_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12784__A1 (.DIODE(_04508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12541__A1 (.DIODE(_04508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12402__A1 (.DIODE(_04508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12333__A1 (.DIODE(_04508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__A1 (.DIODE(_04508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12265__A1 (.DIODE(_04508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12161__A1 (.DIODE(_04508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11971__A1 (.DIODE(_04508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09383__A (.DIODE(_04508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08866__A (.DIODE(_04508_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09277__A1 (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09243__A1 (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09174__A1 (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09138__A1 (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09104__A1 (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09033__A1 (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08997__A1 (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08963__A1 (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08927__A1 (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08867__A1 (.DIODE(_04509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12786__A1 (.DIODE(_04511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12543__A1 (.DIODE(_04511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12404__A1 (.DIODE(_04511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12335__A1 (.DIODE(_04511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12301__A1 (.DIODE(_04511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12267__A1 (.DIODE(_04511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12163__A1 (.DIODE(_04511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11973__A1 (.DIODE(_04511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09386__A (.DIODE(_04511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08870__A (.DIODE(_04511_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09279__A1 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09245__A1 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09176__A1 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09140__A1 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09106__A1 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09035__A1 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08999__A1 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08965__A1 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08929__A1 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08871__A1 (.DIODE(_04512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12788__A1 (.DIODE(_04514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12545__A1 (.DIODE(_04514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12406__A1 (.DIODE(_04514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12337__A1 (.DIODE(_04514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12303__A1 (.DIODE(_04514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12269__A1 (.DIODE(_04514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12165__A1 (.DIODE(_04514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11975__A1 (.DIODE(_04514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09389__A (.DIODE(_04514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08874__A (.DIODE(_04514_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__A1 (.DIODE(_04515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09247__A1 (.DIODE(_04515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09178__A1 (.DIODE(_04515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09142__A1 (.DIODE(_04515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09108__A1 (.DIODE(_04515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09037__A1 (.DIODE(_04515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09001__A1 (.DIODE(_04515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08967__A1 (.DIODE(_04515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08931__A1 (.DIODE(_04515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08875__A1 (.DIODE(_04515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12790__A1 (.DIODE(_04517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12547__A1 (.DIODE(_04517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12408__A1 (.DIODE(_04517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12339__A1 (.DIODE(_04517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12305__A1 (.DIODE(_04517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12271__A1 (.DIODE(_04517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12167__A1 (.DIODE(_04517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11977__A1 (.DIODE(_04517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09392__A (.DIODE(_04517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08878__A (.DIODE(_04517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__A1 (.DIODE(_04518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09249__A1 (.DIODE(_04518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09180__A1 (.DIODE(_04518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09144__A1 (.DIODE(_04518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09110__A1 (.DIODE(_04518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09039__A1 (.DIODE(_04518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09003__A1 (.DIODE(_04518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08969__A1 (.DIODE(_04518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08933__A1 (.DIODE(_04518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08879__A1 (.DIODE(_04518_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12792__A1 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12549__A1 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12410__A1 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12341__A1 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12307__A1 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12273__A1 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12169__A1 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11979__A1 (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09395__A (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08882__A (.DIODE(_04520_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09285__A1 (.DIODE(_04521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09251__A1 (.DIODE(_04521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09182__A1 (.DIODE(_04521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09146__A1 (.DIODE(_04521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09112__A1 (.DIODE(_04521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09041__A1 (.DIODE(_04521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09005__A1 (.DIODE(_04521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08971__A1 (.DIODE(_04521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08935__A1 (.DIODE(_04521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08883__A1 (.DIODE(_04521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12794__A1 (.DIODE(_04523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12551__A1 (.DIODE(_04523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12412__A1 (.DIODE(_04523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12343__A1 (.DIODE(_04523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__A1 (.DIODE(_04523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12275__A1 (.DIODE(_04523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12171__A1 (.DIODE(_04523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11981__A1 (.DIODE(_04523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09398__A (.DIODE(_04523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08886__A (.DIODE(_04523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09287__A1 (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__A1 (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09184__A1 (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09148__A1 (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09114__A1 (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09043__A1 (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09007__A1 (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08973__A1 (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08937__A1 (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08887__A1 (.DIODE(_04524_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12796__A1 (.DIODE(_04526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12553__A1 (.DIODE(_04526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12414__A1 (.DIODE(_04526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12345__A1 (.DIODE(_04526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12311__A1 (.DIODE(_04526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12277__A1 (.DIODE(_04526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12173__A1 (.DIODE(_04526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11983__A1 (.DIODE(_04526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09401__A (.DIODE(_04526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08890__A (.DIODE(_04526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__A1 (.DIODE(_04527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09255__A1 (.DIODE(_04527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09186__A1 (.DIODE(_04527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09150__A1 (.DIODE(_04527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09116__A1 (.DIODE(_04527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09045__A1 (.DIODE(_04527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09009__A1 (.DIODE(_04527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08975__A1 (.DIODE(_04527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08939__A1 (.DIODE(_04527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08891__A1 (.DIODE(_04527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12798__A1 (.DIODE(_04529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12555__A1 (.DIODE(_04529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12416__A1 (.DIODE(_04529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12347__A1 (.DIODE(_04529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12313__A1 (.DIODE(_04529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12279__A1 (.DIODE(_04529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12175__A1 (.DIODE(_04529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11985__A1 (.DIODE(_04529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09404__A (.DIODE(_04529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08894__A (.DIODE(_04529_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09291__A1 (.DIODE(_04530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__A1 (.DIODE(_04530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09188__A1 (.DIODE(_04530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09152__A1 (.DIODE(_04530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09118__A1 (.DIODE(_04530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09047__A1 (.DIODE(_04530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09011__A1 (.DIODE(_04530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__A1 (.DIODE(_04530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08941__A1 (.DIODE(_04530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08895__A1 (.DIODE(_04530_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12800__A1 (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12557__A1 (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12418__A1 (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12349__A1 (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12315__A1 (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__A1 (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12177__A1 (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11987__A1 (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09407__A (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08898__A (.DIODE(_04532_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09293__A1 (.DIODE(_04533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09259__A1 (.DIODE(_04533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09190__A1 (.DIODE(_04533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09154__A1 (.DIODE(_04533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09120__A1 (.DIODE(_04533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09049__A1 (.DIODE(_04533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09013__A1 (.DIODE(_04533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08979__A1 (.DIODE(_04533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08943__A1 (.DIODE(_04533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08899__A1 (.DIODE(_04533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12802__A1 (.DIODE(_04535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12559__A1 (.DIODE(_04535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12420__A1 (.DIODE(_04535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12351__A1 (.DIODE(_04535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12317__A1 (.DIODE(_04535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12283__A1 (.DIODE(_04535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12179__A1 (.DIODE(_04535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11989__A1 (.DIODE(_04535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09410__A (.DIODE(_04535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08902__A (.DIODE(_04535_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09295__A1 (.DIODE(_04536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09261__A1 (.DIODE(_04536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09192__A1 (.DIODE(_04536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09156__A1 (.DIODE(_04536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09122__A1 (.DIODE(_04536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09051__A1 (.DIODE(_04536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09015__A1 (.DIODE(_04536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08981__A1 (.DIODE(_04536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08945__A1 (.DIODE(_04536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08903__A1 (.DIODE(_04536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12804__A1 (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12561__A1 (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12422__A1 (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12353__A1 (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12319__A1 (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12285__A1 (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12181__A1 (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11991__A1 (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09413__A (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08906__A (.DIODE(_04538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09297__A1 (.DIODE(_04539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09263__A1 (.DIODE(_04539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09194__A1 (.DIODE(_04539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09158__A1 (.DIODE(_04539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09124__A1 (.DIODE(_04539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09053__A1 (.DIODE(_04539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09017__A1 (.DIODE(_04539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08983__A1 (.DIODE(_04539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08947__A1 (.DIODE(_04539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__A1 (.DIODE(_04539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12806__A1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12563__A1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12424__A1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12355__A1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12321__A1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12287__A1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12183__A1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11993__A1 (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09416__A (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08910__A (.DIODE(_04541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09299__A1 (.DIODE(_04542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09265__A1 (.DIODE(_04542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__A1 (.DIODE(_04542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09160__A1 (.DIODE(_04542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__A1 (.DIODE(_04542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09055__A1 (.DIODE(_04542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09019__A1 (.DIODE(_04542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08985__A1 (.DIODE(_04542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08949__A1 (.DIODE(_04542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08911__A1 (.DIODE(_04542_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12808__A1 (.DIODE(_04544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12565__A1 (.DIODE(_04544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12426__A1 (.DIODE(_04544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12357__A1 (.DIODE(_04544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12323__A1 (.DIODE(_04544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12289__A1 (.DIODE(_04544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12185__A1 (.DIODE(_04544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11995__A1 (.DIODE(_04544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09419__A (.DIODE(_04544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08914__A (.DIODE(_04544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__A1 (.DIODE(_04545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__A1 (.DIODE(_04545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09198__A1 (.DIODE(_04545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__A1 (.DIODE(_04545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09128__A1 (.DIODE(_04545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09057__A1 (.DIODE(_04545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09021__A1 (.DIODE(_04545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08987__A1 (.DIODE(_04545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08951__A1 (.DIODE(_04545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08915__A1 (.DIODE(_04545_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12810__A1 (.DIODE(_04547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12567__A1 (.DIODE(_04547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12428__A1 (.DIODE(_04547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12359__A1 (.DIODE(_04547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12325__A1 (.DIODE(_04547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12291__A1 (.DIODE(_04547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12187__A1 (.DIODE(_04547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__A1 (.DIODE(_04547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09422__A (.DIODE(_04547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08918__A (.DIODE(_04547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09303__A1 (.DIODE(_04548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__A1 (.DIODE(_04548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__A1 (.DIODE(_04548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09164__A1 (.DIODE(_04548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09130__A1 (.DIODE(_04548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09059__A1 (.DIODE(_04548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09023__A1 (.DIODE(_04548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08989__A1 (.DIODE(_04548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08953__A1 (.DIODE(_04548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08919__A1 (.DIODE(_04548_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08941__S (.DIODE(_04551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08939__S (.DIODE(_04551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08937__S (.DIODE(_04551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08935__S (.DIODE(_04551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08933__S (.DIODE(_04551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08931__S (.DIODE(_04551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08929__S (.DIODE(_04551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08927__S (.DIODE(_04551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08925__S (.DIODE(_04551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08923__S (.DIODE(_04551_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12396__B (.DIODE(_04569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11826__B (.DIODE(_04569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11258__B (.DIODE(_04569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10676__B (.DIODE(_04569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10092__B (.DIODE(_04569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09989__B (.DIODE(_04569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09527__B (.DIODE(_04569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08957__B (.DIODE(_04569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08989__S (.DIODE(_04570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08987__S (.DIODE(_04570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08985__S (.DIODE(_04570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08983__S (.DIODE(_04570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08981__S (.DIODE(_04570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08979__S (.DIODE(_04570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08958__A (.DIODE(_04570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__S (.DIODE(_04571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08975__S (.DIODE(_04571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08973__S (.DIODE(_04571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08971__S (.DIODE(_04571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08969__S (.DIODE(_04571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08967__S (.DIODE(_04571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08965__S (.DIODE(_04571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08963__S (.DIODE(_04571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08961__S (.DIODE(_04571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08959__S (.DIODE(_04571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09023__S (.DIODE(_04588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09021__S (.DIODE(_04588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09019__S (.DIODE(_04588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09017__S (.DIODE(_04588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09015__S (.DIODE(_04588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09013__S (.DIODE(_04588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08992__A (.DIODE(_04588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09011__S (.DIODE(_04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09009__S (.DIODE(_04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09007__S (.DIODE(_04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09005__S (.DIODE(_04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09003__S (.DIODE(_04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09001__S (.DIODE(_04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08999__S (.DIODE(_04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08997__S (.DIODE(_04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08995__S (.DIODE(_04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08993__S (.DIODE(_04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12465__B (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11895__B (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11327__B (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10744__B (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10710__B (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10177__B (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09595__B (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09027__B (.DIODE(_04607_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09059__S (.DIODE(_04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09057__S (.DIODE(_04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09055__S (.DIODE(_04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09053__S (.DIODE(_04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09051__S (.DIODE(_04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09049__S (.DIODE(_04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09028__A (.DIODE(_04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09047__S (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09045__S (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09043__S (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09041__S (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09039__S (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09037__S (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09035__S (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09033__S (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09031__S (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09029__S (.DIODE(_04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09094__S (.DIODE(_04627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09092__S (.DIODE(_04627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09090__S (.DIODE(_04627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09088__S (.DIODE(_04627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__S (.DIODE(_04627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09084__S (.DIODE(_04627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09063__A (.DIODE(_04627_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09082__S (.DIODE(_04628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__S (.DIODE(_04628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09078__S (.DIODE(_04628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09076__S (.DIODE(_04628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09074__S (.DIODE(_04628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__S (.DIODE(_04628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__S (.DIODE(_04628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09068__S (.DIODE(_04628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09066__S (.DIODE(_04628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09064__S (.DIODE(_04628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__B (.DIODE(_04646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11965__B (.DIODE(_04646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11431__B (.DIODE(_04646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11397__B (.DIODE(_04646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10813__B (.DIODE(_04646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10247__B (.DIODE(_04646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09663__B (.DIODE(_04646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09098__B (.DIODE(_04646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09130__S (.DIODE(_04647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09128__S (.DIODE(_04647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__S (.DIODE(_04647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09124__S (.DIODE(_04647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09122__S (.DIODE(_04647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09120__S (.DIODE(_04647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09099__A (.DIODE(_04647_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09118__S (.DIODE(_04648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09116__S (.DIODE(_04648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09114__S (.DIODE(_04648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09112__S (.DIODE(_04648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09110__S (.DIODE(_04648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09108__S (.DIODE(_04648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09106__S (.DIODE(_04648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09104__S (.DIODE(_04648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09102__S (.DIODE(_04648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09100__S (.DIODE(_04648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09164__S (.DIODE(_04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__S (.DIODE(_04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09160__S (.DIODE(_04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09158__S (.DIODE(_04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09156__S (.DIODE(_04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09154__S (.DIODE(_04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09133__A (.DIODE(_04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09152__S (.DIODE(_04666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09150__S (.DIODE(_04666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09148__S (.DIODE(_04666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09146__S (.DIODE(_04666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09144__S (.DIODE(_04666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09142__S (.DIODE(_04666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09140__S (.DIODE(_04666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09138__S (.DIODE(_04666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09136__S (.DIODE(_04666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09134__S (.DIODE(_04666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12604__B (.DIODE(_04684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12155__B (.DIODE(_04684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12034__B (.DIODE(_04684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11465__B (.DIODE(_04684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10881__B (.DIODE(_04684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10316__B (.DIODE(_04684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09732__B (.DIODE(_04684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09168__B (.DIODE(_04684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09200__S (.DIODE(_04685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09198__S (.DIODE(_04685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__S (.DIODE(_04685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09194__S (.DIODE(_04685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09192__S (.DIODE(_04685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09190__S (.DIODE(_04685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09169__A (.DIODE(_04685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09188__S (.DIODE(_04686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09186__S (.DIODE(_04686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09184__S (.DIODE(_04686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09182__S (.DIODE(_04686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09180__S (.DIODE(_04686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09178__S (.DIODE(_04686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09176__S (.DIODE(_04686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09174__S (.DIODE(_04686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09172__S (.DIODE(_04686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09170__S (.DIODE(_04686_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09235__S (.DIODE(_04704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09233__S (.DIODE(_04704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09231__S (.DIODE(_04704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__S (.DIODE(_04704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09227__S (.DIODE(_04704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09225__S (.DIODE(_04704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09204__A (.DIODE(_04704_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09223__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09221__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09219__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09217__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09215__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09213__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09211__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09209__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09207__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09205__S (.DIODE(_04705_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__S (.DIODE(_04722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__S (.DIODE(_04722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09265__S (.DIODE(_04722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09263__S (.DIODE(_04722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09261__S (.DIODE(_04722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09259__S (.DIODE(_04722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09238__A (.DIODE(_04722_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__S (.DIODE(_04723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09255__S (.DIODE(_04723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__S (.DIODE(_04723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09251__S (.DIODE(_04723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09249__S (.DIODE(_04723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09247__S (.DIODE(_04723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09245__S (.DIODE(_04723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09243__S (.DIODE(_04723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09241__S (.DIODE(_04723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09239__S (.DIODE(_04723_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09291__S (.DIODE(_04741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09289__S (.DIODE(_04741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09287__S (.DIODE(_04741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09285__S (.DIODE(_04741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09283__S (.DIODE(_04741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09281__S (.DIODE(_04741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09279__S (.DIODE(_04741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09277__S (.DIODE(_04741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09275__S (.DIODE(_04741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09273__S (.DIODE(_04741_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09337__S (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09335__S (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09333__S (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09331__S (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09329__S (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09327__S (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09306__A (.DIODE(_04758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09325__S (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09323__S (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09321__S (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09319__S (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09317__S (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09315__S (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__S (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09311__S (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09309__S (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09307__S (.DIODE(_04759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09372__S (.DIODE(_04777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09370__S (.DIODE(_04777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09368__S (.DIODE(_04777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09366__S (.DIODE(_04777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09364__S (.DIODE(_04777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09362__S (.DIODE(_04777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09341__A (.DIODE(_04777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09360__S (.DIODE(_04778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09358__S (.DIODE(_04778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09356__S (.DIODE(_04778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09354__S (.DIODE(_04778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09352__S (.DIODE(_04778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09350__S (.DIODE(_04778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09348__S (.DIODE(_04778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09346__S (.DIODE(_04778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09344__S (.DIODE(_04778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09342__S (.DIODE(_04778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09699__A1 (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09665__A1 (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09631__A1 (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09597__A1 (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09563__A1 (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09529__A1 (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09495__A1 (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09461__A1 (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__A1 (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__A1 (.DIODE(_04795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09732__A (.DIODE(_04796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09697__B (.DIODE(_04796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09663__A (.DIODE(_04796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09595__A (.DIODE(_04796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09561__B (.DIODE(_04796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09527__A (.DIODE(_04796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09493__B (.DIODE(_04796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09459__A (.DIODE(_04796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09425__B (.DIODE(_04796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__A (.DIODE(_04796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__S (.DIODE(_04797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09420__S (.DIODE(_04797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09417__S (.DIODE(_04797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09414__S (.DIODE(_04797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09411__S (.DIODE(_04797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09408__S (.DIODE(_04797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09377__A (.DIODE(_04797_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09405__S (.DIODE(_04798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__S (.DIODE(_04798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09399__S (.DIODE(_04798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09396__S (.DIODE(_04798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09393__S (.DIODE(_04798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09390__S (.DIODE(_04798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__S (.DIODE(_04798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09384__S (.DIODE(_04798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09381__S (.DIODE(_04798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09378__S (.DIODE(_04798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09701__A1 (.DIODE(_04800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09667__A1 (.DIODE(_04800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09633__A1 (.DIODE(_04800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09599__A1 (.DIODE(_04800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09565__A1 (.DIODE(_04800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09531__A1 (.DIODE(_04800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09497__A1 (.DIODE(_04800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09463__A1 (.DIODE(_04800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__A1 (.DIODE(_04800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09381__A1 (.DIODE(_04800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__A1 (.DIODE(_04802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09669__A1 (.DIODE(_04802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09635__A1 (.DIODE(_04802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09601__A1 (.DIODE(_04802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09567__A1 (.DIODE(_04802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09533__A1 (.DIODE(_04802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__A1 (.DIODE(_04802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09465__A1 (.DIODE(_04802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09431__A1 (.DIODE(_04802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09384__A1 (.DIODE(_04802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__A1 (.DIODE(_04804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09671__A1 (.DIODE(_04804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09637__A1 (.DIODE(_04804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__A1 (.DIODE(_04804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09569__A1 (.DIODE(_04804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09535__A1 (.DIODE(_04804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09501__A1 (.DIODE(_04804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09467__A1 (.DIODE(_04804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09433__A1 (.DIODE(_04804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09387__A1 (.DIODE(_04804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__A1 (.DIODE(_04806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09673__A1 (.DIODE(_04806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09639__A1 (.DIODE(_04806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__A1 (.DIODE(_04806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09571__A1 (.DIODE(_04806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09537__A1 (.DIODE(_04806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09503__A1 (.DIODE(_04806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09469__A1 (.DIODE(_04806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09435__A1 (.DIODE(_04806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09390__A1 (.DIODE(_04806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__A1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__A1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09641__A1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__A1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09573__A1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09539__A1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09505__A1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09471__A1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09437__A1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09393__A1 (.DIODE(_04808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09711__A1 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__A1 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09643__A1 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__A1 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09575__A1 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__A1 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09507__A1 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09473__A1 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09439__A1 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09396__A1 (.DIODE(_04810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09713__A1 (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09679__A1 (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09645__A1 (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09611__A1 (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09577__A1 (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__A1 (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09509__A1 (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09475__A1 (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09441__A1 (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09399__A1 (.DIODE(_04812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__A1 (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09681__A1 (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09647__A1 (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09613__A1 (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09579__A1 (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09545__A1 (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__A1 (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09477__A1 (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09443__A1 (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09402__A1 (.DIODE(_04814_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09717__A1 (.DIODE(_04816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09683__A1 (.DIODE(_04816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09649__A1 (.DIODE(_04816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09615__A1 (.DIODE(_04816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__A1 (.DIODE(_04816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09547__A1 (.DIODE(_04816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09513__A1 (.DIODE(_04816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09479__A1 (.DIODE(_04816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__A1 (.DIODE(_04816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09405__A1 (.DIODE(_04816_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09719__A1 (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09685__A1 (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09651__A1 (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09617__A1 (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09583__A1 (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09549__A1 (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__A1 (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09481__A1 (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__A1 (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09408__A1 (.DIODE(_04818_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09721__A1 (.DIODE(_04820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09687__A1 (.DIODE(_04820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09653__A1 (.DIODE(_04820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09619__A1 (.DIODE(_04820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__A1 (.DIODE(_04820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09551__A1 (.DIODE(_04820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09517__A1 (.DIODE(_04820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09483__A1 (.DIODE(_04820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09449__A1 (.DIODE(_04820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09411__A1 (.DIODE(_04820_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09723__A1 (.DIODE(_04822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09689__A1 (.DIODE(_04822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09655__A1 (.DIODE(_04822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09621__A1 (.DIODE(_04822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09587__A1 (.DIODE(_04822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09553__A1 (.DIODE(_04822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09519__A1 (.DIODE(_04822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09485__A1 (.DIODE(_04822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09451__A1 (.DIODE(_04822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09414__A1 (.DIODE(_04822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09725__A1 (.DIODE(_04824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09691__A1 (.DIODE(_04824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09657__A1 (.DIODE(_04824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__A1 (.DIODE(_04824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09589__A1 (.DIODE(_04824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09555__A1 (.DIODE(_04824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09521__A1 (.DIODE(_04824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__A1 (.DIODE(_04824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09453__A1 (.DIODE(_04824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09417__A1 (.DIODE(_04824_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__A1 (.DIODE(_04826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09693__A1 (.DIODE(_04826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__A1 (.DIODE(_04826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__A1 (.DIODE(_04826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09591__A1 (.DIODE(_04826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09557__A1 (.DIODE(_04826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__A1 (.DIODE(_04826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09489__A1 (.DIODE(_04826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09455__A1 (.DIODE(_04826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09420__A1 (.DIODE(_04826_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09729__A1 (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09695__A1 (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09661__A1 (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09627__A1 (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09593__A1 (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09559__A1 (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09525__A1 (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09491__A1 (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09457__A1 (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__A1 (.DIODE(_04828_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09457__S (.DIODE(_04830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09455__S (.DIODE(_04830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09453__S (.DIODE(_04830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09451__S (.DIODE(_04830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09449__S (.DIODE(_04830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__S (.DIODE(_04830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09426__A (.DIODE(_04830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09445__S (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09443__S (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09441__S (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09439__S (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09437__S (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09435__S (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09433__S (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09431__S (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09429__S (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__S (.DIODE(_04831_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09491__S (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09489__S (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__S (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09485__S (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09483__S (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09481__S (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09460__A (.DIODE(_04848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09479__S (.DIODE(_04849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09477__S (.DIODE(_04849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09475__S (.DIODE(_04849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09473__S (.DIODE(_04849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09471__S (.DIODE(_04849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09469__S (.DIODE(_04849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09467__S (.DIODE(_04849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09465__S (.DIODE(_04849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09463__S (.DIODE(_04849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09461__S (.DIODE(_04849_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09525__S (.DIODE(_04866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__S (.DIODE(_04866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09521__S (.DIODE(_04866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09519__S (.DIODE(_04866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09517__S (.DIODE(_04866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__S (.DIODE(_04866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09494__A (.DIODE(_04866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09513__S (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__S (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09509__S (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09507__S (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09505__S (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09503__S (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09501__S (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__S (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09497__S (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09495__S (.DIODE(_04867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09559__S (.DIODE(_04884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09557__S (.DIODE(_04884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09555__S (.DIODE(_04884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09553__S (.DIODE(_04884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09551__S (.DIODE(_04884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09549__S (.DIODE(_04884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09528__A (.DIODE(_04884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09547__S (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09545__S (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__S (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__S (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09539__S (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09537__S (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09535__S (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09533__S (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09531__S (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09529__S (.DIODE(_04885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09593__S (.DIODE(_04902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09591__S (.DIODE(_04902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09589__S (.DIODE(_04902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09587__S (.DIODE(_04902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09585__S (.DIODE(_04902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09583__S (.DIODE(_04902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09562__A (.DIODE(_04902_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09581__S (.DIODE(_04903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09579__S (.DIODE(_04903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09577__S (.DIODE(_04903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09575__S (.DIODE(_04903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09573__S (.DIODE(_04903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09571__S (.DIODE(_04903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09569__S (.DIODE(_04903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09567__S (.DIODE(_04903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09565__S (.DIODE(_04903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09563__S (.DIODE(_04903_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09627__S (.DIODE(_04920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09625__S (.DIODE(_04920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__S (.DIODE(_04920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09621__S (.DIODE(_04920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09619__S (.DIODE(_04920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09617__S (.DIODE(_04920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09596__A (.DIODE(_04920_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09615__S (.DIODE(_04921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09613__S (.DIODE(_04921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09611__S (.DIODE(_04921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__S (.DIODE(_04921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09607__S (.DIODE(_04921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__S (.DIODE(_04921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09603__S (.DIODE(_04921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09601__S (.DIODE(_04921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09599__S (.DIODE(_04921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09597__S (.DIODE(_04921_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09695__S (.DIODE(_04956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09693__S (.DIODE(_04956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09691__S (.DIODE(_04956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09689__S (.DIODE(_04956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09687__S (.DIODE(_04956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09685__S (.DIODE(_04956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09664__A (.DIODE(_04956_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09683__S (.DIODE(_04957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09681__S (.DIODE(_04957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09679__S (.DIODE(_04957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09677__S (.DIODE(_04957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__S (.DIODE(_04957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09673__S (.DIODE(_04957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09671__S (.DIODE(_04957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09669__S (.DIODE(_04957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09667__S (.DIODE(_04957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09665__S (.DIODE(_04957_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09729__S (.DIODE(_04974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__S (.DIODE(_04974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09725__S (.DIODE(_04974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09723__S (.DIODE(_04974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09721__S (.DIODE(_04974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09719__S (.DIODE(_04974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__A (.DIODE(_04974_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09717__S (.DIODE(_04975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__S (.DIODE(_04975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09713__S (.DIODE(_04975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09711__S (.DIODE(_04975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09709__S (.DIODE(_04975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__S (.DIODE(_04975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09705__S (.DIODE(_04975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__S (.DIODE(_04975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09701__S (.DIODE(_04975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09699__S (.DIODE(_04975_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10560__A1 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10526__A1 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10353__A1 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__A1 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__A1 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10025__A1 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09991__A1 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09957__A1 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09819__A1 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09734__A1 (.DIODE(_04992_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__S (.DIODE(_04993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09776__S (.DIODE(_04993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09773__S (.DIODE(_04993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09770__S (.DIODE(_04993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09767__S (.DIODE(_04993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09764__S (.DIODE(_04993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09733__A (.DIODE(_04993_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09761__S (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09758__S (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09755__S (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09752__S (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__S (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09746__S (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09743__S (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09740__S (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09737__S (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09734__S (.DIODE(_04994_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10562__A1 (.DIODE(_04996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10528__A1 (.DIODE(_04996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10355__A1 (.DIODE(_04996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10251__A1 (.DIODE(_04996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10096__A1 (.DIODE(_04996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10027__A1 (.DIODE(_04996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09993__A1 (.DIODE(_04996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09959__A1 (.DIODE(_04996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09821__A1 (.DIODE(_04996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09737__A1 (.DIODE(_04996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__A1 (.DIODE(_04998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10530__A1 (.DIODE(_04998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__A1 (.DIODE(_04998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10253__A1 (.DIODE(_04998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10098__A1 (.DIODE(_04998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10029__A1 (.DIODE(_04998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09995__A1 (.DIODE(_04998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09961__A1 (.DIODE(_04998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09823__A1 (.DIODE(_04998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09740__A1 (.DIODE(_04998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10566__A1 (.DIODE(_05000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10532__A1 (.DIODE(_05000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__A1 (.DIODE(_05000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10255__A1 (.DIODE(_05000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10100__A1 (.DIODE(_05000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10031__A1 (.DIODE(_05000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09997__A1 (.DIODE(_05000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09963__A1 (.DIODE(_05000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__A1 (.DIODE(_05000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09743__A1 (.DIODE(_05000_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10568__A1 (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10534__A1 (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10361__A1 (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10257__A1 (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10102__A1 (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10033__A1 (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09999__A1 (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09965__A1 (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09827__A1 (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09746__A1 (.DIODE(_05002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10570__A1 (.DIODE(_05004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10536__A1 (.DIODE(_05004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10363__A1 (.DIODE(_05004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10259__A1 (.DIODE(_05004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10104__A1 (.DIODE(_05004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10035__A1 (.DIODE(_05004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10001__A1 (.DIODE(_05004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09967__A1 (.DIODE(_05004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09829__A1 (.DIODE(_05004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__A1 (.DIODE(_05004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10572__A1 (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10538__A1 (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10365__A1 (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10261__A1 (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10106__A1 (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10037__A1 (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10003__A1 (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09969__A1 (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09831__A1 (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09752__A1 (.DIODE(_05006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10574__A1 (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10540__A1 (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10367__A1 (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10263__A1 (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10108__A1 (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10039__A1 (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10005__A1 (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09971__A1 (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09833__A1 (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09755__A1 (.DIODE(_05008_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10576__A1 (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10542__A1 (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10369__A1 (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10265__A1 (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10110__A1 (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10041__A1 (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__A1 (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09973__A1 (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09835__A1 (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09758__A1 (.DIODE(_05010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10578__A1 (.DIODE(_05012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10544__A1 (.DIODE(_05012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10371__A1 (.DIODE(_05012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10267__A1 (.DIODE(_05012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10112__A1 (.DIODE(_05012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__A1 (.DIODE(_05012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10009__A1 (.DIODE(_05012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09975__A1 (.DIODE(_05012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09837__A1 (.DIODE(_05012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09761__A1 (.DIODE(_05012_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10580__A1 (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10546__A1 (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10373__A1 (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10269__A1 (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10114__A1 (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10045__A1 (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10011__A1 (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09977__A1 (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09839__A1 (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09764__A1 (.DIODE(_05014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10582__A1 (.DIODE(_05016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10548__A1 (.DIODE(_05016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__A1 (.DIODE(_05016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10271__A1 (.DIODE(_05016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10116__A1 (.DIODE(_05016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10047__A1 (.DIODE(_05016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10013__A1 (.DIODE(_05016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09979__A1 (.DIODE(_05016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09841__A1 (.DIODE(_05016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09767__A1 (.DIODE(_05016_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10584__A1 (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10550__A1 (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10377__A1 (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10273__A1 (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10118__A1 (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10049__A1 (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10015__A1 (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09981__A1 (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09843__A1 (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09770__A1 (.DIODE(_05018_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10586__A1 (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10552__A1 (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__A1 (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10275__A1 (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10120__A1 (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10051__A1 (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10017__A1 (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09983__A1 (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09845__A1 (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09773__A1 (.DIODE(_05020_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10588__A1 (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10554__A1 (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10381__A1 (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10277__A1 (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10122__A1 (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10053__A1 (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10019__A1 (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09985__A1 (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09847__A1 (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09776__A1 (.DIODE(_05022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10590__A1 (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10556__A1 (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10383__A1 (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10279__A1 (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10124__A1 (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10055__A1 (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10021__A1 (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09987__A1 (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09849__A1 (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__A1 (.DIODE(_05024_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11655__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11500__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11362__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11069__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10916__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10778__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10489__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10212__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09920__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09782__B (.DIODE(_05026_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09815__S (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09813__S (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09811__S (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09809__S (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09807__S (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__S (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09784__A (.DIODE(_05028_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09803__S (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__S (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09799__S (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09797__S (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__S (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09793__S (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09791__S (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09789__S (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09787__S (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09785__S (.DIODE(_05029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09849__S (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09847__S (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09845__S (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09843__S (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09841__S (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09839__S (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09818__A (.DIODE(_05046_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09837__S (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09835__S (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09833__S (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09831__S (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09829__S (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09827__S (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09825__S (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09823__S (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09821__S (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09819__S (.DIODE(_05047_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09884__S (.DIODE(_05065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09882__S (.DIODE(_05065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09880__S (.DIODE(_05065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09878__S (.DIODE(_05065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09876__S (.DIODE(_05065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09874__S (.DIODE(_05065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09853__A (.DIODE(_05065_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09872__S (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09870__S (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09868__S (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09866__S (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09864__S (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09862__S (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09860__S (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09858__S (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09856__S (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09854__S (.DIODE(_05066_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09918__S (.DIODE(_05083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09916__S (.DIODE(_05083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09914__S (.DIODE(_05083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09912__S (.DIODE(_05083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__S (.DIODE(_05083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09908__S (.DIODE(_05083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09887__A (.DIODE(_05083_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09906__S (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09904__S (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09902__S (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__S (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09898__S (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09896__S (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09894__S (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09892__S (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09890__S (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09888__S (.DIODE(_05084_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09953__S (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__S (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__S (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09947__S (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09945__S (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09943__S (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09922__A (.DIODE(_05102_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__S (.DIODE(_05103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__S (.DIODE(_05103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09937__S (.DIODE(_05103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__S (.DIODE(_05103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09933__S (.DIODE(_05103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09931__S (.DIODE(_05103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09929__S (.DIODE(_05103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09927__S (.DIODE(_05103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09925__S (.DIODE(_05103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09923__S (.DIODE(_05103_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09975__S (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09973__S (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09971__S (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09969__S (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09967__S (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09965__S (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09963__S (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09961__S (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09959__S (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09957__S (.DIODE(_05121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10021__S (.DIODE(_05138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10019__S (.DIODE(_05138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10017__S (.DIODE(_05138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10015__S (.DIODE(_05138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10013__S (.DIODE(_05138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10011__S (.DIODE(_05138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09990__A (.DIODE(_05138_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10009__S (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__S (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10005__S (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10003__S (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10001__S (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09999__S (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09997__S (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09995__S (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09993__S (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09991__S (.DIODE(_05139_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10043__S (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10041__S (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10039__S (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10037__S (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10035__S (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10033__S (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10031__S (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10029__S (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10027__S (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10025__S (.DIODE(_05157_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10078__S (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10076__S (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10074__S (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10072__S (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10070__S (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10068__S (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10066__S (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10064__S (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10062__S (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10060__S (.DIODE(_05176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10124__S (.DIODE(_05193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10122__S (.DIODE(_05193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10120__S (.DIODE(_05193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10118__S (.DIODE(_05193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10116__S (.DIODE(_05193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10114__S (.DIODE(_05193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10093__A (.DIODE(_05193_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10112__S (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10110__S (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10108__S (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10106__S (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10104__S (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10102__S (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10100__S (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10098__S (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10096__S (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10094__S (.DIODE(_05194_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10781__A0 (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__A0 (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10457__A0 (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10423__A0 (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10388__A0 (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10319__A0 (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10284__A0 (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10215__A0 (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10180__A0 (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10130__A0 (.DIODE(_05211_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10175__S (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10172__S (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10169__S (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10166__S (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10163__S (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10160__S (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10129__A (.DIODE(_05213_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10157__S (.DIODE(_05214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__S (.DIODE(_05214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__S (.DIODE(_05214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10148__S (.DIODE(_05214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10145__S (.DIODE(_05214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10142__S (.DIODE(_05214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10139__S (.DIODE(_05214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10136__S (.DIODE(_05214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10133__S (.DIODE(_05214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10130__S (.DIODE(_05214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10783__A0 (.DIODE(_05216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10494__A0 (.DIODE(_05216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10459__A0 (.DIODE(_05216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10425__A0 (.DIODE(_05216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10390__A0 (.DIODE(_05216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10321__A0 (.DIODE(_05216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10286__A0 (.DIODE(_05216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10217__A0 (.DIODE(_05216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10182__A0 (.DIODE(_05216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10133__A0 (.DIODE(_05216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10785__A0 (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10496__A0 (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10461__A0 (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10427__A0 (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10392__A0 (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10323__A0 (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10288__A0 (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10219__A0 (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10184__A0 (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10136__A0 (.DIODE(_05218_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10787__A0 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10498__A0 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10463__A0 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10429__A0 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10394__A0 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10325__A0 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10290__A0 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10221__A0 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10186__A0 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10139__A0 (.DIODE(_05220_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10789__A0 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10500__A0 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10465__A0 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10431__A0 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10396__A0 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__A0 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10292__A0 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10223__A0 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__A0 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10142__A0 (.DIODE(_05222_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10791__A0 (.DIODE(_05224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__A0 (.DIODE(_05224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10467__A0 (.DIODE(_05224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10433__A0 (.DIODE(_05224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10398__A0 (.DIODE(_05224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__A0 (.DIODE(_05224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10294__A0 (.DIODE(_05224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10225__A0 (.DIODE(_05224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10190__A0 (.DIODE(_05224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10145__A0 (.DIODE(_05224_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10793__A0 (.DIODE(_05226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10504__A0 (.DIODE(_05226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10469__A0 (.DIODE(_05226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10435__A0 (.DIODE(_05226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10400__A0 (.DIODE(_05226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10331__A0 (.DIODE(_05226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10296__A0 (.DIODE(_05226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10227__A0 (.DIODE(_05226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10192__A0 (.DIODE(_05226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10148__A0 (.DIODE(_05226_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10795__A0 (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10506__A0 (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10471__A0 (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10437__A0 (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10402__A0 (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10333__A0 (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__A0 (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10229__A0 (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__A0 (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__A0 (.DIODE(_05228_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10797__A0 (.DIODE(_05230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__A0 (.DIODE(_05230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10473__A0 (.DIODE(_05230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10439__A0 (.DIODE(_05230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10404__A0 (.DIODE(_05230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__A0 (.DIODE(_05230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10300__A0 (.DIODE(_05230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__A0 (.DIODE(_05230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__A0 (.DIODE(_05230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__A0 (.DIODE(_05230_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10799__A0 (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10510__A0 (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10475__A0 (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10441__A0 (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__A0 (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10337__A0 (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10302__A0 (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__A0 (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10198__A0 (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10157__A0 (.DIODE(_05232_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10801__A0 (.DIODE(_05234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10512__A0 (.DIODE(_05234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10477__A0 (.DIODE(_05234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__A0 (.DIODE(_05234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10408__A0 (.DIODE(_05234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10339__A0 (.DIODE(_05234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10304__A0 (.DIODE(_05234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10235__A0 (.DIODE(_05234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10200__A0 (.DIODE(_05234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10160__A0 (.DIODE(_05234_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10803__A0 (.DIODE(_05236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10514__A0 (.DIODE(_05236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10479__A0 (.DIODE(_05236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10445__A0 (.DIODE(_05236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10410__A0 (.DIODE(_05236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10341__A0 (.DIODE(_05236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10306__A0 (.DIODE(_05236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10237__A0 (.DIODE(_05236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10202__A0 (.DIODE(_05236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10163__A0 (.DIODE(_05236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10805__A0 (.DIODE(_05238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10516__A0 (.DIODE(_05238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10481__A0 (.DIODE(_05238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__A0 (.DIODE(_05238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10412__A0 (.DIODE(_05238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10343__A0 (.DIODE(_05238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10308__A0 (.DIODE(_05238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10239__A0 (.DIODE(_05238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10204__A0 (.DIODE(_05238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10166__A0 (.DIODE(_05238_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10807__A0 (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10518__A0 (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10483__A0 (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10449__A0 (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10414__A0 (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10345__A0 (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10310__A0 (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10241__A0 (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10206__A0 (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10169__A0 (.DIODE(_05240_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10809__A0 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10520__A0 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10485__A0 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10451__A0 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10416__A0 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10347__A0 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10312__A0 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10243__A0 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10208__A0 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10172__A0 (.DIODE(_05242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__A0 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10522__A0 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10487__A0 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10453__A0 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__A0 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10349__A0 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10314__A0 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10245__A0 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10210__A0 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10175__A0 (.DIODE(_05244_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10210__S (.DIODE(_05247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10208__S (.DIODE(_05247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10206__S (.DIODE(_05247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10204__S (.DIODE(_05247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10202__S (.DIODE(_05247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10200__S (.DIODE(_05247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10179__A (.DIODE(_05247_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10198__S (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__S (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__S (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10192__S (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10190__S (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10188__S (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10186__S (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10184__S (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10182__S (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10180__S (.DIODE(_05248_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10245__S (.DIODE(_05266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10243__S (.DIODE(_05266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10241__S (.DIODE(_05266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10239__S (.DIODE(_05266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10237__S (.DIODE(_05266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10235__S (.DIODE(_05266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10214__A (.DIODE(_05266_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__S (.DIODE(_05267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__S (.DIODE(_05267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10229__S (.DIODE(_05267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10227__S (.DIODE(_05267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10225__S (.DIODE(_05267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10223__S (.DIODE(_05267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10221__S (.DIODE(_05267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10219__S (.DIODE(_05267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10217__S (.DIODE(_05267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10215__S (.DIODE(_05267_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10267__S (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10265__S (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10263__S (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10261__S (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10259__S (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10257__S (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10255__S (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10253__S (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10251__S (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__S (.DIODE(_05285_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10302__S (.DIODE(_05304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10300__S (.DIODE(_05304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__S (.DIODE(_05304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10296__S (.DIODE(_05304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10294__S (.DIODE(_05304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10292__S (.DIODE(_05304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10290__S (.DIODE(_05304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10288__S (.DIODE(_05304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10286__S (.DIODE(_05304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10284__S (.DIODE(_05304_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10349__S (.DIODE(_05322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10347__S (.DIODE(_05322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10345__S (.DIODE(_05322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10343__S (.DIODE(_05322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10341__S (.DIODE(_05322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10339__S (.DIODE(_05322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10318__A (.DIODE(_05322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10337__S (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__S (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10333__S (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10331__S (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__S (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__S (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10325__S (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10323__S (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10321__S (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10319__S (.DIODE(_05323_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10383__S (.DIODE(_05340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10381__S (.DIODE(_05340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__S (.DIODE(_05340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10377__S (.DIODE(_05340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__S (.DIODE(_05340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10373__S (.DIODE(_05340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10352__A (.DIODE(_05340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__S (.DIODE(_05359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10416__S (.DIODE(_05359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10414__S (.DIODE(_05359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10412__S (.DIODE(_05359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10410__S (.DIODE(_05359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10408__S (.DIODE(_05359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10387__A (.DIODE(_05359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__S (.DIODE(_05360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10404__S (.DIODE(_05360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10402__S (.DIODE(_05360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10400__S (.DIODE(_05360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10398__S (.DIODE(_05360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10396__S (.DIODE(_05360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10394__S (.DIODE(_05360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10392__S (.DIODE(_05360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10390__S (.DIODE(_05360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10388__S (.DIODE(_05360_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10453__S (.DIODE(_05378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10451__S (.DIODE(_05378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10449__S (.DIODE(_05378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__S (.DIODE(_05378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10445__S (.DIODE(_05378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__S (.DIODE(_05378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10422__A (.DIODE(_05378_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10441__S (.DIODE(_05379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10439__S (.DIODE(_05379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10437__S (.DIODE(_05379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10435__S (.DIODE(_05379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10433__S (.DIODE(_05379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10431__S (.DIODE(_05379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10429__S (.DIODE(_05379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10427__S (.DIODE(_05379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10425__S (.DIODE(_05379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10423__S (.DIODE(_05379_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10487__S (.DIODE(_05396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10485__S (.DIODE(_05396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10483__S (.DIODE(_05396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10481__S (.DIODE(_05396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10479__S (.DIODE(_05396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10477__S (.DIODE(_05396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10456__A (.DIODE(_05396_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10475__S (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10473__S (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10471__S (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10469__S (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10467__S (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10465__S (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10463__S (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10461__S (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10459__S (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10457__S (.DIODE(_05397_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10522__S (.DIODE(_05415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10520__S (.DIODE(_05415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10518__S (.DIODE(_05415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10516__S (.DIODE(_05415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10514__S (.DIODE(_05415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10512__S (.DIODE(_05415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10491__A (.DIODE(_05415_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10510__S (.DIODE(_05416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__S (.DIODE(_05416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10506__S (.DIODE(_05416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10504__S (.DIODE(_05416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__S (.DIODE(_05416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10500__S (.DIODE(_05416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10498__S (.DIODE(_05416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10496__S (.DIODE(_05416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10494__S (.DIODE(_05416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__S (.DIODE(_05416_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10556__S (.DIODE(_05433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10554__S (.DIODE(_05433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10552__S (.DIODE(_05433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10550__S (.DIODE(_05433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10548__S (.DIODE(_05433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10546__S (.DIODE(_05433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10525__A (.DIODE(_05433_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10544__S (.DIODE(_05434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10542__S (.DIODE(_05434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10540__S (.DIODE(_05434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10538__S (.DIODE(_05434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10536__S (.DIODE(_05434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10534__S (.DIODE(_05434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10532__S (.DIODE(_05434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10530__S (.DIODE(_05434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10528__S (.DIODE(_05434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10526__S (.DIODE(_05434_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10590__S (.DIODE(_05451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10588__S (.DIODE(_05451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10586__S (.DIODE(_05451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10584__S (.DIODE(_05451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10582__S (.DIODE(_05451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10580__S (.DIODE(_05451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10559__A (.DIODE(_05451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10578__S (.DIODE(_05452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10576__S (.DIODE(_05452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10574__S (.DIODE(_05452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10572__S (.DIODE(_05452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10570__S (.DIODE(_05452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10568__S (.DIODE(_05452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10566__S (.DIODE(_05452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__S (.DIODE(_05452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10562__S (.DIODE(_05452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10560__S (.DIODE(_05452_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11107__A1 (.DIODE(_05469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10968__A1 (.DIODE(_05469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10883__A1 (.DIODE(_05469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__A1 (.DIODE(_05469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10815__A1 (.DIODE(_05469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10746__A1 (.DIODE(_05469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10712__A1 (.DIODE(_05469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__A1 (.DIODE(_05469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__A1 (.DIODE(_05469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__A1 (.DIODE(_05469_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10622__S (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10619__S (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10616__S (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10613__S (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10610__S (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__S (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10604__S (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10601__S (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10598__S (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__S (.DIODE(_05471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11109__A1 (.DIODE(_05473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10970__A1 (.DIODE(_05473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10885__A1 (.DIODE(_05473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10851__A1 (.DIODE(_05473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10817__A1 (.DIODE(_05473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10748__A1 (.DIODE(_05473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10714__A1 (.DIODE(_05473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10680__A1 (.DIODE(_05473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10646__A1 (.DIODE(_05473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10598__A1 (.DIODE(_05473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11111__A1 (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10972__A1 (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10887__A1 (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10853__A1 (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10819__A1 (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10750__A1 (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__A1 (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10682__A1 (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__A1 (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10601__A1 (.DIODE(_05475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11113__A1 (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10974__A1 (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10889__A1 (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10855__A1 (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10821__A1 (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10752__A1 (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10718__A1 (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10684__A1 (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10650__A1 (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10604__A1 (.DIODE(_05477_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11115__A1 (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10976__A1 (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10891__A1 (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10857__A1 (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10823__A1 (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10754__A1 (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10720__A1 (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10686__A1 (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10652__A1 (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__A1 (.DIODE(_05479_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11117__A1 (.DIODE(_05481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10978__A1 (.DIODE(_05481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10893__A1 (.DIODE(_05481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10859__A1 (.DIODE(_05481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10825__A1 (.DIODE(_05481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10756__A1 (.DIODE(_05481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10722__A1 (.DIODE(_05481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10688__A1 (.DIODE(_05481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__A1 (.DIODE(_05481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10610__A1 (.DIODE(_05481_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11119__A1 (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__A1 (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10895__A1 (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10861__A1 (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10827__A1 (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10758__A1 (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10724__A1 (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10690__A1 (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10656__A1 (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10613__A1 (.DIODE(_05483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11121__A1 (.DIODE(_05485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10982__A1 (.DIODE(_05485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10897__A1 (.DIODE(_05485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10863__A1 (.DIODE(_05485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10829__A1 (.DIODE(_05485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10760__A1 (.DIODE(_05485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10726__A1 (.DIODE(_05485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10692__A1 (.DIODE(_05485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10658__A1 (.DIODE(_05485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10616__A1 (.DIODE(_05485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11123__A1 (.DIODE(_05487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10984__A1 (.DIODE(_05487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10899__A1 (.DIODE(_05487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10865__A1 (.DIODE(_05487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10831__A1 (.DIODE(_05487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10762__A1 (.DIODE(_05487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10728__A1 (.DIODE(_05487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10694__A1 (.DIODE(_05487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10660__A1 (.DIODE(_05487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10619__A1 (.DIODE(_05487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11125__A1 (.DIODE(_05489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10986__A1 (.DIODE(_05489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10901__A1 (.DIODE(_05489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10867__A1 (.DIODE(_05489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10833__A1 (.DIODE(_05489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10764__A1 (.DIODE(_05489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10730__A1 (.DIODE(_05489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10696__A1 (.DIODE(_05489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10662__A1 (.DIODE(_05489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10622__A1 (.DIODE(_05489_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11127__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10988__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10903__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10869__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10835__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10766__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10732__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10698__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10664__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10625__A1 (.DIODE(_05491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11129__A1 (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10990__A1 (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10905__A1 (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10871__A1 (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10837__A1 (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10768__A1 (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10734__A1 (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__A1 (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__A1 (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__A1 (.DIODE(_05493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11131__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10992__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10907__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10873__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10839__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10770__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10736__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10702__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10668__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10631__A1 (.DIODE(_05495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11133__A1 (.DIODE(_05497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10994__A1 (.DIODE(_05497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10909__A1 (.DIODE(_05497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10875__A1 (.DIODE(_05497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10841__A1 (.DIODE(_05497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10772__A1 (.DIODE(_05497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10738__A1 (.DIODE(_05497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10704__A1 (.DIODE(_05497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10670__A1 (.DIODE(_05497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10634__A1 (.DIODE(_05497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11135__A1 (.DIODE(_05499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10996__A1 (.DIODE(_05499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10911__A1 (.DIODE(_05499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10877__A1 (.DIODE(_05499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10843__A1 (.DIODE(_05499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10774__A1 (.DIODE(_05499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10740__A1 (.DIODE(_05499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__A1 (.DIODE(_05499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10672__A1 (.DIODE(_05499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10637__A1 (.DIODE(_05499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11137__A1 (.DIODE(_05501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10998__A1 (.DIODE(_05501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10913__A1 (.DIODE(_05501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10879__A1 (.DIODE(_05501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10845__A1 (.DIODE(_05501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10776__A1 (.DIODE(_05501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10742__A1 (.DIODE(_05501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10708__A1 (.DIODE(_05501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__A1 (.DIODE(_05501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10640__A1 (.DIODE(_05501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10662__S (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10660__S (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10658__S (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10656__S (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__S (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10652__S (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10650__S (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__S (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10646__S (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__S (.DIODE(_05504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10708__S (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__S (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10704__S (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10702__S (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10700__S (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10698__S (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10677__A (.DIODE(_05521_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10696__S (.DIODE(_05522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10694__S (.DIODE(_05522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10692__S (.DIODE(_05522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10690__S (.DIODE(_05522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10688__S (.DIODE(_05522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10686__S (.DIODE(_05522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10684__S (.DIODE(_05522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10682__S (.DIODE(_05522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10680__S (.DIODE(_05522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__S (.DIODE(_05522_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10742__S (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10740__S (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10738__S (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10736__S (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10734__S (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10732__S (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10711__A (.DIODE(_05539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10730__S (.DIODE(_05540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10728__S (.DIODE(_05540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10726__S (.DIODE(_05540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10724__S (.DIODE(_05540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10722__S (.DIODE(_05540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10720__S (.DIODE(_05540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10718__S (.DIODE(_05540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__S (.DIODE(_05540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10714__S (.DIODE(_05540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10712__S (.DIODE(_05540_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10776__S (.DIODE(_05557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10774__S (.DIODE(_05557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10772__S (.DIODE(_05557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10770__S (.DIODE(_05557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10768__S (.DIODE(_05557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10766__S (.DIODE(_05557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10745__A (.DIODE(_05557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10764__S (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10762__S (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10760__S (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10758__S (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10756__S (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10754__S (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10752__S (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10750__S (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10748__S (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10746__S (.DIODE(_05558_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10811__S (.DIODE(_05576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10809__S (.DIODE(_05576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10807__S (.DIODE(_05576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10805__S (.DIODE(_05576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10803__S (.DIODE(_05576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10801__S (.DIODE(_05576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10780__A (.DIODE(_05576_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10799__S (.DIODE(_05577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10797__S (.DIODE(_05577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10795__S (.DIODE(_05577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10793__S (.DIODE(_05577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10791__S (.DIODE(_05577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10789__S (.DIODE(_05577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10787__S (.DIODE(_05577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10785__S (.DIODE(_05577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10783__S (.DIODE(_05577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10781__S (.DIODE(_05577_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10845__S (.DIODE(_05594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10843__S (.DIODE(_05594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10841__S (.DIODE(_05594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10839__S (.DIODE(_05594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10837__S (.DIODE(_05594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10835__S (.DIODE(_05594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10814__A (.DIODE(_05594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10833__S (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10831__S (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10829__S (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10827__S (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10825__S (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10823__S (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10821__S (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10819__S (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10817__S (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10815__S (.DIODE(_05595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10879__S (.DIODE(_05612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10877__S (.DIODE(_05612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10875__S (.DIODE(_05612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10873__S (.DIODE(_05612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10871__S (.DIODE(_05612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10869__S (.DIODE(_05612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10848__A (.DIODE(_05612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10867__S (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10865__S (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10863__S (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10861__S (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10859__S (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10857__S (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10855__S (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10853__S (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10851__S (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10849__S (.DIODE(_05613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10913__S (.DIODE(_05630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10911__S (.DIODE(_05630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10909__S (.DIODE(_05630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10907__S (.DIODE(_05630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10905__S (.DIODE(_05630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10903__S (.DIODE(_05630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10882__A (.DIODE(_05630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10901__S (.DIODE(_05631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10899__S (.DIODE(_05631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10897__S (.DIODE(_05631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10895__S (.DIODE(_05631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10893__S (.DIODE(_05631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10891__S (.DIODE(_05631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10889__S (.DIODE(_05631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10887__S (.DIODE(_05631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10885__S (.DIODE(_05631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10883__S (.DIODE(_05631_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11503__A0 (.DIODE(_05648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11468__A0 (.DIODE(_05648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11365__A0 (.DIODE(_05648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11330__A0 (.DIODE(_05648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11295__A0 (.DIODE(_05648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11226__A0 (.DIODE(_05648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11072__A0 (.DIODE(_05648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11037__A0 (.DIODE(_05648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11003__A0 (.DIODE(_05648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__A0 (.DIODE(_05648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10964__S (.DIODE(_05650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10961__S (.DIODE(_05650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10958__S (.DIODE(_05650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__S (.DIODE(_05650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10952__S (.DIODE(_05650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10949__S (.DIODE(_05650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10918__A (.DIODE(_05650_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10946__S (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__S (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__S (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10937__S (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10934__S (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10931__S (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10928__S (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10925__S (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10922__S (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__S (.DIODE(_05651_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11505__A0 (.DIODE(_05653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11470__A0 (.DIODE(_05653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11367__A0 (.DIODE(_05653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11332__A0 (.DIODE(_05653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11297__A0 (.DIODE(_05653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11228__A0 (.DIODE(_05653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11074__A0 (.DIODE(_05653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11039__A0 (.DIODE(_05653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11005__A0 (.DIODE(_05653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10922__A0 (.DIODE(_05653_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11507__A0 (.DIODE(_05655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11472__A0 (.DIODE(_05655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11369__A0 (.DIODE(_05655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11334__A0 (.DIODE(_05655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11299__A0 (.DIODE(_05655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11230__A0 (.DIODE(_05655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11076__A0 (.DIODE(_05655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__A0 (.DIODE(_05655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11007__A0 (.DIODE(_05655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10925__A0 (.DIODE(_05655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11509__A0 (.DIODE(_05657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11474__A0 (.DIODE(_05657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11371__A0 (.DIODE(_05657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11336__A0 (.DIODE(_05657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11301__A0 (.DIODE(_05657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11232__A0 (.DIODE(_05657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11078__A0 (.DIODE(_05657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11043__A0 (.DIODE(_05657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11009__A0 (.DIODE(_05657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10928__A0 (.DIODE(_05657_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11511__A0 (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__A0 (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11373__A0 (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11338__A0 (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11303__A0 (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11234__A0 (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11080__A0 (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11045__A0 (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11011__A0 (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10931__A0 (.DIODE(_05659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11513__A0 (.DIODE(_05661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11478__A0 (.DIODE(_05661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11375__A0 (.DIODE(_05661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11340__A0 (.DIODE(_05661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11305__A0 (.DIODE(_05661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11236__A0 (.DIODE(_05661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11082__A0 (.DIODE(_05661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11047__A0 (.DIODE(_05661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11013__A0 (.DIODE(_05661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10934__A0 (.DIODE(_05661_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11515__A0 (.DIODE(_05663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11480__A0 (.DIODE(_05663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__A0 (.DIODE(_05663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11342__A0 (.DIODE(_05663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11307__A0 (.DIODE(_05663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11238__A0 (.DIODE(_05663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11084__A0 (.DIODE(_05663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11049__A0 (.DIODE(_05663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11015__A0 (.DIODE(_05663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10937__A0 (.DIODE(_05663_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__A0 (.DIODE(_05665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11482__A0 (.DIODE(_05665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11379__A0 (.DIODE(_05665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11344__A0 (.DIODE(_05665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11309__A0 (.DIODE(_05665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11240__A0 (.DIODE(_05665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11086__A0 (.DIODE(_05665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11051__A0 (.DIODE(_05665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11017__A0 (.DIODE(_05665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__A0 (.DIODE(_05665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11519__A0 (.DIODE(_05667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11484__A0 (.DIODE(_05667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11381__A0 (.DIODE(_05667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11346__A0 (.DIODE(_05667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11311__A0 (.DIODE(_05667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11242__A0 (.DIODE(_05667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11088__A0 (.DIODE(_05667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11053__A0 (.DIODE(_05667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11019__A0 (.DIODE(_05667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__A0 (.DIODE(_05667_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11521__A0 (.DIODE(_05669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11486__A0 (.DIODE(_05669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__A0 (.DIODE(_05669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11348__A0 (.DIODE(_05669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11313__A0 (.DIODE(_05669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11244__A0 (.DIODE(_05669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11090__A0 (.DIODE(_05669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11055__A0 (.DIODE(_05669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11021__A0 (.DIODE(_05669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10946__A0 (.DIODE(_05669_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11523__A0 (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11488__A0 (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11385__A0 (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11350__A0 (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11315__A0 (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11246__A0 (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11092__A0 (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11057__A0 (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11023__A0 (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10949__A0 (.DIODE(_05671_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11525__A0 (.DIODE(_05673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11490__A0 (.DIODE(_05673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11387__A0 (.DIODE(_05673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11352__A0 (.DIODE(_05673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11317__A0 (.DIODE(_05673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11248__A0 (.DIODE(_05673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11094__A0 (.DIODE(_05673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11059__A0 (.DIODE(_05673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11025__A0 (.DIODE(_05673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10952__A0 (.DIODE(_05673_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11527__A0 (.DIODE(_05675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11492__A0 (.DIODE(_05675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11389__A0 (.DIODE(_05675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11354__A0 (.DIODE(_05675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11319__A0 (.DIODE(_05675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11250__A0 (.DIODE(_05675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11096__A0 (.DIODE(_05675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11061__A0 (.DIODE(_05675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11027__A0 (.DIODE(_05675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__A0 (.DIODE(_05675_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11529__A0 (.DIODE(_05677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11494__A0 (.DIODE(_05677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11391__A0 (.DIODE(_05677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11356__A0 (.DIODE(_05677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11321__A0 (.DIODE(_05677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11252__A0 (.DIODE(_05677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11098__A0 (.DIODE(_05677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11063__A0 (.DIODE(_05677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11029__A0 (.DIODE(_05677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10958__A0 (.DIODE(_05677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11531__A0 (.DIODE(_05679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__A0 (.DIODE(_05679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11393__A0 (.DIODE(_05679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11358__A0 (.DIODE(_05679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11323__A0 (.DIODE(_05679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11254__A0 (.DIODE(_05679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11100__A0 (.DIODE(_05679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11065__A0 (.DIODE(_05679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11031__A0 (.DIODE(_05679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10961__A0 (.DIODE(_05679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11533__A0 (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11498__A0 (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11395__A0 (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11360__A0 (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11325__A0 (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11256__A0 (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11102__A0 (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11067__A0 (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11033__A0 (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10964__A0 (.DIODE(_05681_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10998__S (.DIODE(_05683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10996__S (.DIODE(_05683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10994__S (.DIODE(_05683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10992__S (.DIODE(_05683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10990__S (.DIODE(_05683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10988__S (.DIODE(_05683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10967__A (.DIODE(_05683_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10986__S (.DIODE(_05684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10984__S (.DIODE(_05684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10982__S (.DIODE(_05684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__S (.DIODE(_05684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10978__S (.DIODE(_05684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10976__S (.DIODE(_05684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10974__S (.DIODE(_05684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10972__S (.DIODE(_05684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10970__S (.DIODE(_05684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10968__S (.DIODE(_05684_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11021__S (.DIODE(_05703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11019__S (.DIODE(_05703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11017__S (.DIODE(_05703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11015__S (.DIODE(_05703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11013__S (.DIODE(_05703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11011__S (.DIODE(_05703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11009__S (.DIODE(_05703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11007__S (.DIODE(_05703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11005__S (.DIODE(_05703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11003__S (.DIODE(_05703_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11067__S (.DIODE(_05720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11065__S (.DIODE(_05720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11063__S (.DIODE(_05720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11061__S (.DIODE(_05720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11059__S (.DIODE(_05720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11057__S (.DIODE(_05720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__A (.DIODE(_05720_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11055__S (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11053__S (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11051__S (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11049__S (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11047__S (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11045__S (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11043__S (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__S (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11039__S (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11037__S (.DIODE(_05721_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11102__S (.DIODE(_05739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11100__S (.DIODE(_05739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11098__S (.DIODE(_05739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11096__S (.DIODE(_05739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11094__S (.DIODE(_05739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11092__S (.DIODE(_05739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11071__A (.DIODE(_05739_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11090__S (.DIODE(_05740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11088__S (.DIODE(_05740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11086__S (.DIODE(_05740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11084__S (.DIODE(_05740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11082__S (.DIODE(_05740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11080__S (.DIODE(_05740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11078__S (.DIODE(_05740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11076__S (.DIODE(_05740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11074__S (.DIODE(_05740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11072__S (.DIODE(_05740_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11137__S (.DIODE(_05758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11135__S (.DIODE(_05758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11133__S (.DIODE(_05758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11131__S (.DIODE(_05758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11129__S (.DIODE(_05758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11127__S (.DIODE(_05758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11106__A (.DIODE(_05758_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11125__S (.DIODE(_05759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11123__S (.DIODE(_05759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11121__S (.DIODE(_05759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11119__S (.DIODE(_05759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11117__S (.DIODE(_05759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11115__S (.DIODE(_05759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11113__S (.DIODE(_05759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11111__S (.DIODE(_05759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11109__S (.DIODE(_05759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11107__S (.DIODE(_05759_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11828__A1 (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11794__A1 (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11760__A1 (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11726__A1 (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__A1 (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11433__A1 (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11399__A1 (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__A1 (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__A1 (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11142__A1 (.DIODE(_05776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11187__S (.DIODE(_05777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11184__S (.DIODE(_05777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11181__S (.DIODE(_05777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11178__S (.DIODE(_05777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11175__S (.DIODE(_05777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__S (.DIODE(_05777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11141__A (.DIODE(_05777_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11169__S (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__S (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11163__S (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11160__S (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11157__S (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__S (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11151__S (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11148__S (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11145__S (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11142__S (.DIODE(_05778_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11830__A1 (.DIODE(_05780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11796__A1 (.DIODE(_05780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11762__A1 (.DIODE(_05780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__A1 (.DIODE(_05780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11694__A1 (.DIODE(_05780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11435__A1 (.DIODE(_05780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11401__A1 (.DIODE(_05780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11262__A1 (.DIODE(_05780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11193__A1 (.DIODE(_05780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11145__A1 (.DIODE(_05780_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11832__A1 (.DIODE(_05782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11798__A1 (.DIODE(_05782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11764__A1 (.DIODE(_05782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11730__A1 (.DIODE(_05782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11696__A1 (.DIODE(_05782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11437__A1 (.DIODE(_05782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11403__A1 (.DIODE(_05782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11264__A1 (.DIODE(_05782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11195__A1 (.DIODE(_05782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11148__A1 (.DIODE(_05782_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11834__A1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11800__A1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11766__A1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11732__A1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11698__A1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11439__A1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11405__A1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11266__A1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11197__A1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11151__A1 (.DIODE(_05784_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11836__A1 (.DIODE(_05786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11802__A1 (.DIODE(_05786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11768__A1 (.DIODE(_05786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11734__A1 (.DIODE(_05786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11700__A1 (.DIODE(_05786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11441__A1 (.DIODE(_05786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11407__A1 (.DIODE(_05786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11268__A1 (.DIODE(_05786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11199__A1 (.DIODE(_05786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__A1 (.DIODE(_05786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11838__A1 (.DIODE(_05788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11804__A1 (.DIODE(_05788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11770__A1 (.DIODE(_05788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11736__A1 (.DIODE(_05788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11702__A1 (.DIODE(_05788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11443__A1 (.DIODE(_05788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11409__A1 (.DIODE(_05788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11270__A1 (.DIODE(_05788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11201__A1 (.DIODE(_05788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11157__A1 (.DIODE(_05788_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11840__A1 (.DIODE(_05790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11806__A1 (.DIODE(_05790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11772__A1 (.DIODE(_05790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11738__A1 (.DIODE(_05790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__A1 (.DIODE(_05790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11445__A1 (.DIODE(_05790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11411__A1 (.DIODE(_05790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__A1 (.DIODE(_05790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11203__A1 (.DIODE(_05790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11160__A1 (.DIODE(_05790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11842__A1 (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11808__A1 (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11774__A1 (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__A1 (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11706__A1 (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11447__A1 (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11413__A1 (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11274__A1 (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11205__A1 (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11163__A1 (.DIODE(_05792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11844__A1 (.DIODE(_05794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11810__A1 (.DIODE(_05794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11776__A1 (.DIODE(_05794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11742__A1 (.DIODE(_05794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11708__A1 (.DIODE(_05794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11449__A1 (.DIODE(_05794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11415__A1 (.DIODE(_05794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11276__A1 (.DIODE(_05794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11207__A1 (.DIODE(_05794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__A1 (.DIODE(_05794_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11846__A1 (.DIODE(_05796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11812__A1 (.DIODE(_05796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11778__A1 (.DIODE(_05796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11744__A1 (.DIODE(_05796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11710__A1 (.DIODE(_05796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11451__A1 (.DIODE(_05796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11417__A1 (.DIODE(_05796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11278__A1 (.DIODE(_05796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11209__A1 (.DIODE(_05796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11169__A1 (.DIODE(_05796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11848__A1 (.DIODE(_05798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11814__A1 (.DIODE(_05798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11780__A1 (.DIODE(_05798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11746__A1 (.DIODE(_05798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11712__A1 (.DIODE(_05798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11453__A1 (.DIODE(_05798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11419__A1 (.DIODE(_05798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__A1 (.DIODE(_05798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11211__A1 (.DIODE(_05798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__A1 (.DIODE(_05798_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11850__A1 (.DIODE(_05800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11816__A1 (.DIODE(_05800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11782__A1 (.DIODE(_05800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11748__A1 (.DIODE(_05800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11714__A1 (.DIODE(_05800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11455__A1 (.DIODE(_05800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11421__A1 (.DIODE(_05800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11282__A1 (.DIODE(_05800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11213__A1 (.DIODE(_05800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11175__A1 (.DIODE(_05800_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11852__A1 (.DIODE(_05802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11818__A1 (.DIODE(_05802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11784__A1 (.DIODE(_05802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11750__A1 (.DIODE(_05802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11716__A1 (.DIODE(_05802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11457__A1 (.DIODE(_05802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11423__A1 (.DIODE(_05802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11284__A1 (.DIODE(_05802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11215__A1 (.DIODE(_05802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11178__A1 (.DIODE(_05802_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11854__A1 (.DIODE(_05804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11820__A1 (.DIODE(_05804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11786__A1 (.DIODE(_05804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11752__A1 (.DIODE(_05804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11718__A1 (.DIODE(_05804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11459__A1 (.DIODE(_05804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11425__A1 (.DIODE(_05804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11286__A1 (.DIODE(_05804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11217__A1 (.DIODE(_05804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11181__A1 (.DIODE(_05804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11856__A1 (.DIODE(_05806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11822__A1 (.DIODE(_05806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11788__A1 (.DIODE(_05806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11754__A1 (.DIODE(_05806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__A1 (.DIODE(_05806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11461__A1 (.DIODE(_05806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11427__A1 (.DIODE(_05806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11288__A1 (.DIODE(_05806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11219__A1 (.DIODE(_05806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11184__A1 (.DIODE(_05806_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11858__A1 (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11824__A1 (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11790__A1 (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__A1 (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11722__A1 (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11463__A1 (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11429__A1 (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11290__A1 (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11221__A1 (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11187__A1 (.DIODE(_05808_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11221__S (.DIODE(_05810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11219__S (.DIODE(_05810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11217__S (.DIODE(_05810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11215__S (.DIODE(_05810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11213__S (.DIODE(_05810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11211__S (.DIODE(_05810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11190__A (.DIODE(_05810_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11209__S (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11207__S (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11205__S (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11203__S (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11201__S (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11199__S (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11197__S (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11195__S (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11193__S (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__S (.DIODE(_05811_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11256__S (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11254__S (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11252__S (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11250__S (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11248__S (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11246__S (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__A (.DIODE(_05829_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11244__S (.DIODE(_05830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11242__S (.DIODE(_05830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11240__S (.DIODE(_05830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11238__S (.DIODE(_05830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11236__S (.DIODE(_05830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11234__S (.DIODE(_05830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11232__S (.DIODE(_05830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11230__S (.DIODE(_05830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11228__S (.DIODE(_05830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11226__S (.DIODE(_05830_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11290__S (.DIODE(_05847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11288__S (.DIODE(_05847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11286__S (.DIODE(_05847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11284__S (.DIODE(_05847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11282__S (.DIODE(_05847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__S (.DIODE(_05847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11259__A (.DIODE(_05847_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11278__S (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11276__S (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11274__S (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__S (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11270__S (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11268__S (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11266__S (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11264__S (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11262__S (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__S (.DIODE(_05848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11325__S (.DIODE(_05866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11323__S (.DIODE(_05866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11321__S (.DIODE(_05866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11319__S (.DIODE(_05866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11317__S (.DIODE(_05866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11315__S (.DIODE(_05866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11294__A (.DIODE(_05866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11313__S (.DIODE(_05867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11311__S (.DIODE(_05867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11309__S (.DIODE(_05867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11307__S (.DIODE(_05867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11305__S (.DIODE(_05867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11303__S (.DIODE(_05867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11301__S (.DIODE(_05867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11299__S (.DIODE(_05867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11297__S (.DIODE(_05867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11295__S (.DIODE(_05867_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11360__S (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11358__S (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11356__S (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11354__S (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11352__S (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11350__S (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11329__A (.DIODE(_05885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11348__S (.DIODE(_05886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11346__S (.DIODE(_05886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11344__S (.DIODE(_05886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11342__S (.DIODE(_05886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11340__S (.DIODE(_05886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11338__S (.DIODE(_05886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11336__S (.DIODE(_05886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11334__S (.DIODE(_05886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11332__S (.DIODE(_05886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11330__S (.DIODE(_05886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11395__S (.DIODE(_05904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11393__S (.DIODE(_05904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11391__S (.DIODE(_05904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11389__S (.DIODE(_05904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11387__S (.DIODE(_05904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11385__S (.DIODE(_05904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11364__A (.DIODE(_05904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11383__S (.DIODE(_05905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11381__S (.DIODE(_05905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11379__S (.DIODE(_05905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11377__S (.DIODE(_05905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11375__S (.DIODE(_05905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11373__S (.DIODE(_05905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11371__S (.DIODE(_05905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11369__S (.DIODE(_05905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11367__S (.DIODE(_05905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11365__S (.DIODE(_05905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11429__S (.DIODE(_05922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11427__S (.DIODE(_05922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11425__S (.DIODE(_05922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11423__S (.DIODE(_05922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11421__S (.DIODE(_05922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11419__S (.DIODE(_05922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11398__A (.DIODE(_05922_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11417__S (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11415__S (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11413__S (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11411__S (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11409__S (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11407__S (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11405__S (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11403__S (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11401__S (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11399__S (.DIODE(_05923_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11451__S (.DIODE(_05941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11449__S (.DIODE(_05941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11447__S (.DIODE(_05941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11445__S (.DIODE(_05941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11443__S (.DIODE(_05941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11441__S (.DIODE(_05941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11439__S (.DIODE(_05941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11437__S (.DIODE(_05941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11435__S (.DIODE(_05941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11433__S (.DIODE(_05941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11498__S (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__S (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11494__S (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11492__S (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11490__S (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11488__S (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11467__A (.DIODE(_05959_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11486__S (.DIODE(_05960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11484__S (.DIODE(_05960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11482__S (.DIODE(_05960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11480__S (.DIODE(_05960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11478__S (.DIODE(_05960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__S (.DIODE(_05960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11474__S (.DIODE(_05960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11472__S (.DIODE(_05960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11470__S (.DIODE(_05960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11468__S (.DIODE(_05960_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11533__S (.DIODE(_05978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11531__S (.DIODE(_05978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11529__S (.DIODE(_05978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11527__S (.DIODE(_05978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11525__S (.DIODE(_05978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11523__S (.DIODE(_05978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11502__A (.DIODE(_05978_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11521__S (.DIODE(_05979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11519__S (.DIODE(_05979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__S (.DIODE(_05979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11515__S (.DIODE(_05979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11513__S (.DIODE(_05979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11511__S (.DIODE(_05979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11509__S (.DIODE(_05979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11507__S (.DIODE(_05979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11505__S (.DIODE(_05979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11503__S (.DIODE(_05979_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12072__A0 (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12037__A0 (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12002__A0 (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11933__A0 (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11898__A0 (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__A0 (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11658__A0 (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11623__A0 (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11589__A0 (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11539__A0 (.DIODE(_05996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11584__S (.DIODE(_05998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11581__S (.DIODE(_05998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11578__S (.DIODE(_05998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11575__S (.DIODE(_05998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11572__S (.DIODE(_05998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11569__S (.DIODE(_05998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11538__A (.DIODE(_05998_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11566__S (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__S (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11560__S (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11557__S (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11554__S (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11551__S (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11548__S (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11545__S (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11542__S (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11539__S (.DIODE(_05999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12074__A0 (.DIODE(_06001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12039__A0 (.DIODE(_06001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__A0 (.DIODE(_06001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11935__A0 (.DIODE(_06001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11900__A0 (.DIODE(_06001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11865__A0 (.DIODE(_06001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11660__A0 (.DIODE(_06001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11625__A0 (.DIODE(_06001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11591__A0 (.DIODE(_06001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11542__A0 (.DIODE(_06001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12076__A0 (.DIODE(_06003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12041__A0 (.DIODE(_06003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__A0 (.DIODE(_06003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11937__A0 (.DIODE(_06003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11902__A0 (.DIODE(_06003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__A0 (.DIODE(_06003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11662__A0 (.DIODE(_06003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11627__A0 (.DIODE(_06003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11593__A0 (.DIODE(_06003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11545__A0 (.DIODE(_06003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12078__A0 (.DIODE(_06005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12043__A0 (.DIODE(_06005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12008__A0 (.DIODE(_06005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11939__A0 (.DIODE(_06005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11904__A0 (.DIODE(_06005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11869__A0 (.DIODE(_06005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11664__A0 (.DIODE(_06005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11629__A0 (.DIODE(_06005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11595__A0 (.DIODE(_06005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11548__A0 (.DIODE(_06005_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12080__A0 (.DIODE(_06007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12045__A0 (.DIODE(_06007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12010__A0 (.DIODE(_06007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11941__A0 (.DIODE(_06007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11906__A0 (.DIODE(_06007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11871__A0 (.DIODE(_06007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11666__A0 (.DIODE(_06007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11631__A0 (.DIODE(_06007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11597__A0 (.DIODE(_06007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11551__A0 (.DIODE(_06007_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12082__A0 (.DIODE(_06009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12047__A0 (.DIODE(_06009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12012__A0 (.DIODE(_06009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11943__A0 (.DIODE(_06009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11908__A0 (.DIODE(_06009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11873__A0 (.DIODE(_06009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11668__A0 (.DIODE(_06009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11633__A0 (.DIODE(_06009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11599__A0 (.DIODE(_06009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11554__A0 (.DIODE(_06009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12084__A0 (.DIODE(_06011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12049__A0 (.DIODE(_06011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12014__A0 (.DIODE(_06011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11945__A0 (.DIODE(_06011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11910__A0 (.DIODE(_06011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11875__A0 (.DIODE(_06011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__A0 (.DIODE(_06011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11635__A0 (.DIODE(_06011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11601__A0 (.DIODE(_06011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11557__A0 (.DIODE(_06011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12086__A0 (.DIODE(_06013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12051__A0 (.DIODE(_06013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12016__A0 (.DIODE(_06013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11947__A0 (.DIODE(_06013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11912__A0 (.DIODE(_06013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11877__A0 (.DIODE(_06013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11672__A0 (.DIODE(_06013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__A0 (.DIODE(_06013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11603__A0 (.DIODE(_06013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11560__A0 (.DIODE(_06013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12088__A0 (.DIODE(_06015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12053__A0 (.DIODE(_06015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12018__A0 (.DIODE(_06015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11949__A0 (.DIODE(_06015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11914__A0 (.DIODE(_06015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11879__A0 (.DIODE(_06015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11674__A0 (.DIODE(_06015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__A0 (.DIODE(_06015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11605__A0 (.DIODE(_06015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__A0 (.DIODE(_06015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12090__A0 (.DIODE(_06017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12055__A0 (.DIODE(_06017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12020__A0 (.DIODE(_06017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11951__A0 (.DIODE(_06017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11916__A0 (.DIODE(_06017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11881__A0 (.DIODE(_06017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11676__A0 (.DIODE(_06017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11641__A0 (.DIODE(_06017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11607__A0 (.DIODE(_06017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11566__A0 (.DIODE(_06017_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12092__A0 (.DIODE(_06019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12057__A0 (.DIODE(_06019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12022__A0 (.DIODE(_06019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__A0 (.DIODE(_06019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11918__A0 (.DIODE(_06019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11883__A0 (.DIODE(_06019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11678__A0 (.DIODE(_06019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11643__A0 (.DIODE(_06019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11609__A0 (.DIODE(_06019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11569__A0 (.DIODE(_06019_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12094__A0 (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12059__A0 (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12024__A0 (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11955__A0 (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11920__A0 (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11885__A0 (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11680__A0 (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11645__A0 (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11611__A0 (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11572__A0 (.DIODE(_06021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12096__A0 (.DIODE(_06023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12061__A0 (.DIODE(_06023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12026__A0 (.DIODE(_06023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11957__A0 (.DIODE(_06023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11922__A0 (.DIODE(_06023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11887__A0 (.DIODE(_06023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11682__A0 (.DIODE(_06023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11647__A0 (.DIODE(_06023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11613__A0 (.DIODE(_06023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11575__A0 (.DIODE(_06023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12098__A0 (.DIODE(_06025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12063__A0 (.DIODE(_06025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12028__A0 (.DIODE(_06025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11959__A0 (.DIODE(_06025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11924__A0 (.DIODE(_06025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11889__A0 (.DIODE(_06025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11684__A0 (.DIODE(_06025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11649__A0 (.DIODE(_06025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11615__A0 (.DIODE(_06025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11578__A0 (.DIODE(_06025_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12100__A0 (.DIODE(_06027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12065__A0 (.DIODE(_06027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12030__A0 (.DIODE(_06027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11961__A0 (.DIODE(_06027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11926__A0 (.DIODE(_06027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11891__A0 (.DIODE(_06027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11686__A0 (.DIODE(_06027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11651__A0 (.DIODE(_06027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11617__A0 (.DIODE(_06027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11581__A0 (.DIODE(_06027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12102__A0 (.DIODE(_06029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12067__A0 (.DIODE(_06029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12032__A0 (.DIODE(_06029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11963__A0 (.DIODE(_06029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11928__A0 (.DIODE(_06029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11893__A0 (.DIODE(_06029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11688__A0 (.DIODE(_06029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11653__A0 (.DIODE(_06029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11619__A0 (.DIODE(_06029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11584__A0 (.DIODE(_06029_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11619__S (.DIODE(_06032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11617__S (.DIODE(_06032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11615__S (.DIODE(_06032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11613__S (.DIODE(_06032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11611__S (.DIODE(_06032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11609__S (.DIODE(_06032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11588__A (.DIODE(_06032_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11607__S (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11605__S (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11603__S (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11601__S (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11599__S (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11597__S (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11595__S (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11593__S (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11591__S (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11589__S (.DIODE(_06033_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11653__S (.DIODE(_06050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11651__S (.DIODE(_06050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11649__S (.DIODE(_06050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11647__S (.DIODE(_06050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11645__S (.DIODE(_06050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11643__S (.DIODE(_06050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11622__A (.DIODE(_06050_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11641__S (.DIODE(_06051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11639__S (.DIODE(_06051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__S (.DIODE(_06051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11635__S (.DIODE(_06051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11633__S (.DIODE(_06051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11631__S (.DIODE(_06051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11629__S (.DIODE(_06051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11627__S (.DIODE(_06051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11625__S (.DIODE(_06051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11623__S (.DIODE(_06051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11688__S (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11686__S (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11684__S (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11682__S (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11680__S (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11678__S (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11657__A (.DIODE(_06069_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11676__S (.DIODE(_06070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11674__S (.DIODE(_06070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11672__S (.DIODE(_06070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__S (.DIODE(_06070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11668__S (.DIODE(_06070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11666__S (.DIODE(_06070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11664__S (.DIODE(_06070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11662__S (.DIODE(_06070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11660__S (.DIODE(_06070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11658__S (.DIODE(_06070_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11722__S (.DIODE(_06087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__S (.DIODE(_06087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11718__S (.DIODE(_06087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11716__S (.DIODE(_06087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11714__S (.DIODE(_06087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11712__S (.DIODE(_06087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11691__A (.DIODE(_06087_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11710__S (.DIODE(_06088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11708__S (.DIODE(_06088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11706__S (.DIODE(_06088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__S (.DIODE(_06088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11702__S (.DIODE(_06088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11700__S (.DIODE(_06088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11698__S (.DIODE(_06088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11696__S (.DIODE(_06088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11694__S (.DIODE(_06088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11692__S (.DIODE(_06088_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__S (.DIODE(_06105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11754__S (.DIODE(_06105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11752__S (.DIODE(_06105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11750__S (.DIODE(_06105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11748__S (.DIODE(_06105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11746__S (.DIODE(_06105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11725__A (.DIODE(_06105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11744__S (.DIODE(_06106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11742__S (.DIODE(_06106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__S (.DIODE(_06106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11738__S (.DIODE(_06106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11736__S (.DIODE(_06106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11734__S (.DIODE(_06106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11732__S (.DIODE(_06106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11730__S (.DIODE(_06106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11728__S (.DIODE(_06106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11726__S (.DIODE(_06106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11790__S (.DIODE(_06123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11788__S (.DIODE(_06123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11786__S (.DIODE(_06123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11784__S (.DIODE(_06123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11782__S (.DIODE(_06123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11780__S (.DIODE(_06123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11759__A (.DIODE(_06123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11778__S (.DIODE(_06124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11776__S (.DIODE(_06124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11774__S (.DIODE(_06124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11772__S (.DIODE(_06124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11770__S (.DIODE(_06124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11768__S (.DIODE(_06124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11766__S (.DIODE(_06124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11764__S (.DIODE(_06124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11762__S (.DIODE(_06124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11760__S (.DIODE(_06124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11812__S (.DIODE(_06142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11810__S (.DIODE(_06142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11808__S (.DIODE(_06142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11806__S (.DIODE(_06142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11804__S (.DIODE(_06142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11802__S (.DIODE(_06142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11800__S (.DIODE(_06142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11798__S (.DIODE(_06142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11796__S (.DIODE(_06142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11794__S (.DIODE(_06142_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11858__S (.DIODE(_06159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11856__S (.DIODE(_06159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11854__S (.DIODE(_06159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11852__S (.DIODE(_06159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11850__S (.DIODE(_06159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11848__S (.DIODE(_06159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11827__A (.DIODE(_06159_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11846__S (.DIODE(_06160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11844__S (.DIODE(_06160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11842__S (.DIODE(_06160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11840__S (.DIODE(_06160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11838__S (.DIODE(_06160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11836__S (.DIODE(_06160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11834__S (.DIODE(_06160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11832__S (.DIODE(_06160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11830__S (.DIODE(_06160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11828__S (.DIODE(_06160_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11893__S (.DIODE(_06178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11891__S (.DIODE(_06178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11889__S (.DIODE(_06178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11887__S (.DIODE(_06178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11885__S (.DIODE(_06178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11883__S (.DIODE(_06178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11862__A (.DIODE(_06178_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11881__S (.DIODE(_06179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11879__S (.DIODE(_06179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11877__S (.DIODE(_06179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11875__S (.DIODE(_06179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11873__S (.DIODE(_06179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11871__S (.DIODE(_06179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11869__S (.DIODE(_06179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11867__S (.DIODE(_06179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11865__S (.DIODE(_06179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__S (.DIODE(_06179_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11928__S (.DIODE(_06197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11926__S (.DIODE(_06197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11924__S (.DIODE(_06197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11922__S (.DIODE(_06197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11920__S (.DIODE(_06197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11918__S (.DIODE(_06197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11897__A (.DIODE(_06197_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11916__S (.DIODE(_06198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11914__S (.DIODE(_06198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11912__S (.DIODE(_06198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11910__S (.DIODE(_06198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11908__S (.DIODE(_06198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11906__S (.DIODE(_06198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11904__S (.DIODE(_06198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11902__S (.DIODE(_06198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11900__S (.DIODE(_06198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11898__S (.DIODE(_06198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11963__S (.DIODE(_06216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11961__S (.DIODE(_06216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11959__S (.DIODE(_06216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11957__S (.DIODE(_06216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11955__S (.DIODE(_06216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11953__S (.DIODE(_06216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11932__A (.DIODE(_06216_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11951__S (.DIODE(_06217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11949__S (.DIODE(_06217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11947__S (.DIODE(_06217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11945__S (.DIODE(_06217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11943__S (.DIODE(_06217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11941__S (.DIODE(_06217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11939__S (.DIODE(_06217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11937__S (.DIODE(_06217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11935__S (.DIODE(_06217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11933__S (.DIODE(_06217_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11985__S (.DIODE(_06235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11983__S (.DIODE(_06235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11981__S (.DIODE(_06235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11979__S (.DIODE(_06235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11977__S (.DIODE(_06235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11975__S (.DIODE(_06235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11973__S (.DIODE(_06235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11971__S (.DIODE(_06235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11969__S (.DIODE(_06235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11967__S (.DIODE(_06235_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12020__S (.DIODE(_06254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12018__S (.DIODE(_06254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12016__S (.DIODE(_06254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12014__S (.DIODE(_06254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12012__S (.DIODE(_06254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12010__S (.DIODE(_06254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12008__S (.DIODE(_06254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__S (.DIODE(_06254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__S (.DIODE(_06254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12002__S (.DIODE(_06254_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12055__S (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12053__S (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12051__S (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12049__S (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12047__S (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12045__S (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12043__S (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12041__S (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12039__S (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12037__S (.DIODE(_06273_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12102__S (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12100__S (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12098__S (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12096__S (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12094__S (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12092__S (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12071__A (.DIODE(_06291_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12090__S (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12088__S (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12086__S (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12084__S (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12082__S (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12080__S (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12078__S (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12076__S (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12074__S (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12072__S (.DIODE(_06292_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12642__A0 (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12607__A0 (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12572__A0 (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12503__A0 (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12468__A0 (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12433__A0 (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12364__A0 (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12226__A0 (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12191__A0 (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12108__A0 (.DIODE(_06309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12135__S (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12132__S (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12129__S (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12126__S (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12123__S (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12120__S (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12117__S (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12114__S (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12111__S (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12108__S (.DIODE(_06312_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12644__A0 (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12609__A0 (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12574__A0 (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12505__A0 (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12470__A0 (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12435__A0 (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12366__A0 (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12228__A0 (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12193__A0 (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12111__A0 (.DIODE(_06314_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12646__A0 (.DIODE(_06316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12611__A0 (.DIODE(_06316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12576__A0 (.DIODE(_06316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12507__A0 (.DIODE(_06316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12472__A0 (.DIODE(_06316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12437__A0 (.DIODE(_06316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12368__A0 (.DIODE(_06316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12230__A0 (.DIODE(_06316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12195__A0 (.DIODE(_06316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12114__A0 (.DIODE(_06316_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12648__A0 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12613__A0 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12578__A0 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12509__A0 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12474__A0 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12439__A0 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12370__A0 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12232__A0 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12197__A0 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12117__A0 (.DIODE(_06318_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12650__A0 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12615__A0 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12580__A0 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12511__A0 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12476__A0 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12441__A0 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12372__A0 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12234__A0 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12199__A0 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12120__A0 (.DIODE(_06320_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12652__A0 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12617__A0 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12582__A0 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12513__A0 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12478__A0 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12443__A0 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12374__A0 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12236__A0 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12201__A0 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12123__A0 (.DIODE(_06322_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12654__A0 (.DIODE(_06324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12619__A0 (.DIODE(_06324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12584__A0 (.DIODE(_06324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12515__A0 (.DIODE(_06324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12480__A0 (.DIODE(_06324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12445__A0 (.DIODE(_06324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12376__A0 (.DIODE(_06324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12238__A0 (.DIODE(_06324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12203__A0 (.DIODE(_06324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12126__A0 (.DIODE(_06324_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12656__A0 (.DIODE(_06326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12621__A0 (.DIODE(_06326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12586__A0 (.DIODE(_06326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12517__A0 (.DIODE(_06326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12482__A0 (.DIODE(_06326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12447__A0 (.DIODE(_06326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12378__A0 (.DIODE(_06326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12240__A0 (.DIODE(_06326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12205__A0 (.DIODE(_06326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12129__A0 (.DIODE(_06326_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12658__A0 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12623__A0 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12588__A0 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12519__A0 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12484__A0 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12449__A0 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12380__A0 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12242__A0 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12207__A0 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12132__A0 (.DIODE(_06328_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12660__A0 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12625__A0 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12590__A0 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12521__A0 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12486__A0 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12451__A0 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12382__A0 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12244__A0 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12209__A0 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12135__A0 (.DIODE(_06330_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12662__A0 (.DIODE(_06332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12627__A0 (.DIODE(_06332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12592__A0 (.DIODE(_06332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12523__A0 (.DIODE(_06332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12488__A0 (.DIODE(_06332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12453__A0 (.DIODE(_06332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12384__A0 (.DIODE(_06332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12246__A0 (.DIODE(_06332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12211__A0 (.DIODE(_06332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12138__A0 (.DIODE(_06332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12664__A0 (.DIODE(_06334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12629__A0 (.DIODE(_06334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12594__A0 (.DIODE(_06334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12525__A0 (.DIODE(_06334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12490__A0 (.DIODE(_06334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12455__A0 (.DIODE(_06334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12386__A0 (.DIODE(_06334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12248__A0 (.DIODE(_06334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12213__A0 (.DIODE(_06334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12141__A0 (.DIODE(_06334_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12666__A0 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12631__A0 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12596__A0 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12527__A0 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12492__A0 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12457__A0 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12388__A0 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12250__A0 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12215__A0 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12144__A0 (.DIODE(_06336_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12668__A0 (.DIODE(_06338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12633__A0 (.DIODE(_06338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12598__A0 (.DIODE(_06338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12529__A0 (.DIODE(_06338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12494__A0 (.DIODE(_06338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12459__A0 (.DIODE(_06338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12390__A0 (.DIODE(_06338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__A0 (.DIODE(_06338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12217__A0 (.DIODE(_06338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12147__A0 (.DIODE(_06338_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12670__A0 (.DIODE(_06340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12635__A0 (.DIODE(_06340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12600__A0 (.DIODE(_06340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12531__A0 (.DIODE(_06340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12496__A0 (.DIODE(_06340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12461__A0 (.DIODE(_06340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12392__A0 (.DIODE(_06340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12254__A0 (.DIODE(_06340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12219__A0 (.DIODE(_06340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12150__A0 (.DIODE(_06340_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12672__A0 (.DIODE(_06342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12637__A0 (.DIODE(_06342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12602__A0 (.DIODE(_06342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12533__A0 (.DIODE(_06342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12498__A0 (.DIODE(_06342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12463__A0 (.DIODE(_06342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12394__A0 (.DIODE(_06342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12256__A0 (.DIODE(_06342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12221__A0 (.DIODE(_06342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12153__A0 (.DIODE(_06342_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12187__S (.DIODE(_06344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12185__S (.DIODE(_06344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12183__S (.DIODE(_06344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12181__S (.DIODE(_06344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12179__S (.DIODE(_06344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12177__S (.DIODE(_06344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12156__A (.DIODE(_06344_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12175__S (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12173__S (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12171__S (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12169__S (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12167__S (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12165__S (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12163__S (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12161__S (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12159__S (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12157__S (.DIODE(_06345_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12209__S (.DIODE(_06363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12207__S (.DIODE(_06363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12205__S (.DIODE(_06363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12203__S (.DIODE(_06363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12201__S (.DIODE(_06363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12199__S (.DIODE(_06363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12197__S (.DIODE(_06363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12195__S (.DIODE(_06363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12193__S (.DIODE(_06363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12191__S (.DIODE(_06363_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12256__S (.DIODE(_06381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12254__S (.DIODE(_06381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__S (.DIODE(_06381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12250__S (.DIODE(_06381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12248__S (.DIODE(_06381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12246__S (.DIODE(_06381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12225__A (.DIODE(_06381_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12244__S (.DIODE(_06382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12242__S (.DIODE(_06382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12240__S (.DIODE(_06382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12238__S (.DIODE(_06382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12236__S (.DIODE(_06382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12234__S (.DIODE(_06382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12232__S (.DIODE(_06382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12230__S (.DIODE(_06382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12228__S (.DIODE(_06382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12226__S (.DIODE(_06382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12291__S (.DIODE(_06400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12289__S (.DIODE(_06400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12287__S (.DIODE(_06400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12285__S (.DIODE(_06400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12283__S (.DIODE(_06400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__S (.DIODE(_06400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12260__A (.DIODE(_06400_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12279__S (.DIODE(_06401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12277__S (.DIODE(_06401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12275__S (.DIODE(_06401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12273__S (.DIODE(_06401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12271__S (.DIODE(_06401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12269__S (.DIODE(_06401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12267__S (.DIODE(_06401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12265__S (.DIODE(_06401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12263__S (.DIODE(_06401_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12261__S (.DIODE(_06401_));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(i_addr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(i_addr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(i_addr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(i_addr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(i_addr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(i_addr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(i_addr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_i_clk_A (.DIODE(i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(i_data[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(i_data[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(i_data[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(i_data[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(i_data[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(i_data[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(i_data[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(i_data[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(i_data[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(i_data[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(i_data[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(i_data[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(i_data[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(i_data[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(i_data[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(i_data[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(i_we));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2029_A (.DIODE(\mem[3][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06486__B2 (.DIODE(\mem[3][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2034_A (.DIODE(\mem[3][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07614__B2 (.DIODE(\mem[3][10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2040_A (.DIODE(\mem[3][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__B2 (.DIODE(\mem[3][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2047_A (.DIODE(\mem[3][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07973__B2 (.DIODE(\mem[3][14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2039_A (.DIODE(\mem[3][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08063__B2 (.DIODE(\mem[3][15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2042_A (.DIODE(\mem[49][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06544__A1 (.DIODE(\mem[49][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2044_A (.DIODE(\mem[49][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06889__A1 (.DIODE(\mem[49][2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2045_A (.DIODE(\mem[49][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06992__A1 (.DIODE(\mem[49][3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2048_A (.DIODE(\mem[49][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07090__A1 (.DIODE(\mem[49][4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2030_A (.DIODE(\mem[49][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__A1 (.DIODE(\mem[49][5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2037_A (.DIODE(\mem[49][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07270__A1 (.DIODE(\mem[49][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2046_A (.DIODE(\mem[49][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__A1 (.DIODE(\mem[49][7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2041_A (.DIODE(\mem[49][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07453__A1 (.DIODE(\mem[49][8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2033_A (.DIODE(\mem[5][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06502__A1 (.DIODE(\mem[5][0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2032_A (.DIODE(\mem[69][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06744__A1 (.DIODE(\mem[69][1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2036_A (.DIODE(\mem[71][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07892__B2 (.DIODE(\mem[71][13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2035_A (.DIODE(\mem[80][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07824__A1 (.DIODE(\mem[80][12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2043_A (.DIODE(\mem[85][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07291__A1 (.DIODE(\mem[85][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2038_A (.DIODE(\mem[86][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07290__A1 (.DIODE(\mem[86][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2031_A (.DIODE(\mem[87][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07290__B2 (.DIODE(\mem[87][6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06419__A_N (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06411__A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA__06439__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__06410__A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__06432__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__06415__A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA__06659__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__06556__B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__06548__A_N (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__06545__B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__06534__B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__06529__A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__06466__A_N (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__06447__B_N (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__06433__B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__06415__B (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__08625__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__08480__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__08140__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__06471__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__06408__A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA__08625__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__08300__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__08212__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__08140__B (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__06560__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__06406__A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA__08211__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__08141__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__06685__A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA__08853__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA__08901__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__08188__A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA__08909__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__08196__A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA__08861__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__08148__A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA__08865__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__08152__A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA__08869__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__08156__A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__08873__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__08160__A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__08877__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__08164__A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__08881__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__08168__A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__08172__A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__08889__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__08176__A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__08893__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__08180__A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA__08211__B (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__08141__B_N (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_output25_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_output26_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_output27_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_output28_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_output29_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_output30_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_output31_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_output32_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_output33_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_output34_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_output35_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_output36_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_output37_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_output38_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_output39_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_output40_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_1_0_i_clk_A (.DIODE(clknet_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_1_0_0_i_clk_A (.DIODE(clknet_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1_0_i_clk_A (.DIODE(clknet_1_0_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0_0_i_clk_A (.DIODE(clknet_1_0_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3_0_i_clk_A (.DIODE(clknet_1_1_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2_0_i_clk_A (.DIODE(clknet_1_1_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1_0_i_clk_A (.DIODE(clknet_2_0_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0_0_i_clk_A (.DIODE(clknet_2_0_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3_0_i_clk_A (.DIODE(clknet_2_1_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2_0_i_clk_A (.DIODE(clknet_2_1_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5_0_i_clk_A (.DIODE(clknet_2_2_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4_0_i_clk_A (.DIODE(clknet_2_2_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7_0_i_clk_A (.DIODE(clknet_2_3_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6_0_i_clk_A (.DIODE(clknet_2_3_1_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1_0_i_clk_A (.DIODE(clknet_3_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0_0_i_clk_A (.DIODE(clknet_3_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3_0_i_clk_A (.DIODE(clknet_3_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2_0_i_clk_A (.DIODE(clknet_3_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5_0_i_clk_A (.DIODE(clknet_3_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4_0_i_clk_A (.DIODE(clknet_3_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7_0_i_clk_A (.DIODE(clknet_3_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6_0_i_clk_A (.DIODE(clknet_3_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9_0_i_clk_A (.DIODE(clknet_3_4_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8_0_i_clk_A (.DIODE(clknet_3_4_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11_0_i_clk_A (.DIODE(clknet_3_5_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10_0_i_clk_A (.DIODE(clknet_3_5_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13_0_i_clk_A (.DIODE(clknet_3_6_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12_0_i_clk_A (.DIODE(clknet_3_6_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15_0_i_clk_A (.DIODE(clknet_3_7_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14_0_i_clk_A (.DIODE(clknet_3_7_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_288_i_clk_A (.DIODE(clknet_5_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_287_i_clk_A (.DIODE(clknet_5_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_i_clk_A (.DIODE(clknet_5_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_i_clk_A (.DIODE(clknet_5_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_i_clk_A (.DIODE(clknet_5_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_i_clk_A (.DIODE(clknet_5_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_i_clk_A (.DIODE(clknet_5_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_i_clk_A (.DIODE(clknet_5_0_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_286_i_clk_A (.DIODE(clknet_5_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_285_i_clk_A (.DIODE(clknet_5_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_284_i_clk_A (.DIODE(clknet_5_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_283_i_clk_A (.DIODE(clknet_5_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_282_i_clk_A (.DIODE(clknet_5_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_281_i_clk_A (.DIODE(clknet_5_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_280_i_clk_A (.DIODE(clknet_5_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_i_clk_A (.DIODE(clknet_5_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_i_clk_A (.DIODE(clknet_5_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_i_clk_A (.DIODE(clknet_5_1_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_i_clk_A (.DIODE(clknet_5_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_i_clk_A (.DIODE(clknet_5_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_i_clk_A (.DIODE(clknet_5_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_i_clk_A (.DIODE(clknet_5_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_i_clk_A (.DIODE(clknet_5_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_i_clk_A (.DIODE(clknet_5_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_i_clk_A (.DIODE(clknet_5_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_i_clk_A (.DIODE(clknet_5_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_i_clk_A (.DIODE(clknet_5_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_i_clk_A (.DIODE(clknet_5_2_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_i_clk_A (.DIODE(clknet_5_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_i_clk_A (.DIODE(clknet_5_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_i_clk_A (.DIODE(clknet_5_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_i_clk_A (.DIODE(clknet_5_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_i_clk_A (.DIODE(clknet_5_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_i_clk_A (.DIODE(clknet_5_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_i_clk_A (.DIODE(clknet_5_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_i_clk_A (.DIODE(clknet_5_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_i_clk_A (.DIODE(clknet_5_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_i_clk_A (.DIODE(clknet_5_3_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_279_i_clk_A (.DIODE(clknet_5_4_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_278_i_clk_A (.DIODE(clknet_5_4_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_277_i_clk_A (.DIODE(clknet_5_4_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_276_i_clk_A (.DIODE(clknet_5_4_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_275_i_clk_A (.DIODE(clknet_5_4_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_274_i_clk_A (.DIODE(clknet_5_4_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_273_i_clk_A (.DIODE(clknet_5_4_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_263_i_clk_A (.DIODE(clknet_5_4_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_262_i_clk_A (.DIODE(clknet_5_4_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_272_i_clk_A (.DIODE(clknet_5_5_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_271_i_clk_A (.DIODE(clknet_5_5_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_270_i_clk_A (.DIODE(clknet_5_5_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_269_i_clk_A (.DIODE(clknet_5_5_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_268_i_clk_A (.DIODE(clknet_5_5_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_267_i_clk_A (.DIODE(clknet_5_5_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_266_i_clk_A (.DIODE(clknet_5_5_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_265_i_clk_A (.DIODE(clknet_5_5_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_264_i_clk_A (.DIODE(clknet_5_5_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_261_i_clk_A (.DIODE(clknet_5_6_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_260_i_clk_A (.DIODE(clknet_5_6_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_i_clk_A (.DIODE(clknet_5_6_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_i_clk_A (.DIODE(clknet_5_6_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_i_clk_A (.DIODE(clknet_5_6_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_i_clk_A (.DIODE(clknet_5_6_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_i_clk_A (.DIODE(clknet_5_6_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_i_clk_A (.DIODE(clknet_5_6_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_i_clk_A (.DIODE(clknet_5_6_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_259_i_clk_A (.DIODE(clknet_5_7_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_258_i_clk_A (.DIODE(clknet_5_7_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_257_i_clk_A (.DIODE(clknet_5_7_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_256_i_clk_A (.DIODE(clknet_5_7_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_255_i_clk_A (.DIODE(clknet_5_7_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_254_i_clk_A (.DIODE(clknet_5_7_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_253_i_clk_A (.DIODE(clknet_5_7_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_252_i_clk_A (.DIODE(clknet_5_7_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_i_clk_A (.DIODE(clknet_5_7_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_i_clk_A (.DIODE(clknet_5_7_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_i_clk_A (.DIODE(clknet_5_7_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_65_i_clk_A (.DIODE(clknet_5_8_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_64_i_clk_A (.DIODE(clknet_5_8_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_i_clk_A (.DIODE(clknet_5_8_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_i_clk_A (.DIODE(clknet_5_8_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_61_i_clk_A (.DIODE(clknet_5_8_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_i_clk_A (.DIODE(clknet_5_8_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_i_clk_A (.DIODE(clknet_5_8_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_i_clk_A (.DIODE(clknet_5_8_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_i_clk_A (.DIODE(clknet_5_8_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_i_clk_A (.DIODE(clknet_5_8_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_i_clk_A (.DIODE(clknet_5_8_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_69_i_clk_A (.DIODE(clknet_5_9_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_68_i_clk_A (.DIODE(clknet_5_9_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_i_clk_A (.DIODE(clknet_5_9_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_i_clk_A (.DIODE(clknet_5_9_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_i_clk_A (.DIODE(clknet_5_9_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_i_clk_A (.DIODE(clknet_5_9_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_52_i_clk_A (.DIODE(clknet_5_9_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_i_clk_A (.DIODE(clknet_5_9_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_50_i_clk_A (.DIODE(clknet_5_9_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_i_clk_A (.DIODE(clknet_5_9_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_i_clk_A (.DIODE(clknet_5_9_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_78_i_clk_A (.DIODE(clknet_5_10_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_77_i_clk_A (.DIODE(clknet_5_10_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_76_i_clk_A (.DIODE(clknet_5_10_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_75_i_clk_A (.DIODE(clknet_5_10_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_74_i_clk_A (.DIODE(clknet_5_10_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_73_i_clk_A (.DIODE(clknet_5_10_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_72_i_clk_A (.DIODE(clknet_5_10_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_85_i_clk_A (.DIODE(clknet_5_11_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_84_i_clk_A (.DIODE(clknet_5_11_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_83_i_clk_A (.DIODE(clknet_5_11_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_82_i_clk_A (.DIODE(clknet_5_11_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_81_i_clk_A (.DIODE(clknet_5_11_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_80_i_clk_A (.DIODE(clknet_5_11_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_79_i_clk_A (.DIODE(clknet_5_11_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_71_i_clk_A (.DIODE(clknet_5_11_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_70_i_clk_A (.DIODE(clknet_5_11_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_105_i_clk_A (.DIODE(clknet_5_12_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_104_i_clk_A (.DIODE(clknet_5_12_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_i_clk_A (.DIODE(clknet_5_12_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_i_clk_A (.DIODE(clknet_5_12_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_i_clk_A (.DIODE(clknet_5_12_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_i_clk_A (.DIODE(clknet_5_12_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_i_clk_A (.DIODE(clknet_5_12_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_i_clk_A (.DIODE(clknet_5_12_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_i_clk_A (.DIODE(clknet_5_12_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_112_i_clk_A (.DIODE(clknet_5_13_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_111_i_clk_A (.DIODE(clknet_5_13_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_110_i_clk_A (.DIODE(clknet_5_13_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_109_i_clk_A (.DIODE(clknet_5_13_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_108_i_clk_A (.DIODE(clknet_5_13_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_107_i_clk_A (.DIODE(clknet_5_13_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_106_i_clk_A (.DIODE(clknet_5_13_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_i_clk_A (.DIODE(clknet_5_13_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_i_clk_A (.DIODE(clknet_5_13_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_103_i_clk_A (.DIODE(clknet_5_14_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_102_i_clk_A (.DIODE(clknet_5_14_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_101_i_clk_A (.DIODE(clknet_5_14_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_92_i_clk_A (.DIODE(clknet_5_14_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_91_i_clk_A (.DIODE(clknet_5_14_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_90_i_clk_A (.DIODE(clknet_5_14_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_89_i_clk_A (.DIODE(clknet_5_14_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_88_i_clk_A (.DIODE(clknet_5_14_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_87_i_clk_A (.DIODE(clknet_5_14_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_86_i_clk_A (.DIODE(clknet_5_14_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_100_i_clk_A (.DIODE(clknet_5_15_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_99_i_clk_A (.DIODE(clknet_5_15_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_98_i_clk_A (.DIODE(clknet_5_15_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_97_i_clk_A (.DIODE(clknet_5_15_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_96_i_clk_A (.DIODE(clknet_5_15_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_95_i_clk_A (.DIODE(clknet_5_15_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_94_i_clk_A (.DIODE(clknet_5_15_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_93_i_clk_A (.DIODE(clknet_5_15_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_241_i_clk_A (.DIODE(clknet_5_16_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_240_i_clk_A (.DIODE(clknet_5_16_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_239_i_clk_A (.DIODE(clknet_5_16_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_238_i_clk_A (.DIODE(clknet_5_16_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_237_i_clk_A (.DIODE(clknet_5_16_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_236_i_clk_A (.DIODE(clknet_5_16_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_235_i_clk_A (.DIODE(clknet_5_16_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_234_i_clk_A (.DIODE(clknet_5_16_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_242_i_clk_A (.DIODE(clknet_5_17_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_233_i_clk_A (.DIODE(clknet_5_17_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_232_i_clk_A (.DIODE(clknet_5_17_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_231_i_clk_A (.DIODE(clknet_5_17_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_230_i_clk_A (.DIODE(clknet_5_17_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_229_i_clk_A (.DIODE(clknet_5_17_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_228_i_clk_A (.DIODE(clknet_5_17_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_227_i_clk_A (.DIODE(clknet_5_17_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_251_i_clk_A (.DIODE(clknet_5_18_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_250_i_clk_A (.DIODE(clknet_5_18_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_249_i_clk_A (.DIODE(clknet_5_18_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_248_i_clk_A (.DIODE(clknet_5_18_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_247_i_clk_A (.DIODE(clknet_5_18_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_246_i_clk_A (.DIODE(clknet_5_18_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_182_i_clk_A (.DIODE(clknet_5_18_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_181_i_clk_A (.DIODE(clknet_5_18_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_245_i_clk_A (.DIODE(clknet_5_19_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_244_i_clk_A (.DIODE(clknet_5_19_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_243_i_clk_A (.DIODE(clknet_5_19_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_189_i_clk_A (.DIODE(clknet_5_19_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_188_i_clk_A (.DIODE(clknet_5_19_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_187_i_clk_A (.DIODE(clknet_5_19_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_186_i_clk_A (.DIODE(clknet_5_19_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_185_i_clk_A (.DIODE(clknet_5_19_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_184_i_clk_A (.DIODE(clknet_5_19_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_183_i_clk_A (.DIODE(clknet_5_19_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_226_i_clk_A (.DIODE(clknet_5_20_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_225_i_clk_A (.DIODE(clknet_5_20_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_224_i_clk_A (.DIODE(clknet_5_20_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_223_i_clk_A (.DIODE(clknet_5_20_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_222_i_clk_A (.DIODE(clknet_5_20_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_221_i_clk_A (.DIODE(clknet_5_20_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_210_i_clk_A (.DIODE(clknet_5_20_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_209_i_clk_A (.DIODE(clknet_5_20_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_220_i_clk_A (.DIODE(clknet_5_21_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_219_i_clk_A (.DIODE(clknet_5_21_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_218_i_clk_A (.DIODE(clknet_5_21_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_217_i_clk_A (.DIODE(clknet_5_21_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_216_i_clk_A (.DIODE(clknet_5_21_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_215_i_clk_A (.DIODE(clknet_5_21_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_214_i_clk_A (.DIODE(clknet_5_21_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_213_i_clk_A (.DIODE(clknet_5_21_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_212_i_clk_A (.DIODE(clknet_5_21_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_211_i_clk_A (.DIODE(clknet_5_21_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_208_i_clk_A (.DIODE(clknet_5_22_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_207_i_clk_A (.DIODE(clknet_5_22_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_196_i_clk_A (.DIODE(clknet_5_22_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_195_i_clk_A (.DIODE(clknet_5_22_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_194_i_clk_A (.DIODE(clknet_5_22_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_193_i_clk_A (.DIODE(clknet_5_22_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_192_i_clk_A (.DIODE(clknet_5_22_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_191_i_clk_A (.DIODE(clknet_5_22_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_190_i_clk_A (.DIODE(clknet_5_22_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_206_i_clk_A (.DIODE(clknet_5_23_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_205_i_clk_A (.DIODE(clknet_5_23_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_204_i_clk_A (.DIODE(clknet_5_23_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_203_i_clk_A (.DIODE(clknet_5_23_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_202_i_clk_A (.DIODE(clknet_5_23_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_201_i_clk_A (.DIODE(clknet_5_23_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_200_i_clk_A (.DIODE(clknet_5_23_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_199_i_clk_A (.DIODE(clknet_5_23_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_198_i_clk_A (.DIODE(clknet_5_23_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_197_i_clk_A (.DIODE(clknet_5_23_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_180_i_clk_A (.DIODE(clknet_5_24_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_179_i_clk_A (.DIODE(clknet_5_24_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_118_i_clk_A (.DIODE(clknet_5_24_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_117_i_clk_A (.DIODE(clknet_5_24_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_116_i_clk_A (.DIODE(clknet_5_24_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_115_i_clk_A (.DIODE(clknet_5_24_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_114_i_clk_A (.DIODE(clknet_5_24_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_113_i_clk_A (.DIODE(clknet_5_24_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_178_i_clk_A (.DIODE(clknet_5_25_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_177_i_clk_A (.DIODE(clknet_5_25_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_176_i_clk_A (.DIODE(clknet_5_25_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_175_i_clk_A (.DIODE(clknet_5_25_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_174_i_clk_A (.DIODE(clknet_5_25_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_173_i_clk_A (.DIODE(clknet_5_25_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_120_i_clk_A (.DIODE(clknet_5_25_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_119_i_clk_A (.DIODE(clknet_5_25_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_132_i_clk_A (.DIODE(clknet_5_26_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_131_i_clk_A (.DIODE(clknet_5_26_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_130_i_clk_A (.DIODE(clknet_5_26_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_129_i_clk_A (.DIODE(clknet_5_26_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_128_i_clk_A (.DIODE(clknet_5_26_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_127_i_clk_A (.DIODE(clknet_5_26_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_126_i_clk_A (.DIODE(clknet_5_26_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_125_i_clk_A (.DIODE(clknet_5_26_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_124_i_clk_A (.DIODE(clknet_5_26_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_139_i_clk_A (.DIODE(clknet_5_27_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_138_i_clk_A (.DIODE(clknet_5_27_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_137_i_clk_A (.DIODE(clknet_5_27_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_136_i_clk_A (.DIODE(clknet_5_27_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_135_i_clk_A (.DIODE(clknet_5_27_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_134_i_clk_A (.DIODE(clknet_5_27_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_133_i_clk_A (.DIODE(clknet_5_27_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_123_i_clk_A (.DIODE(clknet_5_27_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_122_i_clk_A (.DIODE(clknet_5_27_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_121_i_clk_A (.DIODE(clknet_5_27_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_172_i_clk_A (.DIODE(clknet_5_28_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_171_i_clk_A (.DIODE(clknet_5_28_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_170_i_clk_A (.DIODE(clknet_5_28_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_169_i_clk_A (.DIODE(clknet_5_28_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_168_i_clk_A (.DIODE(clknet_5_28_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_159_i_clk_A (.DIODE(clknet_5_28_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_158_i_clk_A (.DIODE(clknet_5_28_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_167_i_clk_A (.DIODE(clknet_5_29_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_166_i_clk_A (.DIODE(clknet_5_29_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_165_i_clk_A (.DIODE(clknet_5_29_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_164_i_clk_A (.DIODE(clknet_5_29_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_163_i_clk_A (.DIODE(clknet_5_29_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_162_i_clk_A (.DIODE(clknet_5_29_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_161_i_clk_A (.DIODE(clknet_5_29_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_160_i_clk_A (.DIODE(clknet_5_29_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_157_i_clk_A (.DIODE(clknet_5_30_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_156_i_clk_A (.DIODE(clknet_5_30_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_146_i_clk_A (.DIODE(clknet_5_30_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_145_i_clk_A (.DIODE(clknet_5_30_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_144_i_clk_A (.DIODE(clknet_5_30_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_143_i_clk_A (.DIODE(clknet_5_30_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_142_i_clk_A (.DIODE(clknet_5_30_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_141_i_clk_A (.DIODE(clknet_5_30_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_140_i_clk_A (.DIODE(clknet_5_30_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_155_i_clk_A (.DIODE(clknet_5_31_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_154_i_clk_A (.DIODE(clknet_5_31_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_153_i_clk_A (.DIODE(clknet_5_31_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_152_i_clk_A (.DIODE(clknet_5_31_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_151_i_clk_A (.DIODE(clknet_5_31_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_150_i_clk_A (.DIODE(clknet_5_31_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_149_i_clk_A (.DIODE(clknet_5_31_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_148_i_clk_A (.DIODE(clknet_5_31_0_i_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_147_i_clk_A (.DIODE(clknet_5_31_0_i_clk));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_770 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1016 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_868 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_396 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1105 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1106 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1140 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1019 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_750 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_988 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1129 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_779 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_980 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1141 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_946 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1124 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_760 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_227 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1014 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_690 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1111 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_1164 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1008 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1123 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_820 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_959 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_994 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_570 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_802 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_308 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_756 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_863 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1059 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1116 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_236 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1099 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1124 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_910 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1136 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1155 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_396 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1000 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1094 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_1098 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1134 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1136 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1082 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1002 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1059 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1106 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1058 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_346 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_999 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1108 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_521 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_859 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1084 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1091 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_899 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_968 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_529 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_935 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1150 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1156 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1061 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1067 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1134 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_240 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_990 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1152 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_950 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1139 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_226 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_900 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_264 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_1142 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1162 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_951 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1025 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1042 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1083 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1104 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1117 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_270 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1030 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1083 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1151 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_336 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1054 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_339 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_938 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1112 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1124 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_822 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_871 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_986 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1042 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_850 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_891 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1120 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_974 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1106 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_745 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1016 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1124 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_927 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_1036 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_1130 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_799 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_788 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1019 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1115 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1088 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_955 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1115 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1040 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_1107 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1111 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1117 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1025 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_326 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_850 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1159 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1163 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_810 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_913 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1022 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_888 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1078 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1082 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1112 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_833 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_967 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_984 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_619 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_790 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_954 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1056 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1072 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_323 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_870 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1001 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1126 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_115 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_451 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1130 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1025 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_861 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_30 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1114 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_1142 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1012 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_574 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1050 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1073 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1108 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1053 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_366 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1141 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1162 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_632 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1012 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1056 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1073 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_123 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_804 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1162 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_103 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_282 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_840 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_956 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_703 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_709 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_704 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_914 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_939 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_1138 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_746 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1002 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_1141 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_463 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1069 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_864 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_945 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_994 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1102 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1108 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1059 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1071 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1166 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1140 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1144 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_392 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_24 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_28 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_700 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_803 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1052 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1102 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1142 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1018 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1048 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_10 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_200 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_858 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1035 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1104 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1143 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1166 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_456 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1124 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1130 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_142 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1002 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1087 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1125 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1111 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_28 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_88 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_861 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1104 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1157 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1053 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1111 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1154 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1141 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_26 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1012 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1026 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_584 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_802 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1079 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1103 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1041 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_1144 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1167 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_821 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_970 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1028 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1040 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_103 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_672 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_679 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_955 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1013 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1113 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1092 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_960 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1011 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_12 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_146 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1041 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_12 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_990 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1088 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1123 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1166 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_298 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_827 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1011 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1122 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_129 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_984 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1136 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1148 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1010 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1113 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1052 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1083 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1141 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_778 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1006 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1074 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1111 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1131 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_511 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1050 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1081 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1148 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_570 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_843 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1141 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_1165 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_998 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1088 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1094 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1114 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_22 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_252 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_497 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1079 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1098 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1120 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_758 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_951 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_975 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1020 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_914 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_958 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1018 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_918 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_983 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1024 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_680 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_904 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_995 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1132 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1159 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_103 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_598 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_918 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_924 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1095 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1167 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1138 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_143 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_863 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1041 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1060 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1082 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1118 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1126 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1136 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_189 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_578 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_636 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_799 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_820 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1028 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1128 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1140 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_952 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_956 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1128 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_79 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_303 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_950 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_982 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_995 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1083 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1118 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1137 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_497 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_687 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1010 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1022 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1088 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_969 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1018 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1024 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1087 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1016 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1035 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1097 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1129 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1133 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_259 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_409 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_412 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_653 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_860 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_877 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_940 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1076 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1134 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1147 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1151 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1155 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_864 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1001 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1111 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1126 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_311 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_329 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_772 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_863 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1004 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1078 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1144 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_532 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1036 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1046 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1076 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1137 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_1154 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_270 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_398 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1001 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1050 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1079 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1147 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_104 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1042 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1107 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1147 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1164 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_998 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1046 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1111 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1143 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_88 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_700 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1040 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1145 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_451 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1090 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_131 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_367 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_662 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_901 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_984 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1026 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1030 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1051 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1095 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_1107 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1115 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1139 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_106 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_883 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_987 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1127 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_134 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_370 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_928 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_995 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1075 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1135 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1142 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1162 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_115 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_752 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1060 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1066 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1115 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1137 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1153 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1165 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1088 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1095 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1139 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1151 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_508 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_892 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1022 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1051 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1064 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1072 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1114 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1121 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_817 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1096 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1142 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_226 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_817 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_908 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_955 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_961 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1055 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1114 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1120 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1126 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1130 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_368 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_872 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1026 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_1135 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1149 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_133 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_896 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1088 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1136 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_814 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_861 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_942 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1075 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1109 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1118 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1141 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_453 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1024 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1123 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_11 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_84 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1043 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1054 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_824 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_852 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_954 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1048 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1056 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1068 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1129 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_973 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1053 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1090 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1094 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1100 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1133 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_394 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_774 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_847 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_898 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1006 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1012 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1054 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_892 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1038 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1156 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_180 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_297 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_775 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_858 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_200 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_873 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_971 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_984 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1139 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1143 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_964 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1098 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1104 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1110 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1118 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_31 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_879 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1032 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_1145 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_1165 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1047 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1062 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1082 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1138 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1166 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1027 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1054 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1061 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1079 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_1117 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1139 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1150 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1166 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_11 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_790 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_943 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_964 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1001 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1078 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1118 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1124 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1140 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_590 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_718 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1062 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1135 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_523 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_680 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_733 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_800 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1128 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1154 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_470 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_886 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_964 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1028 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1045 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1051 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1082 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1167 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_923 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1052 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1097 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1100 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1106 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1110 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1116 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_587 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_702 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_992 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1044 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1086 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1092 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1096 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1105 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1111 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_1117 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1129 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1142 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_1158 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_20 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_544 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_851 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_945 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_958 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1103 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1107 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1147 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_582 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1119 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_211 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_948 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1047 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1063 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1088 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_87 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_928 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1051 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1069 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1096 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1121 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1125 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_116 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_134 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_619 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_728 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_899 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_912 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_954 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_966 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_978 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1000 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1008 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1034 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1084 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_49 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_591 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_816 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_872 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_967 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_994 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1041 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1108 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1112 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1116 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1125 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1131 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1137 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_886 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1104 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1110 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1162 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_816 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_986 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1055 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1061 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1100 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1132 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_905 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_954 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1051 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1080 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1088 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1121 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_692 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_907 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1044 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1099 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_1106 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1114 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1132 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1144 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_351 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_793 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_956 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_970 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1031 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1109 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1123 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1132 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_248 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_299 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_762 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_949 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_982 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1086 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_1092 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1127 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1138 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_284 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_676 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_728 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_821 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_965 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1003 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1027 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1067 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1133 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1137 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1155 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_805 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1030 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1063 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1082 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_1088 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1096 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1119 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1127 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1131 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1153 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_605 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1004 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1023 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1055 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1064 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1070 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1076 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1080 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1086 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1099 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1109 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1142 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_1165 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_480 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_604 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_970 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1007 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1069 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1112 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1132 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1138 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1146 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_550 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_575 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_780 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_844 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_964 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1011 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1032 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1115 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1135 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1160 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_186 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_311 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_756 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_908 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_982 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1027 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1047 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1116 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1143 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1149 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1157 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_271 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_948 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_960 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1007 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1013 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1054 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1060 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1104 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1116 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1122 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1135 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1147 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1153 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1161 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1166 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_862 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1028 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1037 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1069 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1081 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1097 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1103 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1109 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1115 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1119 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1121 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1127 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1131 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1145 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1153 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1159 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1165 ();
endmodule

