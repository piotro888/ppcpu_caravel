magic
tech sky130B
magscale 1 2
timestamp 1663051562
<< viali >>
rect 4629 47209 4663 47243
rect 9873 47209 9907 47243
rect 10977 47209 11011 47243
rect 13461 47209 13495 47243
rect 15945 47209 15979 47243
rect 18153 47209 18187 47243
rect 20085 47209 20119 47243
rect 20913 47209 20947 47243
rect 22477 47209 22511 47243
rect 27169 47209 27203 47243
rect 27905 47209 27939 47243
rect 30573 47209 30607 47243
rect 31309 47209 31343 47243
rect 32321 47209 32355 47243
rect 36645 47209 36679 47243
rect 2973 47141 3007 47175
rect 6745 47141 6779 47175
rect 19441 47141 19475 47175
rect 28641 47141 28675 47175
rect 1501 47073 1535 47107
rect 7205 47073 7239 47107
rect 14289 47073 14323 47107
rect 23029 47073 23063 47107
rect 24409 47073 24443 47107
rect 32965 47073 32999 47107
rect 34897 47073 34931 47107
rect 37565 47073 37599 47107
rect 2053 47005 2087 47039
rect 3893 47005 3927 47039
rect 4813 47005 4847 47039
rect 5365 47005 5399 47039
rect 6561 47005 6595 47039
rect 7481 47005 7515 47039
rect 9137 47005 9171 47039
rect 10057 47005 10091 47039
rect 10793 47005 10827 47039
rect 11989 47005 12023 47039
rect 12633 47005 12667 47039
rect 13277 47005 13311 47039
rect 14565 47005 14599 47039
rect 16129 47005 16163 47039
rect 16681 47005 16715 47039
rect 16957 47005 16991 47039
rect 17969 47005 18003 47039
rect 19625 47005 19659 47039
rect 20269 47005 20303 47039
rect 20729 47005 20763 47039
rect 22293 47005 22327 47039
rect 23305 47005 23339 47039
rect 24685 47005 24719 47039
rect 26065 47005 26099 47039
rect 26985 47005 27019 47039
rect 27721 47005 27755 47039
rect 28457 47005 28491 47039
rect 29745 47005 29779 47039
rect 30389 47005 30423 47039
rect 31125 47005 31159 47039
rect 32137 47005 32171 47039
rect 33241 47005 33275 47039
rect 35173 47005 35207 47039
rect 36461 47005 36495 47039
rect 37289 47005 37323 47039
rect 2237 46937 2271 46971
rect 2789 46937 2823 46971
rect 4077 46937 4111 46971
rect 5549 46937 5583 46971
rect 9321 46937 9355 46971
rect 25881 46937 25915 46971
rect 12173 46869 12207 46903
rect 12817 46869 12851 46903
rect 29561 46869 29595 46903
rect 3709 46665 3743 46699
rect 5181 46665 5215 46699
rect 5825 46665 5859 46699
rect 7113 46665 7147 46699
rect 7941 46665 7975 46699
rect 10885 46665 10919 46699
rect 13829 46665 13863 46699
rect 15853 46665 15887 46699
rect 17417 46665 17451 46699
rect 19993 46665 20027 46699
rect 21281 46665 21315 46699
rect 23949 46665 23983 46699
rect 25881 46665 25915 46699
rect 35173 46665 35207 46699
rect 36645 46665 36679 46699
rect 2973 46597 3007 46631
rect 15025 46597 15059 46631
rect 32689 46597 32723 46631
rect 2237 46529 2271 46563
rect 3893 46529 3927 46563
rect 4353 46529 4387 46563
rect 6377 46529 6411 46563
rect 8125 46529 8159 46563
rect 8677 46529 8711 46563
rect 9137 46529 9171 46563
rect 11713 46529 11747 46563
rect 13737 46529 13771 46563
rect 14933 46529 14967 46563
rect 16037 46529 16071 46563
rect 17509 46529 17543 46563
rect 18797 46529 18831 46563
rect 21833 46529 21867 46563
rect 22661 46529 22695 46563
rect 23121 46529 23155 46563
rect 24777 46529 24811 46563
rect 25237 46529 25271 46563
rect 28641 46529 28675 46563
rect 29101 46529 29135 46563
rect 29929 46529 29963 46563
rect 30389 46529 30423 46563
rect 33793 46529 33827 46563
rect 34437 46529 34471 46563
rect 34989 46529 35023 46563
rect 35909 46529 35943 46563
rect 36461 46529 36495 46563
rect 37289 46529 37323 46563
rect 12909 46461 12943 46495
rect 14013 46461 14047 46495
rect 15209 46461 15243 46495
rect 17233 46461 17267 46495
rect 37565 46461 37599 46495
rect 2421 46393 2455 46427
rect 9321 46393 9355 46427
rect 24593 46393 24627 46427
rect 29745 46393 29779 46427
rect 34253 46393 34287 46427
rect 35725 46393 35759 46427
rect 1685 46325 1719 46359
rect 3065 46325 3099 46359
rect 4537 46325 4571 46359
rect 6561 46325 6595 46359
rect 10241 46325 10275 46359
rect 11897 46325 11931 46359
rect 13369 46325 13403 46359
rect 14565 46325 14599 46359
rect 17877 46325 17911 46359
rect 18981 46325 19015 46359
rect 22017 46325 22051 46359
rect 22477 46325 22511 46359
rect 27905 46325 27939 46359
rect 28457 46325 28491 46359
rect 30941 46325 30975 46359
rect 31493 46325 31527 46359
rect 32597 46325 32631 46359
rect 33609 46325 33643 46359
rect 2237 46121 2271 46155
rect 2973 46121 3007 46155
rect 4169 46121 4203 46155
rect 4905 46121 4939 46155
rect 6469 46121 6503 46155
rect 8953 46121 8987 46155
rect 11621 46121 11655 46155
rect 12173 46121 12207 46155
rect 15117 46121 15151 46155
rect 19349 46121 19383 46155
rect 24409 46121 24443 46155
rect 29653 46121 29687 46155
rect 32321 46121 32355 46155
rect 32965 46121 32999 46155
rect 33517 46121 33551 46155
rect 34161 46121 34195 46155
rect 36737 46121 36771 46155
rect 5549 46053 5583 46087
rect 13277 46053 13311 46087
rect 14473 46053 14507 46087
rect 36001 46053 36035 46087
rect 16681 45985 16715 46019
rect 16865 45985 16899 46019
rect 37289 45985 37323 46019
rect 1685 45917 1719 45951
rect 2421 45917 2455 45951
rect 3157 45917 3191 45951
rect 12817 45917 12851 45951
rect 13461 45917 13495 45951
rect 14289 45917 14323 45951
rect 14933 45917 14967 45951
rect 16957 45917 16991 45951
rect 18337 45917 18371 45951
rect 35357 45917 35391 45951
rect 35817 45917 35851 45951
rect 36553 45917 36587 45951
rect 37565 45917 37599 45951
rect 8309 45849 8343 45883
rect 1501 45781 1535 45815
rect 16037 45781 16071 45815
rect 17325 45781 17359 45815
rect 18153 45781 18187 45815
rect 35173 45781 35207 45815
rect 18705 45577 18739 45611
rect 35449 45577 35483 45611
rect 4353 45509 4387 45543
rect 12909 45509 12943 45543
rect 13921 45509 13955 45543
rect 17141 45509 17175 45543
rect 34345 45509 34379 45543
rect 37381 45509 37415 45543
rect 1869 45441 1903 45475
rect 2513 45441 2547 45475
rect 4905 45441 4939 45475
rect 17785 45441 17819 45475
rect 33793 45441 33827 45475
rect 36737 45441 36771 45475
rect 37841 45441 37875 45475
rect 3801 45373 3835 45407
rect 2053 45305 2087 45339
rect 2697 45305 2731 45339
rect 17325 45305 17359 45339
rect 17969 45305 18003 45339
rect 36001 45305 36035 45339
rect 3249 45237 3283 45271
rect 14381 45237 14415 45271
rect 15393 45237 15427 45271
rect 16037 45237 16071 45271
rect 34805 45237 34839 45271
rect 36553 45237 36587 45271
rect 38025 45237 38059 45271
rect 3801 45033 3835 45067
rect 16681 45033 16715 45067
rect 18061 45033 18095 45067
rect 36093 45033 36127 45067
rect 37197 44965 37231 44999
rect 33609 44897 33643 44931
rect 35633 44897 35667 44931
rect 2513 44829 2547 44863
rect 3157 44829 3191 44863
rect 33793 44829 33827 44863
rect 36737 44829 36771 44863
rect 37381 44829 37415 44863
rect 38025 44829 38059 44863
rect 1869 44761 1903 44795
rect 32873 44761 32907 44795
rect 33701 44761 33735 44795
rect 35081 44761 35115 44795
rect 1961 44693 1995 44727
rect 2697 44693 2731 44727
rect 16221 44693 16255 44727
rect 34161 44693 34195 44727
rect 37933 44693 37967 44727
rect 2697 44489 2731 44523
rect 3157 44421 3191 44455
rect 1409 44353 1443 44387
rect 2053 44353 2087 44387
rect 22937 44353 22971 44387
rect 37841 44353 37875 44387
rect 21833 44285 21867 44319
rect 22293 44285 22327 44319
rect 22109 44217 22143 44251
rect 23121 44217 23155 44251
rect 38025 44217 38059 44251
rect 1593 44149 1627 44183
rect 33333 44149 33367 44183
rect 35725 44149 35759 44183
rect 36277 44149 36311 44183
rect 37289 44149 37323 44183
rect 22477 43945 22511 43979
rect 36277 43945 36311 43979
rect 1409 43741 1443 43775
rect 2053 43741 2087 43775
rect 34713 43741 34747 43775
rect 37289 43741 37323 43775
rect 37565 43741 37599 43775
rect 1593 43605 1627 43639
rect 26985 43605 27019 43639
rect 34897 43605 34931 43639
rect 36737 43605 36771 43639
rect 26249 43401 26283 43435
rect 27537 43401 27571 43435
rect 1409 43265 1443 43299
rect 2053 43265 2087 43299
rect 5181 43265 5215 43299
rect 26433 43265 26467 43299
rect 27445 43265 27479 43299
rect 37381 43265 37415 43299
rect 38025 43265 38059 43299
rect 4905 43197 4939 43231
rect 27721 43197 27755 43231
rect 1593 43129 1627 43163
rect 37841 43129 37875 43163
rect 27077 43061 27111 43095
rect 4721 42857 4755 42891
rect 27445 42857 27479 42891
rect 4169 42721 4203 42755
rect 4261 42721 4295 42755
rect 27997 42721 28031 42755
rect 1409 42653 1443 42687
rect 2053 42653 2087 42687
rect 26433 42653 26467 42687
rect 27905 42653 27939 42687
rect 37473 42653 37507 42687
rect 38117 42653 38151 42687
rect 4353 42585 4387 42619
rect 27813 42585 27847 42619
rect 1593 42517 1627 42551
rect 5181 42517 5215 42551
rect 26341 42517 26375 42551
rect 37933 42517 37967 42551
rect 20729 42313 20763 42347
rect 27353 42313 27387 42347
rect 27169 42177 27203 42211
rect 1685 41973 1719 42007
rect 3801 41973 3835 42007
rect 27813 41973 27847 42007
rect 22569 41769 22603 41803
rect 37933 41769 37967 41803
rect 20729 41633 20763 41667
rect 21373 41633 21407 41667
rect 1869 41565 1903 41599
rect 21465 41565 21499 41599
rect 22385 41565 22419 41599
rect 37473 41565 37507 41599
rect 38117 41565 38151 41599
rect 2053 41497 2087 41531
rect 21557 41429 21591 41463
rect 21925 41429 21959 41463
rect 27537 41225 27571 41259
rect 28733 41225 28767 41259
rect 27997 41157 28031 41191
rect 27905 41089 27939 41123
rect 37473 41089 37507 41123
rect 38117 41089 38151 41123
rect 1961 41021 1995 41055
rect 2237 41021 2271 41055
rect 2697 41021 2731 41055
rect 26985 41021 27019 41055
rect 28089 41021 28123 41055
rect 37933 40953 37967 40987
rect 20913 40885 20947 40919
rect 37473 40477 37507 40511
rect 38117 40477 38151 40511
rect 1869 40409 1903 40443
rect 2053 40409 2087 40443
rect 2513 40341 2547 40375
rect 37933 40341 37967 40375
rect 37381 40001 37415 40035
rect 37841 40001 37875 40035
rect 1409 39933 1443 39967
rect 1685 39933 1719 39967
rect 38025 39797 38059 39831
rect 22661 39593 22695 39627
rect 1409 39525 1443 39559
rect 20269 39457 20303 39491
rect 19625 39389 19659 39423
rect 20637 39389 20671 39423
rect 22063 39389 22097 39423
rect 21143 39049 21177 39083
rect 21925 38981 21959 39015
rect 1685 38913 1719 38947
rect 2237 38913 2271 38947
rect 19717 38913 19751 38947
rect 22017 38913 22051 38947
rect 22477 38913 22511 38947
rect 37841 38913 37875 38947
rect 19349 38845 19383 38879
rect 1501 38777 1535 38811
rect 38025 38777 38059 38811
rect 37289 38709 37323 38743
rect 20729 38505 20763 38539
rect 21925 38505 21959 38539
rect 1961 38301 1995 38335
rect 2237 38301 2271 38335
rect 2697 38301 2731 38335
rect 20637 38301 20671 38335
rect 21281 38301 21315 38335
rect 37473 38301 37507 38335
rect 38117 38301 38151 38335
rect 37933 38165 37967 38199
rect 8401 37961 8435 37995
rect 8585 37825 8619 37859
rect 37841 37825 37875 37859
rect 1961 37757 1995 37791
rect 2237 37757 2271 37791
rect 2697 37757 2731 37791
rect 38025 37621 38059 37655
rect 9045 37417 9079 37451
rect 22753 37417 22787 37451
rect 9597 37281 9631 37315
rect 1685 37213 1719 37247
rect 9505 37213 9539 37247
rect 22017 37213 22051 37247
rect 37841 37213 37875 37247
rect 38117 37213 38151 37247
rect 9413 37145 9447 37179
rect 10333 37145 10367 37179
rect 1501 37077 1535 37111
rect 2145 37077 2179 37111
rect 22201 37077 22235 37111
rect 22201 36873 22235 36907
rect 22293 36873 22327 36907
rect 23489 36873 23523 36907
rect 38117 36805 38151 36839
rect 22385 36669 22419 36703
rect 9965 36533 9999 36567
rect 21189 36533 21223 36567
rect 21833 36533 21867 36567
rect 22109 36329 22143 36363
rect 23765 36329 23799 36363
rect 24409 36329 24443 36363
rect 23121 36261 23155 36295
rect 21557 36193 21591 36227
rect 1685 36125 1719 36159
rect 21649 36125 21683 36159
rect 37841 36125 37875 36159
rect 1501 35989 1535 36023
rect 20821 35989 20855 36023
rect 21741 35989 21775 36023
rect 22661 35989 22695 36023
rect 38025 35989 38059 36023
rect 6929 35785 6963 35819
rect 7573 35785 7607 35819
rect 22937 35785 22971 35819
rect 24409 35785 24443 35819
rect 24501 35785 24535 35819
rect 22845 35717 22879 35751
rect 1685 35649 1719 35683
rect 7113 35649 7147 35683
rect 7941 35649 7975 35683
rect 37473 35649 37507 35683
rect 38117 35649 38151 35683
rect 8033 35581 8067 35615
rect 8217 35581 8251 35615
rect 21925 35581 21959 35615
rect 23029 35581 23063 35615
rect 24225 35581 24259 35615
rect 25329 35581 25363 35615
rect 1501 35445 1535 35479
rect 2237 35445 2271 35479
rect 8769 35445 8803 35479
rect 9413 35445 9447 35479
rect 22477 35445 22511 35479
rect 24869 35445 24903 35479
rect 37933 35445 37967 35479
rect 2145 35241 2179 35275
rect 22661 35241 22695 35275
rect 23305 35241 23339 35275
rect 22569 35105 22603 35139
rect 1685 35037 1719 35071
rect 2329 35037 2363 35071
rect 21925 35037 21959 35071
rect 22385 35037 22419 35071
rect 22661 35037 22695 35071
rect 24869 35037 24903 35071
rect 21373 34969 21407 35003
rect 25053 34969 25087 35003
rect 1501 34901 1535 34935
rect 22845 34901 22879 34935
rect 23213 34697 23247 34731
rect 27537 34697 27571 34731
rect 37933 34697 37967 34731
rect 22385 34629 22419 34663
rect 1961 34561 1995 34595
rect 22201 34561 22235 34595
rect 27353 34561 27387 34595
rect 37473 34561 37507 34595
rect 38117 34561 38151 34595
rect 2237 34493 2271 34527
rect 2697 34493 2731 34527
rect 2329 34153 2363 34187
rect 22385 34153 22419 34187
rect 27353 34153 27387 34187
rect 23213 34085 23247 34119
rect 1685 34017 1719 34051
rect 21833 34017 21867 34051
rect 26709 34017 26743 34051
rect 1961 33949 1995 33983
rect 21557 33949 21591 33983
rect 22569 33949 22603 33983
rect 26893 33881 26927 33915
rect 1869 33813 1903 33847
rect 2881 33813 2915 33847
rect 25513 33813 25547 33847
rect 26157 33813 26191 33847
rect 26985 33813 27019 33847
rect 1593 33609 1627 33643
rect 5457 33609 5491 33643
rect 17877 33609 17911 33643
rect 22293 33609 22327 33643
rect 22753 33609 22787 33643
rect 1409 33473 1443 33507
rect 2053 33473 2087 33507
rect 5549 33473 5583 33507
rect 6377 33473 6411 33507
rect 17785 33473 17819 33507
rect 22661 33473 22695 33507
rect 37473 33473 37507 33507
rect 38117 33473 38151 33507
rect 5641 33405 5675 33439
rect 17049 33405 17083 33439
rect 17693 33405 17727 33439
rect 22937 33405 22971 33439
rect 23489 33405 23523 33439
rect 21189 33337 21223 33371
rect 37933 33337 37967 33371
rect 5089 33269 5123 33303
rect 18245 33269 18279 33303
rect 5917 33065 5951 33099
rect 17141 33065 17175 33099
rect 22201 33065 22235 33099
rect 29745 33065 29779 33099
rect 23029 32997 23063 33031
rect 22661 32929 22695 32963
rect 1409 32861 1443 32895
rect 2053 32861 2087 32895
rect 22017 32861 22051 32895
rect 29561 32861 29595 32895
rect 37473 32861 37507 32895
rect 38117 32861 38151 32895
rect 23581 32793 23615 32827
rect 1593 32725 1627 32759
rect 21281 32725 21315 32759
rect 23121 32725 23155 32759
rect 37933 32725 37967 32759
rect 20085 32521 20119 32555
rect 22201 32521 22235 32555
rect 22569 32521 22603 32555
rect 23673 32521 23707 32555
rect 24501 32521 24535 32555
rect 29377 32521 29411 32555
rect 37933 32521 37967 32555
rect 22109 32453 22143 32487
rect 23581 32453 23615 32487
rect 1685 32385 1719 32419
rect 21097 32385 21131 32419
rect 29009 32385 29043 32419
rect 37473 32385 37507 32419
rect 38117 32385 38151 32419
rect 21925 32317 21959 32351
rect 23765 32317 23799 32351
rect 28733 32317 28767 32351
rect 28917 32317 28951 32351
rect 29837 32317 29871 32351
rect 21281 32249 21315 32283
rect 28089 32249 28123 32283
rect 1501 32181 1535 32215
rect 23213 32181 23247 32215
rect 2697 31977 2731 32011
rect 21373 31977 21407 32011
rect 21925 31977 21959 32011
rect 23397 31977 23431 32011
rect 15669 31909 15703 31943
rect 17325 31909 17359 31943
rect 1685 31841 1719 31875
rect 17877 31841 17911 31875
rect 20177 31841 20211 31875
rect 20729 31841 20763 31875
rect 20913 31841 20947 31875
rect 23121 31841 23155 31875
rect 23238 31841 23272 31875
rect 37841 31841 37875 31875
rect 1409 31773 1443 31807
rect 2881 31773 2915 31807
rect 15025 31773 15059 31807
rect 15117 31773 15151 31807
rect 16865 31773 16899 31807
rect 18153 31773 18187 31807
rect 22753 31773 22787 31807
rect 28457 31773 28491 31807
rect 37381 31773 37415 31807
rect 38025 31773 38059 31807
rect 23029 31705 23063 31739
rect 16773 31637 16807 31671
rect 21005 31637 21039 31671
rect 24409 31637 24443 31671
rect 2329 31433 2363 31467
rect 20269 31433 20303 31467
rect 21833 31433 21867 31467
rect 23305 31433 23339 31467
rect 23857 31433 23891 31467
rect 1961 31365 1995 31399
rect 2789 31365 2823 31399
rect 22753 31365 22787 31399
rect 5181 31297 5215 31331
rect 14197 31297 14231 31331
rect 1685 31229 1719 31263
rect 1869 31229 1903 31263
rect 14565 31229 14599 31263
rect 15991 31229 16025 31263
rect 17233 31229 17267 31263
rect 22569 31229 22603 31263
rect 4997 31093 5031 31127
rect 16681 31093 16715 31127
rect 24501 31093 24535 31127
rect 1409 30889 1443 30923
rect 14565 30889 14599 30923
rect 17187 30821 17221 30855
rect 15393 30753 15427 30787
rect 15761 30753 15795 30787
rect 23489 30753 23523 30787
rect 23581 30753 23615 30787
rect 22477 30549 22511 30583
rect 23029 30549 23063 30583
rect 23397 30549 23431 30583
rect 24409 30549 24443 30583
rect 22569 30277 22603 30311
rect 24317 30277 24351 30311
rect 1685 30209 1719 30243
rect 2237 30209 2271 30243
rect 23397 30209 23431 30243
rect 24409 30209 24443 30243
rect 25145 30209 25179 30243
rect 27537 30209 27571 30243
rect 37841 30209 37875 30243
rect 24593 30141 24627 30175
rect 22385 30073 22419 30107
rect 23949 30073 23983 30107
rect 1501 30005 1535 30039
rect 23305 30005 23339 30039
rect 25789 30005 25823 30039
rect 26985 30005 27019 30039
rect 27721 30005 27755 30039
rect 38025 30005 38059 30039
rect 20637 29801 20671 29835
rect 23765 29801 23799 29835
rect 27537 29801 27571 29835
rect 34897 29801 34931 29835
rect 22109 29665 22143 29699
rect 26985 29665 27019 29699
rect 1685 29597 1719 29631
rect 20453 29597 20487 29631
rect 22385 29597 22419 29631
rect 34713 29597 34747 29631
rect 37473 29597 37507 29631
rect 38117 29597 38151 29631
rect 24777 29529 24811 29563
rect 25513 29529 25547 29563
rect 1501 29461 1535 29495
rect 22845 29461 22879 29495
rect 26157 29461 26191 29495
rect 27077 29461 27111 29495
rect 27169 29461 27203 29495
rect 27997 29461 28031 29495
rect 37933 29461 37967 29495
rect 19809 29257 19843 29291
rect 22201 29257 22235 29291
rect 27077 29257 27111 29291
rect 34253 29257 34287 29291
rect 16037 29189 16071 29223
rect 22661 29189 22695 29223
rect 24041 29189 24075 29223
rect 33885 29189 33919 29223
rect 1409 29121 1443 29155
rect 2053 29121 2087 29155
rect 15485 29121 15519 29155
rect 20269 29121 20303 29155
rect 22569 29121 22603 29155
rect 37473 29121 37507 29155
rect 38117 29121 38151 29155
rect 16681 29053 16715 29087
rect 20545 29053 20579 29087
rect 22753 29053 22787 29087
rect 33609 29053 33643 29087
rect 33793 29053 33827 29087
rect 1593 28985 1627 29019
rect 23397 28985 23431 29019
rect 32965 28985 32999 29019
rect 37933 28985 37967 29019
rect 20821 28713 20855 28747
rect 33425 28713 33459 28747
rect 21373 28577 21407 28611
rect 22017 28509 22051 28543
rect 21189 28441 21223 28475
rect 22201 28441 22235 28475
rect 4997 28373 5031 28407
rect 19625 28373 19659 28407
rect 20177 28373 20211 28407
rect 21281 28373 21315 28407
rect 22753 28373 22787 28407
rect 1593 28169 1627 28203
rect 4445 28169 4479 28203
rect 4537 28169 4571 28203
rect 5365 28169 5399 28203
rect 19349 28169 19383 28203
rect 20361 28169 20395 28203
rect 21925 28169 21959 28203
rect 22293 28169 22327 28203
rect 20729 28101 20763 28135
rect 1409 28033 1443 28067
rect 2053 28033 2087 28067
rect 19901 28033 19935 28067
rect 20821 28033 20855 28067
rect 25605 28033 25639 28067
rect 37841 28033 37875 28067
rect 4353 27965 4387 27999
rect 20913 27965 20947 27999
rect 22385 27965 22419 27999
rect 22477 27965 22511 27999
rect 23121 27965 23155 27999
rect 25973 27965 26007 27999
rect 37289 27897 37323 27931
rect 38025 27897 38059 27931
rect 4905 27829 4939 27863
rect 23673 27829 23707 27863
rect 27077 27829 27111 27863
rect 21465 27625 21499 27659
rect 23029 27625 23063 27659
rect 1593 27557 1627 27591
rect 21005 27557 21039 27591
rect 22385 27557 22419 27591
rect 19809 27489 19843 27523
rect 21557 27489 21591 27523
rect 1409 27421 1443 27455
rect 2053 27421 2087 27455
rect 5273 27421 5307 27455
rect 21465 27421 21499 27455
rect 21741 27421 21775 27455
rect 37841 27421 37875 27455
rect 5457 27353 5491 27387
rect 18705 27353 18739 27387
rect 20085 27353 20119 27387
rect 19993 27285 20027 27319
rect 20453 27285 20487 27319
rect 21925 27285 21959 27319
rect 37289 27285 37323 27319
rect 38025 27285 38059 27319
rect 18981 27081 19015 27115
rect 22477 27081 22511 27115
rect 1685 26945 1719 26979
rect 2237 26945 2271 26979
rect 20085 26945 20119 26979
rect 20729 26945 20763 26979
rect 21833 26945 21867 26979
rect 37473 26945 37507 26979
rect 38117 26945 38151 26979
rect 21005 26877 21039 26911
rect 20269 26809 20303 26843
rect 1501 26741 1535 26775
rect 19533 26741 19567 26775
rect 23213 26741 23247 26775
rect 37933 26741 37967 26775
rect 18613 26537 18647 26571
rect 20913 26537 20947 26571
rect 22753 26537 22787 26571
rect 22293 26469 22327 26503
rect 38025 26469 38059 26503
rect 1685 26333 1719 26367
rect 21833 26333 21867 26367
rect 22477 26333 22511 26367
rect 22845 26333 22879 26367
rect 27261 26333 27295 26367
rect 37381 26333 37415 26367
rect 37841 26333 37875 26367
rect 1501 26197 1535 26231
rect 23397 26197 23431 26231
rect 27445 26197 27479 26231
rect 19625 25993 19659 26027
rect 20913 25993 20947 26027
rect 23857 25993 23891 26027
rect 26433 25993 26467 26027
rect 27353 25993 27387 26027
rect 27721 25993 27755 26027
rect 18153 25857 18187 25891
rect 19073 25857 19107 25891
rect 22661 25857 22695 25891
rect 22753 25857 22787 25891
rect 18429 25789 18463 25823
rect 22477 25789 22511 25823
rect 22569 25789 22603 25823
rect 27077 25789 27111 25823
rect 27261 25789 27295 25823
rect 23397 25721 23431 25755
rect 1685 25653 1719 25687
rect 20361 25653 20395 25687
rect 22293 25653 22327 25687
rect 25513 25449 25547 25483
rect 37933 25449 37967 25483
rect 24409 25381 24443 25415
rect 19717 25313 19751 25347
rect 19901 25313 19935 25347
rect 21649 25313 21683 25347
rect 21741 25313 21775 25347
rect 22937 25313 22971 25347
rect 1869 25245 1903 25279
rect 17877 25245 17911 25279
rect 19625 25245 19659 25279
rect 23213 25245 23247 25279
rect 23765 25245 23799 25279
rect 37473 25245 37507 25279
rect 38117 25245 38151 25279
rect 2053 25177 2087 25211
rect 18245 25177 18279 25211
rect 25053 25177 25087 25211
rect 19257 25109 19291 25143
rect 20729 25109 20763 25143
rect 21189 25109 21223 25143
rect 21557 25109 21591 25143
rect 26801 25109 26835 25143
rect 22017 24905 22051 24939
rect 22845 24905 22879 24939
rect 23673 24905 23707 24939
rect 1409 24769 1443 24803
rect 2053 24769 2087 24803
rect 17969 24769 18003 24803
rect 19257 24769 19291 24803
rect 21281 24769 21315 24803
rect 21833 24769 21867 24803
rect 24041 24769 24075 24803
rect 25329 24769 25363 24803
rect 37473 24769 37507 24803
rect 38117 24769 38151 24803
rect 18981 24701 19015 24735
rect 21005 24701 21039 24735
rect 22569 24701 22603 24735
rect 22753 24701 22787 24735
rect 24133 24701 24167 24735
rect 24225 24701 24259 24735
rect 25881 24701 25915 24735
rect 1593 24633 1627 24667
rect 19901 24633 19935 24667
rect 37933 24633 37967 24667
rect 23213 24565 23247 24599
rect 27905 24565 27939 24599
rect 18521 24361 18555 24395
rect 19349 24361 19383 24395
rect 23673 24361 23707 24395
rect 24777 24361 24811 24395
rect 29653 24361 29687 24395
rect 21649 24293 21683 24327
rect 23489 24293 23523 24327
rect 17601 24225 17635 24259
rect 20177 24225 20211 24259
rect 21465 24225 21499 24259
rect 23029 24225 23063 24259
rect 24685 24225 24719 24259
rect 25881 24225 25915 24259
rect 28089 24225 28123 24259
rect 28273 24225 28307 24259
rect 13553 24157 13587 24191
rect 17049 24157 17083 24191
rect 18337 24157 18371 24191
rect 18521 24157 18555 24191
rect 19901 24157 19935 24191
rect 21741 24157 21775 24191
rect 22753 24157 22787 24191
rect 24593 24157 24627 24191
rect 24869 24157 24903 24191
rect 37841 24157 37875 24191
rect 1869 24089 1903 24123
rect 2053 24089 2087 24123
rect 18061 24089 18095 24123
rect 23857 24089 23891 24123
rect 27445 24089 27479 24123
rect 28365 24089 28399 24123
rect 2513 24021 2547 24055
rect 13369 24021 13403 24055
rect 18705 24021 18739 24055
rect 21741 24021 21775 24055
rect 23647 24021 23681 24055
rect 24409 24021 24443 24055
rect 25329 24021 25363 24055
rect 28733 24021 28767 24055
rect 38025 24021 38059 24055
rect 13645 23817 13679 23851
rect 21833 23817 21867 23851
rect 24501 23817 24535 23851
rect 27629 23817 27663 23851
rect 28457 23817 28491 23851
rect 29469 23817 29503 23851
rect 37381 23817 37415 23851
rect 2237 23749 2271 23783
rect 17601 23749 17635 23783
rect 18061 23749 18095 23783
rect 1685 23681 1719 23715
rect 14013 23681 14047 23715
rect 21097 23681 21131 23715
rect 21281 23681 21315 23715
rect 22201 23681 22235 23715
rect 23121 23681 23155 23715
rect 29285 23681 29319 23715
rect 37841 23681 37875 23715
rect 13185 23613 13219 23647
rect 14105 23613 14139 23647
rect 14289 23613 14323 23647
rect 18889 23613 18923 23647
rect 19441 23613 19475 23647
rect 19717 23613 19751 23647
rect 22293 23613 22327 23647
rect 22385 23613 22419 23647
rect 23397 23613 23431 23647
rect 28181 23613 28215 23647
rect 28365 23613 28399 23647
rect 21281 23545 21315 23579
rect 28825 23545 28859 23579
rect 1501 23477 1535 23511
rect 14933 23477 14967 23511
rect 24961 23477 24995 23511
rect 29929 23477 29963 23511
rect 38025 23477 38059 23511
rect 18613 23273 18647 23307
rect 19257 23273 19291 23307
rect 20453 23273 20487 23307
rect 24501 23273 24535 23307
rect 27905 23273 27939 23307
rect 23489 23205 23523 23239
rect 10333 23137 10367 23171
rect 19717 23137 19751 23171
rect 19901 23137 19935 23171
rect 21005 23137 21039 23171
rect 22293 23137 22327 23171
rect 22477 23137 22511 23171
rect 10057 23069 10091 23103
rect 16313 23069 16347 23103
rect 16589 23069 16623 23103
rect 28549 23069 28583 23103
rect 19625 23001 19659 23035
rect 22569 23001 22603 23035
rect 14565 22933 14599 22967
rect 20821 22933 20855 22967
rect 20913 22933 20947 22967
rect 21741 22933 21775 22967
rect 22937 22933 22971 22967
rect 28733 22933 28767 22967
rect 38117 22933 38151 22967
rect 10241 22729 10275 22763
rect 16681 22729 16715 22763
rect 18613 22729 18647 22763
rect 19257 22729 19291 22763
rect 20269 22729 20303 22763
rect 21189 22729 21223 22763
rect 21833 22729 21867 22763
rect 22477 22729 22511 22763
rect 23581 22729 23615 22763
rect 19717 22661 19751 22695
rect 24685 22661 24719 22695
rect 1409 22593 1443 22627
rect 2053 22593 2087 22627
rect 9781 22593 9815 22627
rect 10609 22593 10643 22627
rect 10701 22593 10735 22627
rect 11529 22593 11563 22627
rect 17049 22593 17083 22627
rect 22661 22593 22695 22627
rect 22753 22593 22787 22627
rect 22937 22593 22971 22627
rect 23397 22593 23431 22627
rect 10885 22525 10919 22559
rect 17141 22525 17175 22559
rect 17325 22525 17359 22559
rect 17969 22525 18003 22559
rect 25145 22525 25179 22559
rect 37841 22525 37875 22559
rect 38117 22525 38151 22559
rect 1593 22389 1627 22423
rect 22937 22389 22971 22423
rect 24133 22389 24167 22423
rect 37933 22117 37967 22151
rect 11161 22049 11195 22083
rect 20821 22049 20855 22083
rect 21005 22049 21039 22083
rect 21925 22049 21959 22083
rect 22477 22049 22511 22083
rect 1409 21981 1443 22015
rect 2053 21981 2087 22015
rect 37473 21981 37507 22015
rect 38117 21981 38151 22015
rect 19809 21913 19843 21947
rect 20729 21913 20763 21947
rect 1593 21845 1627 21879
rect 17601 21845 17635 21879
rect 20361 21845 20395 21879
rect 22937 21845 22971 21879
rect 23581 21845 23615 21879
rect 6929 21641 6963 21675
rect 1961 21505 1995 21539
rect 20453 21505 20487 21539
rect 37841 21505 37875 21539
rect 2237 21437 2271 21471
rect 20637 21301 20671 21335
rect 21281 21301 21315 21335
rect 38025 21301 38059 21335
rect 2053 21097 2087 21131
rect 37933 21097 37967 21131
rect 6193 20961 6227 20995
rect 1409 20893 1443 20927
rect 6469 20893 6503 20927
rect 37473 20893 37507 20927
rect 38117 20893 38151 20927
rect 6377 20825 6411 20859
rect 7389 20825 7423 20859
rect 1593 20757 1627 20791
rect 6837 20757 6871 20791
rect 7481 20757 7515 20791
rect 7113 20553 7147 20587
rect 32965 20553 32999 20587
rect 1409 20485 1443 20519
rect 3249 20417 3283 20451
rect 33885 20417 33919 20451
rect 3341 20349 3375 20383
rect 3525 20349 3559 20383
rect 33609 20349 33643 20383
rect 4169 20281 4203 20315
rect 2053 20213 2087 20247
rect 2881 20213 2915 20247
rect 12541 20213 12575 20247
rect 3893 20009 3927 20043
rect 12265 20009 12299 20043
rect 14197 20009 14231 20043
rect 21833 20009 21867 20043
rect 37289 19941 37323 19975
rect 13461 19873 13495 19907
rect 33241 19873 33275 19907
rect 1961 19805 1995 19839
rect 2237 19805 2271 19839
rect 2881 19805 2915 19839
rect 13277 19805 13311 19839
rect 33333 19805 33367 19839
rect 37841 19805 37875 19839
rect 32505 19737 32539 19771
rect 33425 19737 33459 19771
rect 2697 19669 2731 19703
rect 12817 19669 12851 19703
rect 13185 19669 13219 19703
rect 33793 19669 33827 19703
rect 38025 19669 38059 19703
rect 3341 19465 3375 19499
rect 33793 19465 33827 19499
rect 23121 19397 23155 19431
rect 1685 19329 1719 19363
rect 3525 19329 3559 19363
rect 12725 19329 12759 19363
rect 22293 19329 22327 19363
rect 22385 19329 22419 19363
rect 33425 19329 33459 19363
rect 34253 19329 34287 19363
rect 22477 19261 22511 19295
rect 33149 19261 33183 19295
rect 33333 19261 33367 19295
rect 32505 19193 32539 19227
rect 1501 19125 1535 19159
rect 12541 19125 12575 19159
rect 21925 19125 21959 19159
rect 23765 19125 23799 19159
rect 34437 19125 34471 19159
rect 32965 18921 32999 18955
rect 21373 18785 21407 18819
rect 1685 18717 1719 18751
rect 21649 18717 21683 18751
rect 37841 18717 37875 18751
rect 1501 18581 1535 18615
rect 33885 18581 33919 18615
rect 38025 18581 38059 18615
rect 14289 18377 14323 18411
rect 25145 18377 25179 18411
rect 2237 18309 2271 18343
rect 1685 18241 1719 18275
rect 13001 18241 13035 18275
rect 26065 18241 26099 18275
rect 26985 18241 27019 18275
rect 37473 18241 37507 18275
rect 38117 18241 38151 18275
rect 25789 18173 25823 18207
rect 25973 18173 26007 18207
rect 37933 18105 37967 18139
rect 1501 18037 1535 18071
rect 26433 18037 26467 18071
rect 3801 17833 3835 17867
rect 16037 17765 16071 17799
rect 4445 17697 4479 17731
rect 26525 17629 26559 17663
rect 36737 17629 36771 17663
rect 38117 17629 38151 17663
rect 14749 17561 14783 17595
rect 4169 17493 4203 17527
rect 4261 17493 4295 17527
rect 4997 17493 5031 17527
rect 14197 17493 14231 17527
rect 26709 17493 26743 17527
rect 37289 17493 37323 17527
rect 37933 17493 37967 17527
rect 1593 17289 1627 17323
rect 4629 17289 4663 17323
rect 37657 17289 37691 17323
rect 37749 17289 37783 17323
rect 36737 17221 36771 17255
rect 1409 17153 1443 17187
rect 2053 17153 2087 17187
rect 37473 17085 37507 17119
rect 38117 16949 38151 16983
rect 1961 16609 1995 16643
rect 25145 16609 25179 16643
rect 25881 16609 25915 16643
rect 25973 16609 26007 16643
rect 36737 16609 36771 16643
rect 2237 16541 2271 16575
rect 26893 16541 26927 16575
rect 37381 16541 37415 16575
rect 38025 16541 38059 16575
rect 26065 16405 26099 16439
rect 26433 16405 26467 16439
rect 27077 16405 27111 16439
rect 37197 16405 37231 16439
rect 37841 16405 37875 16439
rect 2053 16201 2087 16235
rect 26985 16201 27019 16235
rect 37381 16201 37415 16235
rect 1409 16065 1443 16099
rect 15117 16065 15151 16099
rect 37841 16065 37875 16099
rect 14933 15997 14967 16031
rect 15025 15997 15059 16031
rect 1593 15929 1627 15963
rect 14197 15861 14231 15895
rect 15485 15861 15519 15895
rect 16037 15861 16071 15895
rect 38025 15861 38059 15895
rect 1409 15657 1443 15691
rect 15485 15521 15519 15555
rect 15761 15453 15795 15487
rect 37473 15453 37507 15487
rect 38117 15453 38151 15487
rect 37933 15317 37967 15351
rect 27353 15113 27387 15147
rect 34805 15113 34839 15147
rect 28273 15045 28307 15079
rect 4813 14977 4847 15011
rect 34621 14977 34655 15011
rect 28365 14909 28399 14943
rect 28457 14909 28491 14943
rect 4997 14841 5031 14875
rect 27905 14773 27939 14807
rect 38117 14773 38151 14807
rect 26801 14569 26835 14603
rect 27353 14433 27387 14467
rect 37841 14433 37875 14467
rect 1685 14365 1719 14399
rect 2237 14365 2271 14399
rect 27629 14365 27663 14399
rect 38117 14365 38151 14399
rect 1501 14229 1535 14263
rect 33701 14229 33735 14263
rect 4813 14025 4847 14059
rect 33241 14025 33275 14059
rect 34161 14025 34195 14059
rect 34253 14025 34287 14059
rect 34989 14025 35023 14059
rect 1961 13889 1995 13923
rect 4629 13889 4663 13923
rect 27353 13889 27387 13923
rect 37841 13889 37875 13923
rect 2237 13821 2271 13855
rect 26341 13821 26375 13855
rect 27445 13821 27479 13855
rect 27537 13821 27571 13855
rect 34437 13821 34471 13855
rect 26985 13685 27019 13719
rect 33793 13685 33827 13719
rect 38025 13685 38059 13719
rect 2053 13481 2087 13515
rect 4537 13481 4571 13515
rect 34713 13481 34747 13515
rect 37289 13413 37323 13447
rect 3985 13345 4019 13379
rect 35265 13345 35299 13379
rect 1409 13277 1443 13311
rect 2605 13277 2639 13311
rect 4169 13277 4203 13311
rect 26893 13277 26927 13311
rect 33977 13277 34011 13311
rect 35173 13277 35207 13311
rect 37841 13277 37875 13311
rect 4077 13209 4111 13243
rect 1593 13141 1627 13175
rect 4997 13141 5031 13175
rect 27077 13141 27111 13175
rect 34161 13141 34195 13175
rect 35081 13141 35115 13175
rect 38025 13141 38059 13175
rect 13001 12869 13035 12903
rect 1685 12801 1719 12835
rect 37841 12801 37875 12835
rect 38117 12733 38151 12767
rect 1501 12597 1535 12631
rect 14289 12597 14323 12631
rect 34529 12597 34563 12631
rect 10609 12393 10643 12427
rect 38117 12325 38151 12359
rect 11805 12257 11839 12291
rect 10793 12189 10827 12223
rect 1501 12053 1535 12087
rect 11253 12053 11287 12087
rect 11621 12053 11655 12087
rect 11713 12053 11747 12087
rect 37473 12053 37507 12087
rect 4077 11849 4111 11883
rect 4537 11849 4571 11883
rect 2053 11781 2087 11815
rect 11529 11781 11563 11815
rect 1501 11713 1535 11747
rect 4169 11713 4203 11747
rect 14841 11713 14875 11747
rect 3893 11645 3927 11679
rect 10885 11645 10919 11679
rect 14565 11645 14599 11679
rect 37289 11645 37323 11679
rect 37565 11645 37599 11679
rect 4997 11509 5031 11543
rect 1593 11305 1627 11339
rect 37933 11305 37967 11339
rect 1409 11101 1443 11135
rect 2053 11101 2087 11135
rect 37473 11101 37507 11135
rect 38117 11101 38151 11135
rect 8309 10761 8343 10795
rect 7757 10693 7791 10727
rect 9045 10693 9079 10727
rect 15577 10693 15611 10727
rect 1409 10625 1443 10659
rect 2053 10625 2087 10659
rect 9137 10625 9171 10659
rect 14749 10625 14783 10659
rect 37473 10625 37507 10659
rect 38117 10625 38151 10659
rect 8861 10557 8895 10591
rect 14565 10557 14599 10591
rect 14657 10557 14691 10591
rect 13829 10489 13863 10523
rect 37933 10489 37967 10523
rect 1593 10421 1627 10455
rect 9505 10421 9539 10455
rect 15117 10421 15151 10455
rect 37933 10217 37967 10251
rect 12357 10149 12391 10183
rect 1409 10013 1443 10047
rect 2053 10013 2087 10047
rect 12173 10013 12207 10047
rect 15853 10013 15887 10047
rect 37381 10013 37415 10047
rect 38117 10013 38151 10047
rect 1593 9877 1627 9911
rect 16037 9877 16071 9911
rect 15485 9537 15519 9571
rect 14657 9469 14691 9503
rect 15577 9469 15611 9503
rect 15669 9469 15703 9503
rect 15117 9401 15151 9435
rect 16773 9333 16807 9367
rect 38117 9333 38151 9367
rect 37841 8993 37875 9027
rect 1685 8925 1719 8959
rect 38117 8925 38151 8959
rect 2237 8857 2271 8891
rect 1501 8789 1535 8823
rect 15669 8585 15703 8619
rect 1961 8449 1995 8483
rect 15761 8449 15795 8483
rect 37289 8449 37323 8483
rect 37841 8449 37875 8483
rect 2237 8381 2271 8415
rect 2697 8381 2731 8415
rect 15577 8381 15611 8415
rect 16773 8313 16807 8347
rect 38025 8313 38059 8347
rect 16129 8245 16163 8279
rect 1961 7905 1995 7939
rect 16313 7905 16347 7939
rect 2237 7837 2271 7871
rect 16589 7837 16623 7871
rect 37841 7837 37875 7871
rect 38025 7701 38059 7735
rect 2053 7497 2087 7531
rect 1409 7361 1443 7395
rect 22569 7361 22603 7395
rect 37381 7361 37415 7395
rect 38025 7361 38059 7395
rect 37841 7293 37875 7327
rect 1593 7225 1627 7259
rect 22753 7225 22787 7259
rect 1409 6885 1443 6919
rect 10609 6817 10643 6851
rect 12449 6817 12483 6851
rect 21925 6817 21959 6851
rect 21741 6749 21775 6783
rect 10793 6681 10827 6715
rect 21557 6681 21591 6715
rect 22477 6613 22511 6647
rect 11529 6409 11563 6443
rect 24225 6409 24259 6443
rect 37289 6409 37323 6443
rect 1685 6273 1719 6307
rect 2145 6273 2179 6307
rect 11897 6273 11931 6307
rect 13829 6273 13863 6307
rect 14749 6273 14783 6307
rect 37841 6273 37875 6307
rect 11989 6205 12023 6239
rect 12173 6205 12207 6239
rect 13921 6205 13955 6239
rect 14105 6205 14139 6239
rect 1501 6137 1535 6171
rect 38025 6137 38059 6171
rect 12817 6069 12851 6103
rect 13461 6069 13495 6103
rect 14381 5865 14415 5899
rect 25605 5865 25639 5899
rect 7205 5797 7239 5831
rect 2237 5729 2271 5763
rect 6561 5729 6595 5763
rect 24961 5729 24995 5763
rect 26617 5729 26651 5763
rect 1685 5661 1719 5695
rect 5549 5661 5583 5695
rect 6377 5661 6411 5695
rect 13001 5661 13035 5695
rect 26893 5661 26927 5695
rect 37841 5661 37875 5695
rect 6469 5593 6503 5627
rect 24777 5593 24811 5627
rect 26801 5593 26835 5627
rect 27813 5593 27847 5627
rect 1501 5525 1535 5559
rect 2789 5525 2823 5559
rect 6009 5525 6043 5559
rect 12817 5525 12851 5559
rect 23765 5525 23799 5559
rect 24409 5525 24443 5559
rect 24869 5525 24903 5559
rect 27261 5525 27295 5559
rect 37381 5525 37415 5559
rect 38025 5525 38059 5559
rect 1593 5321 1627 5355
rect 26341 5321 26375 5355
rect 37381 5321 37415 5355
rect 1409 5185 1443 5219
rect 2053 5185 2087 5219
rect 5825 5185 5859 5219
rect 23673 5185 23707 5219
rect 27077 5185 27111 5219
rect 37841 5185 37875 5219
rect 2605 4981 2639 5015
rect 3157 4981 3191 5015
rect 5641 4981 5675 5015
rect 23857 4981 23891 5015
rect 27261 4981 27295 5015
rect 36645 4981 36679 5015
rect 38025 4981 38059 5015
rect 2145 4777 2179 4811
rect 36185 4777 36219 4811
rect 37841 4709 37875 4743
rect 1685 4573 1719 4607
rect 17601 4573 17635 4607
rect 37381 4505 37415 4539
rect 38025 4505 38059 4539
rect 1501 4437 1535 4471
rect 2789 4437 2823 4471
rect 3893 4437 3927 4471
rect 15577 4437 15611 4471
rect 17785 4437 17819 4471
rect 35725 4437 35759 4471
rect 36737 4437 36771 4471
rect 38025 4165 38059 4199
rect 1409 4097 1443 4131
rect 2053 4097 2087 4131
rect 24501 4097 24535 4131
rect 30849 4097 30883 4131
rect 37289 4097 37323 4131
rect 15485 4029 15519 4063
rect 1593 3961 1627 3995
rect 2237 3961 2271 3995
rect 37841 3961 37875 3995
rect 2697 3893 2731 3927
rect 3709 3893 3743 3927
rect 4169 3893 4203 3927
rect 4721 3893 4755 3927
rect 16129 3893 16163 3927
rect 35449 3893 35483 3927
rect 36093 3893 36127 3927
rect 36553 3893 36587 3927
rect 3985 3689 4019 3723
rect 5641 3689 5675 3723
rect 13461 3689 13495 3723
rect 14381 3689 14415 3723
rect 17969 3689 18003 3723
rect 30481 3689 30515 3723
rect 31033 3689 31067 3723
rect 33885 3689 33919 3723
rect 2881 3621 2915 3655
rect 35725 3621 35759 3655
rect 37289 3621 37323 3655
rect 1961 3553 1995 3587
rect 2237 3553 2271 3587
rect 15393 3553 15427 3587
rect 17325 3553 17359 3587
rect 17509 3553 17543 3587
rect 2697 3485 2731 3519
rect 3801 3485 3835 3519
rect 15660 3485 15694 3519
rect 24593 3485 24627 3519
rect 28457 3485 28491 3519
rect 31217 3485 31251 3519
rect 31677 3485 31711 3519
rect 35909 3485 35943 3519
rect 36369 3485 36403 3519
rect 37105 3485 37139 3519
rect 37841 3485 37875 3519
rect 18429 3417 18463 3451
rect 4905 3349 4939 3383
rect 6193 3349 6227 3383
rect 11621 3349 11655 3383
rect 14933 3349 14967 3383
rect 16773 3349 16807 3383
rect 17601 3349 17635 3383
rect 21373 3349 21407 3383
rect 23213 3349 23247 3383
rect 23673 3349 23707 3383
rect 24777 3349 24811 3383
rect 26801 3349 26835 3383
rect 27353 3349 27387 3383
rect 27905 3349 27939 3383
rect 32229 3349 32263 3383
rect 32781 3349 32815 3383
rect 33333 3349 33367 3383
rect 34713 3349 34747 3383
rect 36553 3349 36587 3383
rect 38025 3349 38059 3383
rect 2329 3145 2363 3179
rect 8493 3145 8527 3179
rect 9781 3145 9815 3179
rect 10425 3145 10459 3179
rect 11713 3145 11747 3179
rect 13185 3145 13219 3179
rect 15301 3145 15335 3179
rect 17509 3145 17543 3179
rect 18797 3145 18831 3179
rect 20545 3145 20579 3179
rect 21281 3145 21315 3179
rect 24961 3145 24995 3179
rect 25973 3145 26007 3179
rect 26985 3145 27019 3179
rect 27629 3145 27663 3179
rect 28457 3145 28491 3179
rect 31585 3145 31619 3179
rect 33425 3145 33459 3179
rect 34437 3145 34471 3179
rect 36553 3145 36587 3179
rect 3157 3077 3191 3111
rect 4813 3077 4847 3111
rect 14166 3077 14200 3111
rect 30389 3077 30423 3111
rect 31217 3077 31251 3111
rect 2237 3009 2271 3043
rect 2973 3009 3007 3043
rect 3617 3009 3651 3043
rect 4629 3009 4663 3043
rect 5549 3009 5583 3043
rect 6745 3009 6779 3043
rect 7205 3009 7239 3043
rect 8677 3009 8711 3043
rect 11529 3009 11563 3043
rect 12541 3009 12575 3043
rect 13001 3009 13035 3043
rect 13921 3009 13955 3043
rect 15761 3009 15795 3043
rect 17693 3009 17727 3043
rect 18153 3009 18187 3043
rect 18981 3009 19015 3043
rect 19441 3009 19475 3043
rect 21097 3009 21131 3043
rect 22109 3009 22143 3043
rect 25789 3009 25823 3043
rect 27169 3009 27203 3043
rect 27813 3009 27847 3043
rect 28641 3009 28675 3043
rect 29101 3009 29135 3043
rect 32137 3009 32171 3043
rect 32965 3009 32999 3043
rect 33609 3009 33643 3043
rect 34253 3009 34287 3043
rect 35265 3009 35299 3043
rect 35725 3009 35759 3043
rect 36645 3009 36679 3043
rect 37473 3009 37507 3043
rect 23305 2941 23339 2975
rect 23581 2941 23615 2975
rect 24685 2941 24719 2975
rect 24869 2941 24903 2975
rect 30941 2941 30975 2975
rect 31125 2941 31159 2975
rect 3801 2873 3835 2907
rect 7389 2873 7423 2907
rect 15945 2873 15979 2907
rect 25329 2873 25363 2907
rect 32781 2873 32815 2907
rect 1593 2805 1627 2839
rect 5365 2805 5399 2839
rect 8033 2805 8067 2839
rect 9229 2805 9263 2839
rect 10977 2805 11011 2839
rect 16681 2805 16715 2839
rect 21925 2805 21959 2839
rect 22569 2805 22603 2839
rect 29653 2805 29687 2839
rect 32321 2805 32355 2839
rect 35081 2805 35115 2839
rect 35909 2805 35943 2839
rect 37657 2805 37691 2839
rect 8033 2601 8067 2635
rect 9137 2601 9171 2635
rect 15485 2601 15519 2635
rect 15945 2601 15979 2635
rect 24409 2601 24443 2635
rect 26985 2601 27019 2635
rect 27629 2601 27663 2635
rect 28273 2601 28307 2635
rect 35817 2601 35851 2635
rect 25789 2533 25823 2567
rect 28917 2533 28951 2567
rect 36461 2533 36495 2567
rect 1961 2465 1995 2499
rect 3985 2465 4019 2499
rect 4261 2465 4295 2499
rect 11989 2465 12023 2499
rect 22293 2465 22327 2499
rect 25053 2465 25087 2499
rect 26341 2465 26375 2499
rect 32413 2465 32447 2499
rect 37289 2465 37323 2499
rect 2237 2397 2271 2431
rect 3249 2397 3283 2431
rect 5641 2397 5675 2431
rect 6837 2397 6871 2431
rect 9965 2397 9999 2431
rect 10701 2397 10735 2431
rect 11713 2397 11747 2431
rect 13277 2397 13311 2431
rect 14381 2397 14415 2431
rect 15301 2397 15335 2431
rect 16129 2397 16163 2431
rect 17141 2397 17175 2431
rect 17693 2397 17727 2431
rect 18153 2397 18187 2431
rect 19257 2397 19291 2431
rect 20269 2397 20303 2431
rect 20729 2397 20763 2431
rect 22017 2397 22051 2431
rect 25605 2397 25639 2431
rect 27169 2397 27203 2431
rect 27813 2397 27847 2431
rect 28457 2397 28491 2431
rect 29745 2397 29779 2431
rect 30021 2397 30055 2431
rect 31033 2397 31067 2431
rect 32137 2397 32171 2431
rect 33885 2397 33919 2431
rect 34897 2397 34931 2431
rect 36645 2397 36679 2431
rect 37565 2397 37599 2431
rect 7389 2329 7423 2363
rect 7941 2329 7975 2363
rect 9045 2329 9079 2363
rect 23489 2329 23523 2363
rect 24777 2329 24811 2363
rect 35909 2329 35943 2363
rect 3065 2261 3099 2295
rect 5733 2261 5767 2295
rect 6653 2261 6687 2295
rect 9781 2261 9815 2295
rect 10517 2261 10551 2295
rect 13093 2261 13127 2295
rect 14197 2261 14231 2295
rect 16957 2261 16991 2295
rect 18337 2261 18371 2295
rect 19441 2261 19475 2295
rect 20085 2261 20119 2295
rect 20913 2261 20947 2295
rect 23397 2261 23431 2295
rect 24869 2261 24903 2295
rect 31217 2261 31251 2295
rect 33701 2261 33735 2295
rect 35081 2261 35115 2295
<< metal1 >>
rect 13814 47472 13820 47524
rect 13872 47512 13878 47524
rect 20070 47512 20076 47524
rect 13872 47484 20076 47512
rect 13872 47472 13878 47484
rect 20070 47472 20076 47484
rect 20128 47472 20134 47524
rect 14 47404 20 47456
rect 72 47444 78 47456
rect 934 47444 940 47456
rect 72 47416 940 47444
rect 72 47404 78 47416
rect 934 47404 940 47416
rect 992 47404 998 47456
rect 10962 47404 10968 47456
rect 11020 47444 11026 47456
rect 24302 47444 24308 47456
rect 11020 47416 24308 47444
rect 11020 47404 11026 47416
rect 24302 47404 24308 47416
rect 24360 47404 24366 47456
rect 1104 47354 38824 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 38824 47354
rect 1104 47280 38824 47302
rect 4614 47240 4620 47252
rect 4575 47212 4620 47240
rect 4614 47200 4620 47212
rect 4672 47200 4678 47252
rect 9858 47240 9864 47252
rect 4908 47212 6914 47240
rect 9819 47212 9864 47240
rect 2961 47175 3019 47181
rect 2961 47141 2973 47175
rect 3007 47172 3019 47175
rect 4908 47172 4936 47212
rect 3007 47144 4936 47172
rect 3007 47141 3019 47144
rect 2961 47135 3019 47141
rect 6454 47132 6460 47184
rect 6512 47172 6518 47184
rect 6733 47175 6791 47181
rect 6733 47172 6745 47175
rect 6512 47144 6745 47172
rect 6512 47132 6518 47144
rect 6733 47141 6745 47144
rect 6779 47141 6791 47175
rect 6886 47172 6914 47212
rect 9858 47200 9864 47212
rect 9916 47200 9922 47252
rect 10962 47240 10968 47252
rect 10923 47212 10968 47240
rect 10962 47200 10968 47212
rect 11020 47200 11026 47252
rect 13449 47243 13507 47249
rect 13449 47209 13461 47243
rect 13495 47240 13507 47243
rect 14458 47240 14464 47252
rect 13495 47212 14464 47240
rect 13495 47209 13507 47212
rect 13449 47203 13507 47209
rect 14458 47200 14464 47212
rect 14516 47200 14522 47252
rect 15933 47243 15991 47249
rect 15933 47209 15945 47243
rect 15979 47240 15991 47243
rect 16758 47240 16764 47252
rect 15979 47212 16764 47240
rect 15979 47209 15991 47212
rect 15933 47203 15991 47209
rect 16758 47200 16764 47212
rect 16816 47200 16822 47252
rect 17954 47200 17960 47252
rect 18012 47240 18018 47252
rect 18141 47243 18199 47249
rect 18141 47240 18153 47243
rect 18012 47212 18153 47240
rect 18012 47200 18018 47212
rect 18141 47209 18153 47212
rect 18187 47209 18199 47243
rect 20070 47240 20076 47252
rect 20031 47212 20076 47240
rect 18141 47203 18199 47209
rect 20070 47200 20076 47212
rect 20128 47200 20134 47252
rect 20714 47200 20720 47252
rect 20772 47240 20778 47252
rect 20901 47243 20959 47249
rect 20901 47240 20913 47243
rect 20772 47212 20913 47240
rect 20772 47200 20778 47212
rect 20901 47209 20913 47212
rect 20947 47209 20959 47243
rect 22462 47240 22468 47252
rect 22423 47212 22468 47240
rect 20901 47203 20959 47209
rect 22462 47200 22468 47212
rect 22520 47200 22526 47252
rect 26418 47200 26424 47252
rect 26476 47240 26482 47252
rect 27157 47243 27215 47249
rect 27157 47240 27169 47243
rect 26476 47212 27169 47240
rect 26476 47200 26482 47212
rect 27157 47209 27169 47212
rect 27203 47209 27215 47243
rect 27157 47203 27215 47209
rect 27338 47200 27344 47252
rect 27396 47240 27402 47252
rect 27893 47243 27951 47249
rect 27893 47240 27905 47243
rect 27396 47212 27905 47240
rect 27396 47200 27402 47212
rect 27893 47209 27905 47212
rect 27939 47209 27951 47243
rect 27893 47203 27951 47209
rect 30374 47200 30380 47252
rect 30432 47240 30438 47252
rect 30561 47243 30619 47249
rect 30561 47240 30573 47243
rect 30432 47212 30573 47240
rect 30432 47200 30438 47212
rect 30561 47209 30573 47212
rect 30607 47209 30619 47243
rect 30561 47203 30619 47209
rect 30926 47200 30932 47252
rect 30984 47240 30990 47252
rect 31297 47243 31355 47249
rect 31297 47240 31309 47243
rect 30984 47212 31309 47240
rect 30984 47200 30990 47212
rect 31297 47209 31309 47212
rect 31343 47209 31355 47243
rect 31297 47203 31355 47209
rect 31754 47200 31760 47252
rect 31812 47240 31818 47252
rect 32309 47243 32367 47249
rect 32309 47240 32321 47243
rect 31812 47212 32321 47240
rect 31812 47200 31818 47212
rect 32309 47209 32321 47212
rect 32355 47209 32367 47243
rect 36630 47240 36636 47252
rect 36591 47212 36636 47240
rect 32309 47203 32367 47209
rect 36630 47200 36636 47212
rect 36688 47200 36694 47252
rect 6886 47144 18000 47172
rect 6733 47135 6791 47141
rect 1489 47107 1547 47113
rect 1489 47073 1501 47107
rect 1535 47104 1547 47107
rect 7190 47104 7196 47116
rect 1535 47076 3280 47104
rect 1535 47073 1547 47076
rect 1489 47067 1547 47073
rect 3252 47048 3280 47076
rect 4632 47076 6914 47104
rect 7151 47076 7196 47104
rect 2038 47036 2044 47048
rect 1999 47008 2044 47036
rect 2038 46996 2044 47008
rect 2096 47036 2102 47048
rect 2590 47036 2596 47048
rect 2096 47008 2596 47036
rect 2096 46996 2102 47008
rect 2590 46996 2596 47008
rect 2648 46996 2654 47048
rect 2700 47008 3188 47036
rect 2225 46971 2283 46977
rect 2225 46937 2237 46971
rect 2271 46968 2283 46971
rect 2700 46968 2728 47008
rect 2271 46940 2728 46968
rect 2777 46971 2835 46977
rect 2271 46937 2283 46940
rect 2225 46931 2283 46937
rect 2777 46937 2789 46971
rect 2823 46937 2835 46971
rect 3160 46968 3188 47008
rect 3234 46996 3240 47048
rect 3292 47036 3298 47048
rect 3881 47039 3939 47045
rect 3881 47036 3893 47039
rect 3292 47008 3893 47036
rect 3292 46996 3298 47008
rect 3881 47005 3893 47008
rect 3927 47005 3939 47039
rect 4632 47036 4660 47076
rect 4798 47036 4804 47048
rect 3881 46999 3939 47005
rect 4172 47008 4660 47036
rect 4759 47008 4804 47036
rect 3160 46940 3924 46968
rect 2777 46931 2835 46937
rect 2682 46860 2688 46912
rect 2740 46900 2746 46912
rect 2792 46900 2820 46931
rect 3786 46900 3792 46912
rect 2740 46872 3792 46900
rect 2740 46860 2746 46872
rect 3786 46860 3792 46872
rect 3844 46860 3850 46912
rect 3896 46900 3924 46940
rect 3970 46928 3976 46980
rect 4028 46968 4034 46980
rect 4065 46971 4123 46977
rect 4065 46968 4077 46971
rect 4028 46940 4077 46968
rect 4028 46928 4034 46940
rect 4065 46937 4077 46940
rect 4111 46937 4123 46971
rect 4065 46931 4123 46937
rect 4172 46900 4200 47008
rect 4798 46996 4804 47008
rect 4856 46996 4862 47048
rect 5350 47036 5356 47048
rect 5311 47008 5356 47036
rect 5350 46996 5356 47008
rect 5408 46996 5414 47048
rect 6546 47036 6552 47048
rect 6507 47008 6552 47036
rect 6546 46996 6552 47008
rect 6604 46996 6610 47048
rect 6886 47036 6914 47076
rect 7190 47064 7196 47076
rect 7248 47064 7254 47116
rect 7300 47076 12112 47104
rect 7300 47036 7328 47076
rect 7466 47036 7472 47048
rect 6886 47008 7328 47036
rect 7427 47008 7472 47036
rect 7466 46996 7472 47008
rect 7524 46996 7530 47048
rect 8386 46996 8392 47048
rect 8444 47036 8450 47048
rect 8938 47036 8944 47048
rect 8444 47008 8944 47036
rect 8444 46996 8450 47008
rect 8938 46996 8944 47008
rect 8996 47036 9002 47048
rect 9125 47039 9183 47045
rect 9125 47036 9137 47039
rect 8996 47008 9137 47036
rect 8996 46996 9002 47008
rect 9125 47005 9137 47008
rect 9171 47005 9183 47039
rect 10042 47036 10048 47048
rect 10003 47008 10048 47036
rect 9125 46999 9183 47005
rect 10042 46996 10048 47008
rect 10100 46996 10106 47048
rect 10778 47036 10784 47048
rect 10739 47008 10784 47036
rect 10778 46996 10784 47008
rect 10836 46996 10842 47048
rect 11974 47036 11980 47048
rect 11935 47008 11980 47036
rect 11974 46996 11980 47008
rect 12032 46996 12038 47048
rect 12084 47036 12112 47076
rect 12728 47076 13860 47104
rect 12434 47036 12440 47048
rect 12084 47008 12440 47036
rect 12434 46996 12440 47008
rect 12492 46996 12498 47048
rect 12618 47036 12624 47048
rect 12579 47008 12624 47036
rect 12618 46996 12624 47008
rect 12676 46996 12682 47048
rect 5534 46968 5540 46980
rect 5495 46940 5540 46968
rect 5534 46928 5540 46940
rect 5592 46928 5598 46980
rect 9214 46928 9220 46980
rect 9272 46968 9278 46980
rect 9309 46971 9367 46977
rect 9309 46968 9321 46971
rect 9272 46940 9321 46968
rect 9272 46928 9278 46940
rect 9309 46937 9321 46940
rect 9355 46937 9367 46971
rect 12728 46968 12756 47076
rect 13262 47036 13268 47048
rect 13223 47008 13268 47036
rect 13262 46996 13268 47008
rect 13320 46996 13326 47048
rect 13832 47036 13860 47076
rect 13906 47064 13912 47116
rect 13964 47104 13970 47116
rect 14274 47104 14280 47116
rect 13964 47076 14280 47104
rect 13964 47064 13970 47076
rect 14274 47064 14280 47076
rect 14332 47064 14338 47116
rect 15378 47104 15384 47116
rect 14476 47076 15384 47104
rect 14476 47036 14504 47076
rect 15378 47064 15384 47076
rect 15436 47064 15442 47116
rect 17972 47104 18000 47144
rect 18046 47132 18052 47184
rect 18104 47172 18110 47184
rect 19429 47175 19487 47181
rect 19429 47172 19441 47175
rect 18104 47144 19441 47172
rect 18104 47132 18110 47144
rect 19429 47141 19441 47144
rect 19475 47141 19487 47175
rect 26142 47172 26148 47184
rect 19429 47135 19487 47141
rect 20548 47144 26148 47172
rect 20438 47104 20444 47116
rect 16546 47076 17816 47104
rect 17972 47076 20444 47104
rect 13832 47008 14504 47036
rect 14553 47039 14611 47045
rect 14553 47005 14565 47039
rect 14599 47036 14611 47039
rect 14642 47036 14648 47048
rect 14599 47008 14648 47036
rect 14599 47005 14611 47008
rect 14553 46999 14611 47005
rect 14642 46996 14648 47008
rect 14700 46996 14706 47048
rect 16117 47039 16175 47045
rect 16117 47005 16129 47039
rect 16163 47036 16175 47039
rect 16546 47036 16574 47076
rect 16666 47036 16672 47048
rect 16163 47008 16574 47036
rect 16627 47008 16672 47036
rect 16163 47005 16175 47008
rect 16117 46999 16175 47005
rect 16666 46996 16672 47008
rect 16724 46996 16730 47048
rect 16942 47036 16948 47048
rect 16903 47008 16948 47036
rect 16942 46996 16948 47008
rect 17000 46996 17006 47048
rect 17402 46968 17408 46980
rect 9309 46931 9367 46937
rect 12176 46940 12756 46968
rect 12820 46940 17408 46968
rect 12176 46909 12204 46940
rect 12820 46909 12848 46940
rect 17402 46928 17408 46940
rect 17460 46928 17466 46980
rect 17788 46968 17816 47076
rect 20438 47064 20444 47076
rect 20496 47064 20502 47116
rect 17954 47036 17960 47048
rect 17915 47008 17960 47036
rect 17954 46996 17960 47008
rect 18012 46996 18018 47048
rect 19334 46996 19340 47048
rect 19392 47036 19398 47048
rect 19610 47036 19616 47048
rect 19392 47008 19616 47036
rect 19392 46996 19398 47008
rect 19610 46996 19616 47008
rect 19668 46996 19674 47048
rect 20254 47036 20260 47048
rect 20215 47008 20260 47036
rect 20254 46996 20260 47008
rect 20312 46996 20318 47048
rect 20548 46968 20576 47144
rect 26142 47132 26148 47144
rect 26200 47132 26206 47184
rect 27706 47132 27712 47184
rect 27764 47172 27770 47184
rect 28629 47175 28687 47181
rect 28629 47172 28641 47175
rect 27764 47144 28641 47172
rect 27764 47132 27770 47144
rect 28629 47141 28641 47144
rect 28675 47141 28687 47175
rect 28629 47135 28687 47141
rect 34790 47132 34796 47184
rect 34848 47172 34854 47184
rect 34848 47144 34928 47172
rect 34848 47132 34854 47144
rect 23014 47104 23020 47116
rect 22975 47076 23020 47104
rect 23014 47064 23020 47076
rect 23072 47064 23078 47116
rect 23842 47064 23848 47116
rect 23900 47104 23906 47116
rect 24394 47104 24400 47116
rect 23900 47076 24400 47104
rect 23900 47064 23906 47076
rect 24394 47064 24400 47076
rect 24452 47064 24458 47116
rect 24854 47064 24860 47116
rect 24912 47104 24918 47116
rect 32950 47104 32956 47116
rect 24912 47076 32260 47104
rect 32911 47076 32956 47104
rect 24912 47064 24918 47076
rect 20717 47039 20775 47045
rect 20717 47005 20729 47039
rect 20763 47036 20775 47039
rect 21082 47036 21088 47048
rect 20763 47008 21088 47036
rect 20763 47005 20775 47008
rect 20717 46999 20775 47005
rect 21082 46996 21088 47008
rect 21140 46996 21146 47048
rect 22281 47039 22339 47045
rect 22281 47005 22293 47039
rect 22327 47036 22339 47039
rect 22830 47036 22836 47048
rect 22327 47008 22836 47036
rect 22327 47005 22339 47008
rect 22281 46999 22339 47005
rect 22830 46996 22836 47008
rect 22888 46996 22894 47048
rect 23290 47036 23296 47048
rect 23251 47008 23296 47036
rect 23290 46996 23296 47008
rect 23348 46996 23354 47048
rect 24670 47036 24676 47048
rect 24631 47008 24676 47036
rect 24670 46996 24676 47008
rect 24728 46996 24734 47048
rect 26050 47036 26056 47048
rect 26011 47008 26056 47036
rect 26050 46996 26056 47008
rect 26108 46996 26114 47048
rect 26970 47036 26976 47048
rect 26931 47008 26976 47036
rect 26970 46996 26976 47008
rect 27028 46996 27034 47048
rect 27338 46996 27344 47048
rect 27396 47036 27402 47048
rect 27709 47039 27767 47045
rect 27709 47036 27721 47039
rect 27396 47008 27721 47036
rect 27396 46996 27402 47008
rect 27709 47005 27721 47008
rect 27755 47005 27767 47039
rect 27709 46999 27767 47005
rect 27890 46996 27896 47048
rect 27948 47036 27954 47048
rect 28445 47039 28503 47045
rect 28445 47036 28457 47039
rect 27948 47008 28457 47036
rect 27948 46996 27954 47008
rect 28445 47005 28457 47008
rect 28491 47005 28503 47039
rect 28445 46999 28503 47005
rect 28994 46996 29000 47048
rect 29052 47036 29058 47048
rect 29638 47036 29644 47048
rect 29052 47008 29644 47036
rect 29052 46996 29058 47008
rect 29638 46996 29644 47008
rect 29696 47036 29702 47048
rect 29733 47039 29791 47045
rect 29733 47036 29745 47039
rect 29696 47008 29745 47036
rect 29696 46996 29702 47008
rect 29733 47005 29745 47008
rect 29779 47005 29791 47039
rect 29733 46999 29791 47005
rect 30377 47039 30435 47045
rect 30377 47005 30389 47039
rect 30423 47005 30435 47039
rect 30377 46999 30435 47005
rect 17788 46940 20576 46968
rect 25406 46928 25412 46980
rect 25464 46968 25470 46980
rect 25869 46971 25927 46977
rect 25869 46968 25881 46971
rect 25464 46940 25881 46968
rect 25464 46928 25470 46940
rect 25869 46937 25881 46940
rect 25915 46937 25927 46971
rect 25869 46931 25927 46937
rect 27430 46928 27436 46980
rect 27488 46968 27494 46980
rect 30392 46968 30420 46999
rect 30926 46996 30932 47048
rect 30984 47036 30990 47048
rect 31113 47039 31171 47045
rect 31113 47036 31125 47039
rect 30984 47008 31125 47036
rect 30984 46996 30990 47008
rect 31113 47005 31125 47008
rect 31159 47005 31171 47039
rect 31113 46999 31171 47005
rect 31478 46996 31484 47048
rect 31536 47036 31542 47048
rect 32125 47039 32183 47045
rect 32125 47036 32137 47039
rect 31536 47008 32137 47036
rect 31536 46996 31542 47008
rect 32125 47005 32137 47008
rect 32171 47005 32183 47039
rect 32232 47036 32260 47076
rect 32950 47064 32956 47076
rect 33008 47064 33014 47116
rect 34900 47113 34928 47144
rect 34885 47107 34943 47113
rect 34885 47073 34897 47107
rect 34931 47073 34943 47107
rect 34885 47067 34943 47073
rect 35618 47064 35624 47116
rect 35676 47104 35682 47116
rect 37553 47107 37611 47113
rect 37553 47104 37565 47107
rect 35676 47076 37565 47104
rect 35676 47064 35682 47076
rect 37553 47073 37565 47076
rect 37599 47073 37611 47107
rect 37553 47067 37611 47073
rect 33229 47039 33287 47045
rect 33229 47036 33241 47039
rect 32232 47008 33241 47036
rect 32125 46999 32183 47005
rect 33229 47005 33241 47008
rect 33275 47005 33287 47039
rect 33229 46999 33287 47005
rect 34514 46996 34520 47048
rect 34572 47036 34578 47048
rect 35161 47039 35219 47045
rect 35161 47036 35173 47039
rect 34572 47008 35173 47036
rect 34572 46996 34578 47008
rect 35161 47005 35173 47008
rect 35207 47005 35219 47039
rect 35161 46999 35219 47005
rect 36078 46996 36084 47048
rect 36136 47036 36142 47048
rect 36449 47039 36507 47045
rect 36449 47036 36461 47039
rect 36136 47008 36461 47036
rect 36136 46996 36142 47008
rect 36449 47005 36461 47008
rect 36495 47005 36507 47039
rect 36449 46999 36507 47005
rect 37277 47039 37335 47045
rect 37277 47005 37289 47039
rect 37323 47005 37335 47039
rect 37277 46999 37335 47005
rect 27488 46940 30420 46968
rect 27488 46928 27494 46940
rect 37292 46912 37320 46999
rect 3896 46872 4200 46900
rect 12161 46903 12219 46909
rect 12161 46869 12173 46903
rect 12207 46869 12219 46903
rect 12161 46863 12219 46869
rect 12805 46903 12863 46909
rect 12805 46869 12817 46903
rect 12851 46869 12863 46903
rect 12805 46863 12863 46869
rect 16114 46860 16120 46912
rect 16172 46900 16178 46912
rect 16666 46900 16672 46912
rect 16172 46872 16672 46900
rect 16172 46860 16178 46872
rect 16666 46860 16672 46872
rect 16724 46860 16730 46912
rect 29546 46900 29552 46912
rect 29507 46872 29552 46900
rect 29546 46860 29552 46872
rect 29604 46860 29610 46912
rect 36354 46860 36360 46912
rect 36412 46900 36418 46912
rect 37274 46900 37280 46912
rect 36412 46872 37280 46900
rect 36412 46860 36418 46872
rect 37274 46860 37280 46872
rect 37332 46860 37338 46912
rect 37642 46860 37648 46912
rect 37700 46900 37706 46912
rect 39298 46900 39304 46912
rect 37700 46872 39304 46900
rect 37700 46860 37706 46872
rect 39298 46860 39304 46872
rect 39356 46860 39362 46912
rect 1104 46810 38824 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 38824 46810
rect 1104 46736 38824 46758
rect 658 46656 664 46708
rect 716 46696 722 46708
rect 3697 46699 3755 46705
rect 3697 46696 3709 46699
rect 716 46668 3709 46696
rect 716 46656 722 46668
rect 3697 46665 3709 46668
rect 3743 46665 3755 46699
rect 3697 46659 3755 46665
rect 3878 46656 3884 46708
rect 3936 46656 3942 46708
rect 5169 46699 5227 46705
rect 5169 46665 5181 46699
rect 5215 46696 5227 46699
rect 5350 46696 5356 46708
rect 5215 46668 5356 46696
rect 5215 46665 5227 46668
rect 5169 46659 5227 46665
rect 5350 46656 5356 46668
rect 5408 46656 5414 46708
rect 5810 46696 5816 46708
rect 5771 46668 5816 46696
rect 5810 46656 5816 46668
rect 5868 46656 5874 46708
rect 7101 46699 7159 46705
rect 7101 46665 7113 46699
rect 7147 46696 7159 46699
rect 7190 46696 7196 46708
rect 7147 46668 7196 46696
rect 7147 46665 7159 46668
rect 7101 46659 7159 46665
rect 7190 46656 7196 46668
rect 7248 46656 7254 46708
rect 7926 46696 7932 46708
rect 7887 46668 7932 46696
rect 7926 46656 7932 46668
rect 7984 46656 7990 46708
rect 10778 46656 10784 46708
rect 10836 46696 10842 46708
rect 10873 46699 10931 46705
rect 10873 46696 10885 46699
rect 10836 46668 10885 46696
rect 10836 46656 10842 46668
rect 10873 46665 10885 46668
rect 10919 46665 10931 46699
rect 13814 46696 13820 46708
rect 13775 46668 13820 46696
rect 10873 46659 10931 46665
rect 13814 46656 13820 46668
rect 13872 46656 13878 46708
rect 15470 46656 15476 46708
rect 15528 46696 15534 46708
rect 15841 46699 15899 46705
rect 15841 46696 15853 46699
rect 15528 46668 15853 46696
rect 15528 46656 15534 46668
rect 15841 46665 15853 46668
rect 15887 46665 15899 46699
rect 17402 46696 17408 46708
rect 17363 46668 17408 46696
rect 15841 46659 15899 46665
rect 17402 46656 17408 46668
rect 17460 46656 17466 46708
rect 19981 46699 20039 46705
rect 19981 46665 19993 46699
rect 20027 46696 20039 46699
rect 20254 46696 20260 46708
rect 20027 46668 20260 46696
rect 20027 46665 20039 46668
rect 19981 46659 20039 46665
rect 20254 46656 20260 46668
rect 20312 46656 20318 46708
rect 21266 46696 21272 46708
rect 21227 46668 21272 46696
rect 21266 46656 21272 46668
rect 21324 46656 21330 46708
rect 23014 46656 23020 46708
rect 23072 46696 23078 46708
rect 23937 46699 23995 46705
rect 23937 46696 23949 46699
rect 23072 46668 23949 46696
rect 23072 46656 23078 46668
rect 23937 46665 23949 46668
rect 23983 46665 23995 46699
rect 23937 46659 23995 46665
rect 25869 46699 25927 46705
rect 25869 46665 25881 46699
rect 25915 46696 25927 46699
rect 26050 46696 26056 46708
rect 25915 46668 26056 46696
rect 25915 46665 25927 46668
rect 25869 46659 25927 46665
rect 26050 46656 26056 46668
rect 26108 46656 26114 46708
rect 35161 46699 35219 46705
rect 35161 46665 35173 46699
rect 35207 46696 35219 46699
rect 35434 46696 35440 46708
rect 35207 46668 35440 46696
rect 35207 46665 35219 46668
rect 35161 46659 35219 46665
rect 35434 46656 35440 46668
rect 35492 46656 35498 46708
rect 36633 46699 36691 46705
rect 36633 46665 36645 46699
rect 36679 46696 36691 46699
rect 37366 46696 37372 46708
rect 36679 46668 37372 46696
rect 36679 46665 36691 46668
rect 36633 46659 36691 46665
rect 37366 46656 37372 46668
rect 37424 46656 37430 46708
rect 37458 46656 37464 46708
rect 37516 46656 37522 46708
rect 2961 46631 3019 46637
rect 2961 46597 2973 46631
rect 3007 46628 3019 46631
rect 3050 46628 3056 46640
rect 3007 46600 3056 46628
rect 3007 46597 3019 46600
rect 2961 46591 3019 46597
rect 3050 46588 3056 46600
rect 3108 46588 3114 46640
rect 3896 46628 3924 46656
rect 3896 46600 4384 46628
rect 2225 46563 2283 46569
rect 2225 46529 2237 46563
rect 2271 46560 2283 46563
rect 3142 46560 3148 46572
rect 2271 46532 3148 46560
rect 2271 46529 2283 46532
rect 2225 46523 2283 46529
rect 3142 46520 3148 46532
rect 3200 46520 3206 46572
rect 4356 46569 4384 46600
rect 3881 46563 3939 46569
rect 3881 46529 3893 46563
rect 3927 46529 3939 46563
rect 3881 46523 3939 46529
rect 4341 46563 4399 46569
rect 4341 46529 4353 46563
rect 4387 46529 4399 46563
rect 5828 46560 5856 46656
rect 14366 46588 14372 46640
rect 14424 46628 14430 46640
rect 15013 46631 15071 46637
rect 15013 46628 15025 46631
rect 14424 46600 15025 46628
rect 14424 46588 14430 46600
rect 15013 46597 15025 46600
rect 15059 46597 15071 46631
rect 15013 46591 15071 46597
rect 6365 46563 6423 46569
rect 6365 46560 6377 46563
rect 5828 46532 6377 46560
rect 4341 46523 4399 46529
rect 6365 46529 6377 46532
rect 6411 46529 6423 46563
rect 6365 46523 6423 46529
rect 8113 46563 8171 46569
rect 8113 46529 8125 46563
rect 8159 46560 8171 46563
rect 8294 46560 8300 46572
rect 8159 46532 8300 46560
rect 8159 46529 8171 46532
rect 8113 46523 8171 46529
rect 3896 46492 3924 46523
rect 8294 46520 8300 46532
rect 8352 46520 8358 46572
rect 8665 46563 8723 46569
rect 8665 46529 8677 46563
rect 8711 46560 8723 46563
rect 9122 46560 9128 46572
rect 8711 46532 9128 46560
rect 8711 46529 8723 46532
rect 8665 46523 8723 46529
rect 9122 46520 9128 46532
rect 9180 46520 9186 46572
rect 11698 46560 11704 46572
rect 11659 46532 11704 46560
rect 11698 46520 11704 46532
rect 11756 46520 11762 46572
rect 13722 46560 13728 46572
rect 13683 46532 13728 46560
rect 13722 46520 13728 46532
rect 13780 46520 13786 46572
rect 14921 46563 14979 46569
rect 14921 46529 14933 46563
rect 14967 46560 14979 46563
rect 16025 46563 16083 46569
rect 14967 46532 15792 46560
rect 14967 46529 14979 46532
rect 14921 46523 14979 46529
rect 8386 46492 8392 46504
rect 3896 46464 8392 46492
rect 8386 46452 8392 46464
rect 8444 46452 8450 46504
rect 12897 46495 12955 46501
rect 12897 46461 12909 46495
rect 12943 46492 12955 46495
rect 14001 46495 14059 46501
rect 14001 46492 14013 46495
rect 12943 46464 14013 46492
rect 12943 46461 12955 46464
rect 12897 46455 12955 46461
rect 14001 46461 14013 46464
rect 14047 46492 14059 46495
rect 15197 46495 15255 46501
rect 15197 46492 15209 46495
rect 14047 46464 15209 46492
rect 14047 46461 14059 46464
rect 14001 46455 14059 46461
rect 15197 46461 15209 46464
rect 15243 46492 15255 46495
rect 15286 46492 15292 46504
rect 15243 46464 15292 46492
rect 15243 46461 15255 46464
rect 15197 46455 15255 46461
rect 15286 46452 15292 46464
rect 15344 46452 15350 46504
rect 2409 46427 2467 46433
rect 2409 46393 2421 46427
rect 2455 46424 2467 46427
rect 2498 46424 2504 46436
rect 2455 46396 2504 46424
rect 2455 46393 2467 46396
rect 2409 46387 2467 46393
rect 2498 46384 2504 46396
rect 2556 46384 2562 46436
rect 9309 46427 9367 46433
rect 9309 46393 9321 46427
rect 9355 46424 9367 46427
rect 15764 46424 15792 46532
rect 16025 46529 16037 46563
rect 16071 46560 16083 46563
rect 16206 46560 16212 46572
rect 16071 46532 16212 46560
rect 16071 46529 16083 46532
rect 16025 46523 16083 46529
rect 16206 46520 16212 46532
rect 16264 46520 16270 46572
rect 17497 46563 17555 46569
rect 17497 46529 17509 46563
rect 17543 46529 17555 46563
rect 18782 46560 18788 46572
rect 18743 46532 18788 46560
rect 17497 46523 17555 46529
rect 16482 46452 16488 46504
rect 16540 46492 16546 46504
rect 17221 46495 17279 46501
rect 17221 46492 17233 46495
rect 16540 46464 17233 46492
rect 16540 46452 16546 46464
rect 17221 46461 17233 46464
rect 17267 46461 17279 46495
rect 17512 46492 17540 46523
rect 18782 46520 18788 46532
rect 18840 46520 18846 46572
rect 21284 46560 21312 46656
rect 32214 46588 32220 46640
rect 32272 46628 32278 46640
rect 32677 46631 32735 46637
rect 32677 46628 32689 46631
rect 32272 46600 32689 46628
rect 32272 46588 32278 46600
rect 32677 46597 32689 46600
rect 32723 46597 32735 46631
rect 32677 46591 32735 46597
rect 21821 46563 21879 46569
rect 21821 46560 21833 46563
rect 21284 46532 21833 46560
rect 21821 46529 21833 46532
rect 21867 46529 21879 46563
rect 21821 46523 21879 46529
rect 21910 46520 21916 46572
rect 21968 46560 21974 46572
rect 22649 46563 22707 46569
rect 22649 46560 22661 46563
rect 21968 46532 22661 46560
rect 21968 46520 21974 46532
rect 22649 46529 22661 46532
rect 22695 46560 22707 46563
rect 23109 46563 23167 46569
rect 23109 46560 23121 46563
rect 22695 46532 23121 46560
rect 22695 46529 22707 46532
rect 22649 46523 22707 46529
rect 23109 46529 23121 46532
rect 23155 46529 23167 46563
rect 24762 46560 24768 46572
rect 24723 46532 24768 46560
rect 23109 46523 23167 46529
rect 24762 46520 24768 46532
rect 24820 46560 24826 46572
rect 25225 46563 25283 46569
rect 25225 46560 25237 46563
rect 24820 46532 25237 46560
rect 24820 46520 24826 46532
rect 25225 46529 25237 46532
rect 25271 46529 25283 46563
rect 28626 46560 28632 46572
rect 28587 46532 28632 46560
rect 25225 46523 25283 46529
rect 28626 46520 28632 46532
rect 28684 46560 28690 46572
rect 29089 46563 29147 46569
rect 29089 46560 29101 46563
rect 28684 46532 29101 46560
rect 28684 46520 28690 46532
rect 29089 46529 29101 46532
rect 29135 46529 29147 46563
rect 29914 46560 29920 46572
rect 29875 46532 29920 46560
rect 29089 46523 29147 46529
rect 29914 46520 29920 46532
rect 29972 46560 29978 46572
rect 30377 46563 30435 46569
rect 30377 46560 30389 46563
rect 29972 46532 30389 46560
rect 29972 46520 29978 46532
rect 30377 46529 30389 46532
rect 30423 46529 30435 46563
rect 33778 46560 33784 46572
rect 33739 46532 33784 46560
rect 30377 46523 30435 46529
rect 33778 46520 33784 46532
rect 33836 46520 33842 46572
rect 34422 46560 34428 46572
rect 34383 46532 34428 46560
rect 34422 46520 34428 46532
rect 34480 46520 34486 46572
rect 34790 46520 34796 46572
rect 34848 46560 34854 46572
rect 34977 46563 35035 46569
rect 34977 46560 34989 46563
rect 34848 46532 34989 46560
rect 34848 46520 34854 46532
rect 34977 46529 34989 46532
rect 35023 46529 35035 46563
rect 34977 46523 35035 46529
rect 35894 46520 35900 46572
rect 35952 46560 35958 46572
rect 35952 46532 35997 46560
rect 35952 46520 35958 46532
rect 36262 46520 36268 46572
rect 36320 46560 36326 46572
rect 36449 46563 36507 46569
rect 36449 46560 36461 46563
rect 36320 46532 36461 46560
rect 36320 46520 36326 46532
rect 36449 46529 36461 46532
rect 36495 46529 36507 46563
rect 36449 46523 36507 46529
rect 37277 46563 37335 46569
rect 37277 46529 37289 46563
rect 37323 46560 37335 46563
rect 37476 46560 37504 46656
rect 37323 46532 37504 46560
rect 37323 46529 37335 46532
rect 37277 46523 37335 46529
rect 29546 46492 29552 46504
rect 17512 46464 29552 46492
rect 17221 46455 17279 46461
rect 29546 46452 29552 46464
rect 29604 46452 29610 46504
rect 35526 46452 35532 46504
rect 35584 46492 35590 46504
rect 37292 46492 37320 46523
rect 35584 46464 37320 46492
rect 35584 46452 35590 46464
rect 37458 46452 37464 46504
rect 37516 46492 37522 46504
rect 37553 46495 37611 46501
rect 37553 46492 37565 46495
rect 37516 46464 37565 46492
rect 37516 46452 37522 46464
rect 37553 46461 37565 46464
rect 37599 46461 37611 46495
rect 37553 46455 37611 46461
rect 24581 46427 24639 46433
rect 24581 46424 24593 46427
rect 9355 46396 14872 46424
rect 15764 46396 24593 46424
rect 9355 46393 9367 46396
rect 9309 46387 9367 46393
rect 1673 46359 1731 46365
rect 1673 46325 1685 46359
rect 1719 46356 1731 46359
rect 2314 46356 2320 46368
rect 1719 46328 2320 46356
rect 1719 46325 1731 46328
rect 1673 46319 1731 46325
rect 2314 46316 2320 46328
rect 2372 46316 2378 46368
rect 3050 46356 3056 46368
rect 3011 46328 3056 46356
rect 3050 46316 3056 46328
rect 3108 46316 3114 46368
rect 4525 46359 4583 46365
rect 4525 46325 4537 46359
rect 4571 46356 4583 46359
rect 5350 46356 5356 46368
rect 4571 46328 5356 46356
rect 4571 46325 4583 46328
rect 4525 46319 4583 46325
rect 5350 46316 5356 46328
rect 5408 46316 5414 46368
rect 6546 46356 6552 46368
rect 6507 46328 6552 46356
rect 6546 46316 6552 46328
rect 6604 46316 6610 46368
rect 10042 46316 10048 46368
rect 10100 46356 10106 46368
rect 10229 46359 10287 46365
rect 10229 46356 10241 46359
rect 10100 46328 10241 46356
rect 10100 46316 10106 46328
rect 10229 46325 10241 46328
rect 10275 46356 10287 46359
rect 10686 46356 10692 46368
rect 10275 46328 10692 46356
rect 10275 46325 10287 46328
rect 10229 46319 10287 46325
rect 10686 46316 10692 46328
rect 10744 46316 10750 46368
rect 11885 46359 11943 46365
rect 11885 46325 11897 46359
rect 11931 46356 11943 46359
rect 12710 46356 12716 46368
rect 11931 46328 12716 46356
rect 11931 46325 11943 46328
rect 11885 46319 11943 46325
rect 12710 46316 12716 46328
rect 12768 46316 12774 46368
rect 13357 46359 13415 46365
rect 13357 46325 13369 46359
rect 13403 46356 13415 46359
rect 13446 46356 13452 46368
rect 13403 46328 13452 46356
rect 13403 46325 13415 46328
rect 13357 46319 13415 46325
rect 13446 46316 13452 46328
rect 13504 46316 13510 46368
rect 14274 46316 14280 46368
rect 14332 46356 14338 46368
rect 14553 46359 14611 46365
rect 14553 46356 14565 46359
rect 14332 46328 14565 46356
rect 14332 46316 14338 46328
rect 14553 46325 14565 46328
rect 14599 46325 14611 46359
rect 14844 46356 14872 46396
rect 24581 46393 24593 46396
rect 24627 46393 24639 46427
rect 24581 46387 24639 46393
rect 27154 46384 27160 46436
rect 27212 46424 27218 46436
rect 29733 46427 29791 46433
rect 29733 46424 29745 46427
rect 27212 46396 29745 46424
rect 27212 46384 27218 46396
rect 29733 46393 29745 46396
rect 29779 46393 29791 46427
rect 29733 46387 29791 46393
rect 31570 46384 31576 46436
rect 31628 46424 31634 46436
rect 34241 46427 34299 46433
rect 34241 46424 34253 46427
rect 31628 46396 34253 46424
rect 31628 46384 31634 46396
rect 34241 46393 34253 46396
rect 34287 46393 34299 46427
rect 34241 46387 34299 46393
rect 35434 46384 35440 46436
rect 35492 46424 35498 46436
rect 35713 46427 35771 46433
rect 35713 46424 35725 46427
rect 35492 46396 35725 46424
rect 35492 46384 35498 46396
rect 35713 46393 35725 46396
rect 35759 46393 35771 46427
rect 35713 46387 35771 46393
rect 15194 46356 15200 46368
rect 14844 46328 15200 46356
rect 14553 46319 14611 46325
rect 15194 46316 15200 46328
rect 15252 46316 15258 46368
rect 17770 46316 17776 46368
rect 17828 46356 17834 46368
rect 17865 46359 17923 46365
rect 17865 46356 17877 46359
rect 17828 46328 17877 46356
rect 17828 46316 17834 46328
rect 17865 46325 17877 46328
rect 17911 46325 17923 46359
rect 18966 46356 18972 46368
rect 18927 46328 18972 46356
rect 17865 46319 17923 46325
rect 18966 46316 18972 46328
rect 19024 46316 19030 46368
rect 22005 46359 22063 46365
rect 22005 46325 22017 46359
rect 22051 46356 22063 46359
rect 22094 46356 22100 46368
rect 22051 46328 22100 46356
rect 22051 46325 22063 46328
rect 22005 46319 22063 46325
rect 22094 46316 22100 46328
rect 22152 46316 22158 46368
rect 22186 46316 22192 46368
rect 22244 46356 22250 46368
rect 22465 46359 22523 46365
rect 22465 46356 22477 46359
rect 22244 46328 22477 46356
rect 22244 46316 22250 46328
rect 22465 46325 22477 46328
rect 22511 46325 22523 46359
rect 27890 46356 27896 46368
rect 27851 46328 27896 46356
rect 22465 46319 22523 46325
rect 27890 46316 27896 46328
rect 27948 46316 27954 46368
rect 28442 46356 28448 46368
rect 28403 46328 28448 46356
rect 28442 46316 28448 46328
rect 28500 46316 28506 46368
rect 30926 46356 30932 46368
rect 30887 46328 30932 46356
rect 30926 46316 30932 46328
rect 30984 46316 30990 46368
rect 31478 46356 31484 46368
rect 31439 46328 31484 46356
rect 31478 46316 31484 46328
rect 31536 46316 31542 46368
rect 32582 46356 32588 46368
rect 32543 46328 32588 46356
rect 32582 46316 32588 46328
rect 32640 46316 32646 46368
rect 33594 46356 33600 46368
rect 33555 46328 33600 46356
rect 33594 46316 33600 46328
rect 33652 46316 33658 46368
rect 1104 46266 38824 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 38824 46266
rect 1104 46192 38824 46214
rect 2225 46155 2283 46161
rect 2225 46121 2237 46155
rect 2271 46152 2283 46155
rect 2774 46152 2780 46164
rect 2271 46124 2780 46152
rect 2271 46121 2283 46124
rect 2225 46115 2283 46121
rect 2774 46112 2780 46124
rect 2832 46112 2838 46164
rect 2958 46152 2964 46164
rect 2919 46124 2964 46152
rect 2958 46112 2964 46124
rect 3016 46112 3022 46164
rect 3878 46112 3884 46164
rect 3936 46152 3942 46164
rect 4157 46155 4215 46161
rect 4157 46152 4169 46155
rect 3936 46124 4169 46152
rect 3936 46112 3942 46124
rect 4157 46121 4169 46124
rect 4203 46121 4215 46155
rect 4157 46115 4215 46121
rect 4798 46112 4804 46164
rect 4856 46152 4862 46164
rect 4893 46155 4951 46161
rect 4893 46152 4905 46155
rect 4856 46124 4905 46152
rect 4856 46112 4862 46124
rect 4893 46121 4905 46124
rect 4939 46152 4951 46155
rect 5074 46152 5080 46164
rect 4939 46124 5080 46152
rect 4939 46121 4951 46124
rect 4893 46115 4951 46121
rect 5074 46112 5080 46124
rect 5132 46112 5138 46164
rect 6457 46155 6515 46161
rect 6457 46121 6469 46155
rect 6503 46152 6515 46155
rect 6638 46152 6644 46164
rect 6503 46124 6644 46152
rect 6503 46121 6515 46124
rect 6457 46115 6515 46121
rect 6638 46112 6644 46124
rect 6696 46112 6702 46164
rect 8938 46152 8944 46164
rect 8899 46124 8944 46152
rect 8938 46112 8944 46124
rect 8996 46112 9002 46164
rect 11609 46155 11667 46161
rect 11609 46121 11621 46155
rect 11655 46152 11667 46155
rect 11698 46152 11704 46164
rect 11655 46124 11704 46152
rect 11655 46121 11667 46124
rect 11609 46115 11667 46121
rect 11698 46112 11704 46124
rect 11756 46112 11762 46164
rect 11974 46112 11980 46164
rect 12032 46152 12038 46164
rect 12161 46155 12219 46161
rect 12161 46152 12173 46155
rect 12032 46124 12173 46152
rect 12032 46112 12038 46124
rect 12161 46121 12173 46124
rect 12207 46121 12219 46155
rect 12161 46115 12219 46121
rect 12710 46112 12716 46164
rect 12768 46152 12774 46164
rect 15102 46152 15108 46164
rect 12768 46124 14596 46152
rect 15063 46124 15108 46152
rect 12768 46112 12774 46124
rect 3234 46044 3240 46096
rect 3292 46084 3298 46096
rect 5537 46087 5595 46093
rect 5537 46084 5549 46087
rect 3292 46056 5549 46084
rect 3292 46044 3298 46056
rect 5537 46053 5549 46056
rect 5583 46053 5595 46087
rect 13265 46087 13323 46093
rect 13265 46084 13277 46087
rect 5537 46047 5595 46053
rect 6886 46056 13277 46084
rect 6886 46016 6914 46056
rect 13265 46053 13277 46056
rect 13311 46053 13323 46087
rect 13265 46047 13323 46053
rect 14461 46087 14519 46093
rect 14461 46053 14473 46087
rect 14507 46053 14519 46087
rect 14568 46084 14596 46124
rect 15102 46112 15108 46124
rect 15160 46112 15166 46164
rect 15194 46112 15200 46164
rect 15252 46152 15258 46164
rect 17126 46152 17132 46164
rect 15252 46124 17132 46152
rect 15252 46112 15258 46124
rect 17126 46112 17132 46124
rect 17184 46112 17190 46164
rect 19334 46152 19340 46164
rect 19295 46124 19340 46152
rect 19334 46112 19340 46124
rect 19392 46112 19398 46164
rect 24394 46152 24400 46164
rect 24355 46124 24400 46152
rect 24394 46112 24400 46124
rect 24452 46112 24458 46164
rect 29638 46152 29644 46164
rect 29599 46124 29644 46152
rect 29638 46112 29644 46124
rect 29696 46112 29702 46164
rect 32214 46112 32220 46164
rect 32272 46152 32278 46164
rect 32309 46155 32367 46161
rect 32309 46152 32321 46155
rect 32272 46124 32321 46152
rect 32272 46112 32278 46124
rect 32309 46121 32321 46124
rect 32355 46121 32367 46155
rect 32950 46152 32956 46164
rect 32911 46124 32956 46152
rect 32309 46115 32367 46121
rect 32950 46112 32956 46124
rect 33008 46112 33014 46164
rect 33505 46155 33563 46161
rect 33505 46121 33517 46155
rect 33551 46152 33563 46155
rect 33778 46152 33784 46164
rect 33551 46124 33784 46152
rect 33551 46121 33563 46124
rect 33505 46115 33563 46121
rect 33778 46112 33784 46124
rect 33836 46112 33842 46164
rect 34149 46155 34207 46161
rect 34149 46121 34161 46155
rect 34195 46152 34207 46155
rect 34422 46152 34428 46164
rect 34195 46124 34428 46152
rect 34195 46121 34207 46124
rect 34149 46115 34207 46121
rect 34422 46112 34428 46124
rect 34480 46112 34486 46164
rect 35802 46112 35808 46164
rect 35860 46152 35866 46164
rect 36725 46155 36783 46161
rect 36725 46152 36737 46155
rect 35860 46124 36737 46152
rect 35860 46112 35866 46124
rect 36725 46121 36737 46124
rect 36771 46121 36783 46155
rect 36725 46115 36783 46121
rect 20806 46084 20812 46096
rect 14568 46056 20812 46084
rect 14461 46047 14519 46053
rect 1688 45988 6914 46016
rect 1688 45957 1716 45988
rect 1673 45951 1731 45957
rect 1673 45917 1685 45951
rect 1719 45917 1731 45951
rect 1673 45911 1731 45917
rect 2314 45908 2320 45960
rect 2372 45948 2378 45960
rect 2409 45951 2467 45957
rect 2409 45948 2421 45951
rect 2372 45920 2421 45948
rect 2372 45908 2378 45920
rect 2409 45917 2421 45920
rect 2455 45948 2467 45951
rect 2682 45948 2688 45960
rect 2455 45920 2688 45948
rect 2455 45917 2467 45920
rect 2409 45911 2467 45917
rect 2682 45908 2688 45920
rect 2740 45908 2746 45960
rect 3145 45951 3203 45957
rect 3145 45917 3157 45951
rect 3191 45948 3203 45951
rect 3234 45948 3240 45960
rect 3191 45920 3240 45948
rect 3191 45917 3203 45920
rect 3145 45911 3203 45917
rect 3234 45908 3240 45920
rect 3292 45908 3298 45960
rect 12805 45951 12863 45957
rect 12805 45917 12817 45951
rect 12851 45948 12863 45951
rect 13262 45948 13268 45960
rect 12851 45920 13268 45948
rect 12851 45917 12863 45920
rect 12805 45911 12863 45917
rect 13262 45908 13268 45920
rect 13320 45908 13326 45960
rect 13446 45948 13452 45960
rect 13407 45920 13452 45948
rect 13446 45908 13452 45920
rect 13504 45908 13510 45960
rect 14274 45948 14280 45960
rect 14235 45920 14280 45948
rect 14274 45908 14280 45920
rect 14332 45908 14338 45960
rect 14476 45948 14504 46047
rect 20806 46044 20812 46056
rect 20864 46044 20870 46096
rect 23474 46044 23480 46096
rect 23532 46084 23538 46096
rect 33594 46084 33600 46096
rect 23532 46056 33600 46084
rect 23532 46044 23538 46056
rect 33594 46044 33600 46056
rect 33652 46044 33658 46096
rect 35710 46044 35716 46096
rect 35768 46084 35774 46096
rect 35989 46087 36047 46093
rect 35989 46084 36001 46087
rect 35768 46056 36001 46084
rect 35768 46044 35774 46056
rect 35989 46053 36001 46056
rect 36035 46053 36047 46087
rect 35989 46047 36047 46053
rect 16022 45976 16028 46028
rect 16080 46016 16086 46028
rect 16482 46016 16488 46028
rect 16080 45988 16488 46016
rect 16080 45976 16086 45988
rect 16482 45976 16488 45988
rect 16540 46016 16546 46028
rect 16669 46019 16727 46025
rect 16669 46016 16681 46019
rect 16540 45988 16681 46016
rect 16540 45976 16546 45988
rect 16669 45985 16681 45988
rect 16715 45985 16727 46019
rect 16669 45979 16727 45985
rect 16853 46019 16911 46025
rect 16853 45985 16865 46019
rect 16899 46016 16911 46019
rect 18046 46016 18052 46028
rect 16899 45988 18052 46016
rect 16899 45985 16911 45988
rect 16853 45979 16911 45985
rect 18046 45976 18052 45988
rect 18104 45976 18110 46028
rect 35250 45976 35256 46028
rect 35308 46016 35314 46028
rect 35526 46016 35532 46028
rect 35308 45988 35532 46016
rect 35308 45976 35314 45988
rect 35526 45976 35532 45988
rect 35584 45976 35590 46028
rect 37277 46019 37335 46025
rect 37277 45985 37289 46019
rect 37323 46016 37335 46019
rect 37642 46016 37648 46028
rect 37323 45988 37648 46016
rect 37323 45985 37335 45988
rect 37277 45979 37335 45985
rect 37642 45976 37648 45988
rect 37700 45976 37706 46028
rect 14921 45951 14979 45957
rect 14921 45948 14933 45951
rect 14476 45920 14933 45948
rect 14921 45917 14933 45920
rect 14967 45917 14979 45951
rect 14921 45911 14979 45917
rect 15378 45908 15384 45960
rect 15436 45948 15442 45960
rect 16945 45951 17003 45957
rect 16945 45948 16957 45951
rect 15436 45920 16957 45948
rect 15436 45908 15442 45920
rect 16945 45917 16957 45920
rect 16991 45917 17003 45951
rect 18322 45948 18328 45960
rect 18283 45920 18328 45948
rect 16945 45911 17003 45917
rect 18322 45908 18328 45920
rect 18380 45908 18386 45960
rect 35342 45948 35348 45960
rect 35303 45920 35348 45948
rect 35342 45908 35348 45920
rect 35400 45908 35406 45960
rect 35805 45951 35863 45957
rect 35805 45917 35817 45951
rect 35851 45917 35863 45951
rect 35805 45911 35863 45917
rect 8294 45880 8300 45892
rect 8207 45852 8300 45880
rect 8294 45840 8300 45852
rect 8352 45880 8358 45892
rect 9030 45880 9036 45892
rect 8352 45852 9036 45880
rect 8352 45840 8358 45852
rect 9030 45840 9036 45852
rect 9088 45840 9094 45892
rect 34606 45840 34612 45892
rect 34664 45880 34670 45892
rect 35820 45880 35848 45911
rect 35986 45908 35992 45960
rect 36044 45948 36050 45960
rect 36541 45951 36599 45957
rect 36541 45948 36553 45951
rect 36044 45920 36553 45948
rect 36044 45908 36050 45920
rect 36541 45917 36553 45920
rect 36587 45917 36599 45951
rect 37550 45948 37556 45960
rect 37511 45920 37556 45948
rect 36541 45911 36599 45917
rect 37550 45908 37556 45920
rect 37608 45908 37614 45960
rect 34664 45852 35848 45880
rect 34664 45840 34670 45852
rect 1486 45812 1492 45824
rect 1447 45784 1492 45812
rect 1486 45772 1492 45784
rect 1544 45772 1550 45824
rect 2958 45772 2964 45824
rect 3016 45812 3022 45824
rect 3142 45812 3148 45824
rect 3016 45784 3148 45812
rect 3016 45772 3022 45784
rect 3142 45772 3148 45784
rect 3200 45772 3206 45824
rect 16022 45812 16028 45824
rect 15983 45784 16028 45812
rect 16022 45772 16028 45784
rect 16080 45772 16086 45824
rect 17310 45812 17316 45824
rect 17271 45784 17316 45812
rect 17310 45772 17316 45784
rect 17368 45772 17374 45824
rect 17862 45772 17868 45824
rect 17920 45812 17926 45824
rect 18141 45815 18199 45821
rect 18141 45812 18153 45815
rect 17920 45784 18153 45812
rect 17920 45772 17926 45784
rect 18141 45781 18153 45784
rect 18187 45781 18199 45815
rect 18141 45775 18199 45781
rect 35161 45815 35219 45821
rect 35161 45781 35173 45815
rect 35207 45812 35219 45815
rect 35618 45812 35624 45824
rect 35207 45784 35624 45812
rect 35207 45781 35219 45784
rect 35161 45775 35219 45781
rect 35618 45772 35624 45784
rect 35676 45772 35682 45824
rect 1104 45722 38824 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 38824 45722
rect 1104 45648 38824 45670
rect 18693 45611 18751 45617
rect 18693 45577 18705 45611
rect 18739 45608 18751 45611
rect 18782 45608 18788 45620
rect 18739 45580 18788 45608
rect 18739 45577 18751 45580
rect 18693 45571 18751 45577
rect 18782 45568 18788 45580
rect 18840 45568 18846 45620
rect 35342 45568 35348 45620
rect 35400 45608 35406 45620
rect 35437 45611 35495 45617
rect 35437 45608 35449 45611
rect 35400 45580 35449 45608
rect 35400 45568 35406 45580
rect 35437 45577 35449 45580
rect 35483 45577 35495 45611
rect 35437 45571 35495 45577
rect 14 45500 20 45552
rect 72 45540 78 45552
rect 72 45512 2544 45540
rect 72 45500 78 45512
rect 106 45432 112 45484
rect 164 45472 170 45484
rect 1302 45472 1308 45484
rect 164 45444 1308 45472
rect 164 45432 170 45444
rect 1302 45432 1308 45444
rect 1360 45472 1366 45484
rect 2516 45481 2544 45512
rect 2958 45500 2964 45552
rect 3016 45540 3022 45552
rect 4341 45543 4399 45549
rect 4341 45540 4353 45543
rect 3016 45512 4353 45540
rect 3016 45500 3022 45512
rect 4341 45509 4353 45512
rect 4387 45509 4399 45543
rect 4341 45503 4399 45509
rect 12618 45500 12624 45552
rect 12676 45540 12682 45552
rect 12897 45543 12955 45549
rect 12897 45540 12909 45543
rect 12676 45512 12909 45540
rect 12676 45500 12682 45512
rect 12897 45509 12909 45512
rect 12943 45509 12955 45543
rect 13906 45540 13912 45552
rect 13867 45512 13912 45540
rect 12897 45503 12955 45509
rect 13906 45500 13912 45512
rect 13964 45500 13970 45552
rect 17129 45543 17187 45549
rect 17129 45509 17141 45543
rect 17175 45540 17187 45543
rect 17310 45540 17316 45552
rect 17175 45512 17316 45540
rect 17175 45509 17187 45512
rect 17129 45503 17187 45509
rect 17310 45500 17316 45512
rect 17368 45500 17374 45552
rect 34333 45543 34391 45549
rect 34333 45509 34345 45543
rect 34379 45540 34391 45543
rect 34698 45540 34704 45552
rect 34379 45512 34704 45540
rect 34379 45509 34391 45512
rect 34333 45503 34391 45509
rect 34698 45500 34704 45512
rect 34756 45500 34762 45552
rect 37366 45540 37372 45552
rect 36740 45512 37372 45540
rect 1857 45475 1915 45481
rect 1857 45472 1869 45475
rect 1360 45444 1869 45472
rect 1360 45432 1366 45444
rect 1857 45441 1869 45444
rect 1903 45441 1915 45475
rect 1857 45435 1915 45441
rect 2501 45475 2559 45481
rect 2501 45441 2513 45475
rect 2547 45441 2559 45475
rect 2501 45435 2559 45441
rect 2516 45404 2544 45435
rect 2590 45432 2596 45484
rect 2648 45472 2654 45484
rect 4893 45475 4951 45481
rect 4893 45472 4905 45475
rect 2648 45444 4905 45472
rect 2648 45432 2654 45444
rect 4893 45441 4905 45444
rect 4939 45441 4951 45475
rect 17770 45472 17776 45484
rect 17731 45444 17776 45472
rect 4893 45435 4951 45441
rect 17770 45432 17776 45444
rect 17828 45432 17834 45484
rect 33781 45475 33839 45481
rect 33781 45441 33793 45475
rect 33827 45472 33839 45475
rect 35250 45472 35256 45484
rect 33827 45444 35256 45472
rect 33827 45441 33839 45444
rect 33781 45435 33839 45441
rect 35250 45432 35256 45444
rect 35308 45432 35314 45484
rect 36740 45481 36768 45512
rect 37366 45500 37372 45512
rect 37424 45500 37430 45552
rect 36725 45475 36783 45481
rect 36725 45441 36737 45475
rect 36771 45441 36783 45475
rect 36725 45435 36783 45441
rect 36814 45432 36820 45484
rect 36872 45472 36878 45484
rect 37829 45475 37887 45481
rect 37829 45472 37841 45475
rect 36872 45444 37841 45472
rect 36872 45432 36878 45444
rect 37829 45441 37841 45444
rect 37875 45441 37887 45475
rect 37829 45435 37887 45441
rect 3789 45407 3847 45413
rect 3789 45404 3801 45407
rect 2516 45376 3801 45404
rect 3789 45373 3801 45376
rect 3835 45373 3847 45407
rect 3789 45367 3847 45373
rect 2041 45339 2099 45345
rect 2041 45305 2053 45339
rect 2087 45336 2099 45339
rect 2406 45336 2412 45348
rect 2087 45308 2412 45336
rect 2087 45305 2099 45308
rect 2041 45299 2099 45305
rect 2406 45296 2412 45308
rect 2464 45296 2470 45348
rect 2685 45339 2743 45345
rect 2685 45305 2697 45339
rect 2731 45336 2743 45339
rect 13722 45336 13728 45348
rect 2731 45308 13728 45336
rect 2731 45305 2743 45308
rect 2685 45299 2743 45305
rect 13722 45296 13728 45308
rect 13780 45296 13786 45348
rect 17313 45339 17371 45345
rect 17313 45305 17325 45339
rect 17359 45336 17371 45339
rect 17586 45336 17592 45348
rect 17359 45308 17592 45336
rect 17359 45305 17371 45308
rect 17313 45299 17371 45305
rect 17586 45296 17592 45308
rect 17644 45296 17650 45348
rect 17954 45336 17960 45348
rect 17915 45308 17960 45336
rect 17954 45296 17960 45308
rect 18012 45296 18018 45348
rect 22002 45296 22008 45348
rect 22060 45336 22066 45348
rect 35986 45336 35992 45348
rect 22060 45308 35992 45336
rect 22060 45296 22066 45308
rect 35986 45296 35992 45308
rect 36044 45296 36050 45348
rect 3234 45268 3240 45280
rect 3195 45240 3240 45268
rect 3234 45228 3240 45240
rect 3292 45228 3298 45280
rect 14366 45268 14372 45280
rect 14327 45240 14372 45268
rect 14366 45228 14372 45240
rect 14424 45228 14430 45280
rect 15194 45228 15200 45280
rect 15252 45268 15258 45280
rect 15381 45271 15439 45277
rect 15381 45268 15393 45271
rect 15252 45240 15393 45268
rect 15252 45228 15258 45240
rect 15381 45237 15393 45240
rect 15427 45268 15439 45271
rect 16022 45268 16028 45280
rect 15427 45240 16028 45268
rect 15427 45237 15439 45240
rect 15381 45231 15439 45237
rect 16022 45228 16028 45240
rect 16080 45228 16086 45280
rect 34790 45268 34796 45280
rect 34751 45240 34796 45268
rect 34790 45228 34796 45240
rect 34848 45228 34854 45280
rect 36538 45268 36544 45280
rect 36499 45240 36544 45268
rect 36538 45228 36544 45240
rect 36596 45228 36602 45280
rect 38010 45268 38016 45280
rect 37971 45240 38016 45268
rect 38010 45228 38016 45240
rect 38068 45228 38074 45280
rect 1104 45178 38824 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 38824 45178
rect 1104 45104 38824 45126
rect 3786 45064 3792 45076
rect 3747 45036 3792 45064
rect 3786 45024 3792 45036
rect 3844 45024 3850 45076
rect 16666 45064 16672 45076
rect 16627 45036 16672 45064
rect 16666 45024 16672 45036
rect 16724 45024 16730 45076
rect 18049 45067 18107 45073
rect 18049 45033 18061 45067
rect 18095 45064 18107 45067
rect 18322 45064 18328 45076
rect 18095 45036 18328 45064
rect 18095 45033 18107 45036
rect 18049 45027 18107 45033
rect 18322 45024 18328 45036
rect 18380 45024 18386 45076
rect 35894 45024 35900 45076
rect 35952 45064 35958 45076
rect 36081 45067 36139 45073
rect 36081 45064 36093 45067
rect 35952 45036 36093 45064
rect 35952 45024 35958 45036
rect 36081 45033 36093 45036
rect 36127 45033 36139 45067
rect 36081 45027 36139 45033
rect 30374 44956 30380 45008
rect 30432 44996 30438 45008
rect 37185 44999 37243 45005
rect 37185 44996 37197 44999
rect 30432 44968 37197 44996
rect 30432 44956 30438 44968
rect 37185 44965 37197 44968
rect 37231 44965 37243 44999
rect 37185 44959 37243 44965
rect 33594 44928 33600 44940
rect 33555 44900 33600 44928
rect 33594 44888 33600 44900
rect 33652 44888 33658 44940
rect 35621 44931 35679 44937
rect 35621 44897 35633 44931
rect 35667 44928 35679 44931
rect 38102 44928 38108 44940
rect 35667 44900 38108 44928
rect 35667 44897 35679 44900
rect 35621 44891 35679 44897
rect 2501 44863 2559 44869
rect 2501 44829 2513 44863
rect 2547 44860 2559 44863
rect 2774 44860 2780 44872
rect 2547 44832 2780 44860
rect 2547 44829 2559 44832
rect 2501 44823 2559 44829
rect 2774 44820 2780 44832
rect 2832 44860 2838 44872
rect 3145 44863 3203 44869
rect 3145 44860 3157 44863
rect 2832 44832 3157 44860
rect 2832 44820 2838 44832
rect 3145 44829 3157 44832
rect 3191 44829 3203 44863
rect 3145 44823 3203 44829
rect 33781 44863 33839 44869
rect 33781 44829 33793 44863
rect 33827 44860 33839 44863
rect 36538 44860 36544 44872
rect 33827 44832 36544 44860
rect 33827 44829 33839 44832
rect 33781 44823 33839 44829
rect 36538 44820 36544 44832
rect 36596 44820 36602 44872
rect 36725 44863 36783 44869
rect 36725 44829 36737 44863
rect 36771 44860 36783 44863
rect 37182 44860 37188 44872
rect 36771 44832 37188 44860
rect 36771 44829 36783 44832
rect 36725 44823 36783 44829
rect 37182 44820 37188 44832
rect 37240 44860 37246 44872
rect 38028 44869 38056 44900
rect 38102 44888 38108 44900
rect 38160 44888 38166 44940
rect 37369 44863 37427 44869
rect 37369 44860 37381 44863
rect 37240 44832 37381 44860
rect 37240 44820 37246 44832
rect 37369 44829 37381 44832
rect 37415 44829 37427 44863
rect 37369 44823 37427 44829
rect 38013 44863 38071 44869
rect 38013 44829 38025 44863
rect 38059 44829 38071 44863
rect 38013 44823 38071 44829
rect 1857 44795 1915 44801
rect 1857 44761 1869 44795
rect 1903 44792 1915 44795
rect 2866 44792 2872 44804
rect 1903 44764 2872 44792
rect 1903 44761 1915 44764
rect 1857 44755 1915 44761
rect 2866 44752 2872 44764
rect 2924 44752 2930 44804
rect 7466 44752 7472 44804
rect 7524 44792 7530 44804
rect 32861 44795 32919 44801
rect 32861 44792 32873 44795
rect 7524 44764 32873 44792
rect 7524 44752 7530 44764
rect 32861 44761 32873 44764
rect 32907 44792 32919 44795
rect 33689 44795 33747 44801
rect 33689 44792 33701 44795
rect 32907 44764 33701 44792
rect 32907 44761 32919 44764
rect 32861 44755 32919 44761
rect 33689 44761 33701 44764
rect 33735 44761 33747 44795
rect 33689 44755 33747 44761
rect 35069 44795 35127 44801
rect 35069 44761 35081 44795
rect 35115 44792 35127 44795
rect 37642 44792 37648 44804
rect 35115 44764 37648 44792
rect 35115 44761 35127 44764
rect 35069 44755 35127 44761
rect 37642 44752 37648 44764
rect 37700 44752 37706 44804
rect 1946 44724 1952 44736
rect 1907 44696 1952 44724
rect 1946 44684 1952 44696
rect 2004 44684 2010 44736
rect 2685 44727 2743 44733
rect 2685 44693 2697 44727
rect 2731 44724 2743 44727
rect 4614 44724 4620 44736
rect 2731 44696 4620 44724
rect 2731 44693 2743 44696
rect 2685 44687 2743 44693
rect 4614 44684 4620 44696
rect 4672 44684 4678 44736
rect 16206 44724 16212 44736
rect 16167 44696 16212 44724
rect 16206 44684 16212 44696
rect 16264 44684 16270 44736
rect 34149 44727 34207 44733
rect 34149 44693 34161 44727
rect 34195 44724 34207 44727
rect 34698 44724 34704 44736
rect 34195 44696 34704 44724
rect 34195 44693 34207 44696
rect 34149 44687 34207 44693
rect 34698 44684 34704 44696
rect 34756 44684 34762 44736
rect 37921 44727 37979 44733
rect 37921 44693 37933 44727
rect 37967 44724 37979 44727
rect 38194 44724 38200 44736
rect 37967 44696 38200 44724
rect 37967 44693 37979 44696
rect 37921 44687 37979 44693
rect 38194 44684 38200 44696
rect 38252 44684 38258 44736
rect 1104 44634 38824 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 38824 44634
rect 1104 44560 38824 44582
rect 2685 44523 2743 44529
rect 2685 44489 2697 44523
rect 2731 44520 2743 44523
rect 2866 44520 2872 44532
rect 2731 44492 2872 44520
rect 2731 44489 2743 44492
rect 2685 44483 2743 44489
rect 2866 44480 2872 44492
rect 2924 44480 2930 44532
rect 1302 44412 1308 44464
rect 1360 44452 1366 44464
rect 3145 44455 3203 44461
rect 3145 44452 3157 44455
rect 1360 44424 3157 44452
rect 1360 44412 1366 44424
rect 3145 44421 3157 44424
rect 3191 44421 3203 44455
rect 3145 44415 3203 44421
rect 1394 44384 1400 44396
rect 1355 44356 1400 44384
rect 1394 44344 1400 44356
rect 1452 44384 1458 44396
rect 2041 44387 2099 44393
rect 2041 44384 2053 44387
rect 1452 44356 2053 44384
rect 1452 44344 1458 44356
rect 2041 44353 2053 44356
rect 2087 44353 2099 44387
rect 22925 44387 22983 44393
rect 22925 44384 22937 44387
rect 2041 44347 2099 44353
rect 22296 44356 22937 44384
rect 22296 44325 22324 44356
rect 22925 44353 22937 44356
rect 22971 44353 22983 44387
rect 37829 44387 37887 44393
rect 37829 44384 37841 44387
rect 22925 44347 22983 44353
rect 26206 44356 37841 44384
rect 21821 44319 21879 44325
rect 21821 44285 21833 44319
rect 21867 44285 21879 44319
rect 21821 44279 21879 44285
rect 22281 44319 22339 44325
rect 22281 44285 22293 44319
rect 22327 44285 22339 44319
rect 22281 44279 22339 44285
rect 1581 44183 1639 44189
rect 1581 44149 1593 44183
rect 1627 44180 1639 44183
rect 1762 44180 1768 44192
rect 1627 44152 1768 44180
rect 1627 44149 1639 44152
rect 1581 44143 1639 44149
rect 1762 44140 1768 44152
rect 1820 44140 1826 44192
rect 21836 44180 21864 44279
rect 22094 44248 22100 44260
rect 22055 44220 22100 44248
rect 22094 44208 22100 44220
rect 22152 44208 22158 44260
rect 23109 44251 23167 44257
rect 23109 44217 23121 44251
rect 23155 44248 23167 44251
rect 26206 44248 26234 44356
rect 37829 44353 37841 44356
rect 37875 44353 37887 44387
rect 37829 44347 37887 44353
rect 38010 44248 38016 44260
rect 23155 44220 26234 44248
rect 37971 44220 38016 44248
rect 23155 44217 23167 44220
rect 23109 44211 23167 44217
rect 38010 44208 38016 44220
rect 38068 44208 38074 44260
rect 22462 44180 22468 44192
rect 21836 44152 22468 44180
rect 22462 44140 22468 44152
rect 22520 44180 22526 44192
rect 33321 44183 33379 44189
rect 33321 44180 33333 44183
rect 22520 44152 33333 44180
rect 22520 44140 22526 44152
rect 33321 44149 33333 44152
rect 33367 44180 33379 44183
rect 33594 44180 33600 44192
rect 33367 44152 33600 44180
rect 33367 44149 33379 44152
rect 33321 44143 33379 44149
rect 33594 44140 33600 44152
rect 33652 44140 33658 44192
rect 35526 44140 35532 44192
rect 35584 44180 35590 44192
rect 35713 44183 35771 44189
rect 35713 44180 35725 44183
rect 35584 44152 35725 44180
rect 35584 44140 35590 44152
rect 35713 44149 35725 44152
rect 35759 44180 35771 44183
rect 36078 44180 36084 44192
rect 35759 44152 36084 44180
rect 35759 44149 35771 44152
rect 35713 44143 35771 44149
rect 36078 44140 36084 44152
rect 36136 44140 36142 44192
rect 36262 44180 36268 44192
rect 36223 44152 36268 44180
rect 36262 44140 36268 44152
rect 36320 44140 36326 44192
rect 37274 44180 37280 44192
rect 37235 44152 37280 44180
rect 37274 44140 37280 44152
rect 37332 44140 37338 44192
rect 1104 44090 38824 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 38824 44090
rect 1104 44016 38824 44038
rect 22462 43976 22468 43988
rect 22423 43948 22468 43976
rect 22462 43936 22468 43948
rect 22520 43936 22526 43988
rect 36265 43979 36323 43985
rect 36265 43945 36277 43979
rect 36311 43976 36323 43979
rect 37366 43976 37372 43988
rect 36311 43948 37372 43976
rect 36311 43945 36323 43948
rect 36265 43939 36323 43945
rect 37366 43936 37372 43948
rect 37424 43936 37430 43988
rect 1394 43772 1400 43784
rect 1355 43744 1400 43772
rect 1394 43732 1400 43744
rect 1452 43772 1458 43784
rect 2041 43775 2099 43781
rect 2041 43772 2053 43775
rect 1452 43744 2053 43772
rect 1452 43732 1458 43744
rect 2041 43741 2053 43744
rect 2087 43741 2099 43775
rect 34698 43772 34704 43784
rect 34659 43744 34704 43772
rect 2041 43735 2099 43741
rect 34698 43732 34704 43744
rect 34756 43732 34762 43784
rect 37274 43772 37280 43784
rect 37235 43744 37280 43772
rect 37274 43732 37280 43744
rect 37332 43732 37338 43784
rect 37553 43775 37611 43781
rect 37553 43741 37565 43775
rect 37599 43741 37611 43775
rect 37553 43735 37611 43741
rect 23750 43664 23756 43716
rect 23808 43704 23814 43716
rect 37568 43704 37596 43735
rect 23808 43676 37596 43704
rect 23808 43664 23814 43676
rect 1581 43639 1639 43645
rect 1581 43605 1593 43639
rect 1627 43636 1639 43639
rect 2590 43636 2596 43648
rect 1627 43608 2596 43636
rect 1627 43605 1639 43608
rect 1581 43599 1639 43605
rect 2590 43596 2596 43608
rect 2648 43596 2654 43648
rect 26973 43639 27031 43645
rect 26973 43605 26985 43639
rect 27019 43636 27031 43639
rect 27982 43636 27988 43648
rect 27019 43608 27988 43636
rect 27019 43605 27031 43608
rect 26973 43599 27031 43605
rect 27982 43596 27988 43608
rect 28040 43596 28046 43648
rect 34885 43639 34943 43645
rect 34885 43605 34897 43639
rect 34931 43636 34943 43639
rect 35342 43636 35348 43648
rect 34931 43608 35348 43636
rect 34931 43605 34943 43608
rect 34885 43599 34943 43605
rect 35342 43596 35348 43608
rect 35400 43596 35406 43648
rect 36722 43636 36728 43648
rect 36683 43608 36728 43636
rect 36722 43596 36728 43608
rect 36780 43596 36786 43648
rect 1104 43546 38824 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 38824 43546
rect 1104 43472 38824 43494
rect 26142 43392 26148 43444
rect 26200 43432 26206 43444
rect 26237 43435 26295 43441
rect 26237 43432 26249 43435
rect 26200 43404 26249 43432
rect 26200 43392 26206 43404
rect 26237 43401 26249 43404
rect 26283 43401 26295 43435
rect 26237 43395 26295 43401
rect 27525 43435 27583 43441
rect 27525 43401 27537 43435
rect 27571 43432 27583 43435
rect 31570 43432 31576 43444
rect 27571 43404 31576 43432
rect 27571 43401 27583 43404
rect 27525 43395 27583 43401
rect 31570 43392 31576 43404
rect 31628 43392 31634 43444
rect 35526 43364 35532 43376
rect 6886 43336 35532 43364
rect 1394 43296 1400 43308
rect 1355 43268 1400 43296
rect 1394 43256 1400 43268
rect 1452 43296 1458 43308
rect 2041 43299 2099 43305
rect 2041 43296 2053 43299
rect 1452 43268 2053 43296
rect 1452 43256 1458 43268
rect 2041 43265 2053 43268
rect 2087 43265 2099 43299
rect 2041 43259 2099 43265
rect 5169 43299 5227 43305
rect 5169 43265 5181 43299
rect 5215 43296 5227 43299
rect 6886 43296 6914 43336
rect 35526 43324 35532 43336
rect 35584 43324 35590 43376
rect 26418 43296 26424 43308
rect 5215 43268 6914 43296
rect 26379 43268 26424 43296
rect 5215 43265 5227 43268
rect 5169 43259 5227 43265
rect 26418 43256 26424 43268
rect 26476 43256 26482 43308
rect 27433 43299 27491 43305
rect 27433 43265 27445 43299
rect 27479 43296 27491 43299
rect 30374 43296 30380 43308
rect 27479 43268 30380 43296
rect 27479 43265 27491 43268
rect 27433 43259 27491 43265
rect 30374 43256 30380 43268
rect 30432 43256 30438 43308
rect 37369 43299 37427 43305
rect 37369 43265 37381 43299
rect 37415 43296 37427 43299
rect 38010 43296 38016 43308
rect 37415 43268 38016 43296
rect 37415 43265 37427 43268
rect 37369 43259 37427 43265
rect 38010 43256 38016 43268
rect 38068 43256 38074 43308
rect 4890 43228 4896 43240
rect 4851 43200 4896 43228
rect 4890 43188 4896 43200
rect 4948 43188 4954 43240
rect 27709 43231 27767 43237
rect 27709 43197 27721 43231
rect 27755 43228 27767 43231
rect 27982 43228 27988 43240
rect 27755 43200 27988 43228
rect 27755 43197 27767 43200
rect 27709 43191 27767 43197
rect 27982 43188 27988 43200
rect 28040 43188 28046 43240
rect 1581 43163 1639 43169
rect 1581 43129 1593 43163
rect 1627 43160 1639 43163
rect 4982 43160 4988 43172
rect 1627 43132 4988 43160
rect 1627 43129 1639 43132
rect 1581 43123 1639 43129
rect 4982 43120 4988 43132
rect 5040 43120 5046 43172
rect 37642 43120 37648 43172
rect 37700 43160 37706 43172
rect 37829 43163 37887 43169
rect 37829 43160 37841 43163
rect 37700 43132 37841 43160
rect 37700 43120 37706 43132
rect 37829 43129 37841 43132
rect 37875 43129 37887 43163
rect 37829 43123 37887 43129
rect 27062 43092 27068 43104
rect 27023 43064 27068 43092
rect 27062 43052 27068 43064
rect 27120 43052 27126 43104
rect 1104 43002 38824 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 38824 43002
rect 1104 42928 38824 42950
rect 4709 42891 4767 42897
rect 4709 42857 4721 42891
rect 4755 42888 4767 42891
rect 4890 42888 4896 42900
rect 4755 42860 4896 42888
rect 4755 42857 4767 42860
rect 4709 42851 4767 42857
rect 4890 42848 4896 42860
rect 4948 42848 4954 42900
rect 4982 42848 4988 42900
rect 5040 42888 5046 42900
rect 20622 42888 20628 42900
rect 5040 42860 20628 42888
rect 5040 42848 5046 42860
rect 20622 42848 20628 42860
rect 20680 42848 20686 42900
rect 26418 42848 26424 42900
rect 26476 42888 26482 42900
rect 27433 42891 27491 42897
rect 27433 42888 27445 42891
rect 26476 42860 27445 42888
rect 26476 42848 26482 42860
rect 27433 42857 27445 42860
rect 27479 42857 27491 42891
rect 27433 42851 27491 42857
rect 4157 42755 4215 42761
rect 4157 42721 4169 42755
rect 4203 42721 4215 42755
rect 4157 42715 4215 42721
rect 4249 42755 4307 42761
rect 4249 42721 4261 42755
rect 4295 42752 4307 42755
rect 4614 42752 4620 42764
rect 4295 42724 4620 42752
rect 4295 42721 4307 42724
rect 4249 42715 4307 42721
rect 1394 42684 1400 42696
rect 1355 42656 1400 42684
rect 1394 42644 1400 42656
rect 1452 42684 1458 42696
rect 2041 42687 2099 42693
rect 2041 42684 2053 42687
rect 1452 42656 2053 42684
rect 1452 42644 1458 42656
rect 2041 42653 2053 42656
rect 2087 42653 2099 42687
rect 4172 42684 4200 42715
rect 4614 42712 4620 42724
rect 4672 42712 4678 42764
rect 12434 42712 12440 42764
rect 12492 42752 12498 42764
rect 18506 42752 18512 42764
rect 12492 42724 18512 42752
rect 12492 42712 12498 42724
rect 18506 42712 18512 42724
rect 18564 42712 18570 42764
rect 27982 42752 27988 42764
rect 27943 42724 27988 42752
rect 27982 42712 27988 42724
rect 28040 42712 28046 42764
rect 4706 42684 4712 42696
rect 4172 42656 4712 42684
rect 2041 42647 2099 42653
rect 4706 42644 4712 42656
rect 4764 42644 4770 42696
rect 26421 42687 26479 42693
rect 26421 42653 26433 42687
rect 26467 42684 26479 42687
rect 27062 42684 27068 42696
rect 26467 42656 27068 42684
rect 26467 42653 26479 42656
rect 26421 42647 26479 42653
rect 27062 42644 27068 42656
rect 27120 42644 27126 42696
rect 27893 42687 27951 42693
rect 27893 42653 27905 42687
rect 27939 42684 27951 42687
rect 37366 42684 37372 42696
rect 27939 42656 37372 42684
rect 27939 42653 27951 42656
rect 27893 42647 27951 42653
rect 37366 42644 37372 42656
rect 37424 42644 37430 42696
rect 37461 42687 37519 42693
rect 37461 42653 37473 42687
rect 37507 42684 37519 42687
rect 38102 42684 38108 42696
rect 37507 42656 38108 42684
rect 37507 42653 37519 42656
rect 37461 42647 37519 42653
rect 38102 42644 38108 42656
rect 38160 42644 38166 42696
rect 3694 42576 3700 42628
rect 3752 42616 3758 42628
rect 4341 42619 4399 42625
rect 4341 42616 4353 42619
rect 3752 42588 4353 42616
rect 3752 42576 3758 42588
rect 4341 42585 4353 42588
rect 4387 42585 4399 42619
rect 9490 42616 9496 42628
rect 4341 42579 4399 42585
rect 4448 42588 9496 42616
rect 1581 42551 1639 42557
rect 1581 42517 1593 42551
rect 1627 42548 1639 42551
rect 4448 42548 4476 42588
rect 9490 42576 9496 42588
rect 9548 42576 9554 42628
rect 27801 42619 27859 42625
rect 27801 42585 27813 42619
rect 27847 42616 27859 42619
rect 35618 42616 35624 42628
rect 27847 42588 35624 42616
rect 27847 42585 27859 42588
rect 27801 42579 27859 42585
rect 35618 42576 35624 42588
rect 35676 42576 35682 42628
rect 1627 42520 4476 42548
rect 1627 42517 1639 42520
rect 1581 42511 1639 42517
rect 4706 42508 4712 42560
rect 4764 42548 4770 42560
rect 5169 42551 5227 42557
rect 5169 42548 5181 42551
rect 4764 42520 5181 42548
rect 4764 42508 4770 42520
rect 5169 42517 5181 42520
rect 5215 42517 5227 42551
rect 5169 42511 5227 42517
rect 26329 42551 26387 42557
rect 26329 42517 26341 42551
rect 26375 42548 26387 42551
rect 26602 42548 26608 42560
rect 26375 42520 26608 42548
rect 26375 42517 26387 42520
rect 26329 42511 26387 42517
rect 26602 42508 26608 42520
rect 26660 42508 26666 42560
rect 37826 42508 37832 42560
rect 37884 42548 37890 42560
rect 37921 42551 37979 42557
rect 37921 42548 37933 42551
rect 37884 42520 37933 42548
rect 37884 42508 37890 42520
rect 37921 42517 37933 42520
rect 37967 42517 37979 42551
rect 37921 42511 37979 42517
rect 1104 42458 38824 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 38824 42458
rect 1104 42384 38824 42406
rect 20622 42304 20628 42356
rect 20680 42344 20686 42356
rect 20717 42347 20775 42353
rect 20717 42344 20729 42347
rect 20680 42316 20729 42344
rect 20680 42304 20686 42316
rect 20717 42313 20729 42316
rect 20763 42313 20775 42347
rect 27338 42344 27344 42356
rect 27299 42316 27344 42344
rect 20717 42307 20775 42313
rect 27338 42304 27344 42316
rect 27396 42304 27402 42356
rect 27154 42208 27160 42220
rect 27115 42180 27160 42208
rect 27154 42168 27160 42180
rect 27212 42168 27218 42220
rect 1673 42007 1731 42013
rect 1673 41973 1685 42007
rect 1719 42004 1731 42007
rect 1854 42004 1860 42016
rect 1719 41976 1860 42004
rect 1719 41973 1731 41976
rect 1673 41967 1731 41973
rect 1854 41964 1860 41976
rect 1912 41964 1918 42016
rect 3694 41964 3700 42016
rect 3752 42004 3758 42016
rect 3789 42007 3847 42013
rect 3789 42004 3801 42007
rect 3752 41976 3801 42004
rect 3752 41964 3758 41976
rect 3789 41973 3801 41976
rect 3835 41973 3847 42007
rect 3789 41967 3847 41973
rect 26142 41964 26148 42016
rect 26200 42004 26206 42016
rect 27801 42007 27859 42013
rect 27801 42004 27813 42007
rect 26200 41976 27813 42004
rect 26200 41964 26206 41976
rect 27801 41973 27813 41976
rect 27847 42004 27859 42007
rect 27982 42004 27988 42016
rect 27847 41976 27988 42004
rect 27847 41973 27859 41976
rect 27801 41967 27859 41973
rect 27982 41964 27988 41976
rect 28040 41964 28046 42016
rect 1104 41914 38824 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 38824 41914
rect 1104 41840 38824 41862
rect 22557 41803 22615 41809
rect 22557 41769 22569 41803
rect 22603 41800 22615 41803
rect 26970 41800 26976 41812
rect 22603 41772 26976 41800
rect 22603 41769 22615 41772
rect 22557 41763 22615 41769
rect 26970 41760 26976 41772
rect 27028 41760 27034 41812
rect 37366 41760 37372 41812
rect 37424 41800 37430 41812
rect 37921 41803 37979 41809
rect 37921 41800 37933 41803
rect 37424 41772 37933 41800
rect 37424 41760 37430 41772
rect 37921 41769 37933 41772
rect 37967 41769 37979 41803
rect 37921 41763 37979 41769
rect 20717 41667 20775 41673
rect 20717 41633 20729 41667
rect 20763 41664 20775 41667
rect 21361 41667 21419 41673
rect 21361 41664 21373 41667
rect 20763 41636 21373 41664
rect 20763 41633 20775 41636
rect 20717 41627 20775 41633
rect 21361 41633 21373 41636
rect 21407 41664 21419 41667
rect 21634 41664 21640 41676
rect 21407 41636 21640 41664
rect 21407 41633 21419 41636
rect 21361 41627 21419 41633
rect 21634 41624 21640 41636
rect 21692 41624 21698 41676
rect 1854 41596 1860 41608
rect 1815 41568 1860 41596
rect 1854 41556 1860 41568
rect 1912 41556 1918 41608
rect 20622 41556 20628 41608
rect 20680 41596 20686 41608
rect 21453 41599 21511 41605
rect 21453 41596 21465 41599
rect 20680 41568 21465 41596
rect 20680 41556 20686 41568
rect 21453 41565 21465 41568
rect 21499 41565 21511 41599
rect 22373 41599 22431 41605
rect 22373 41596 22385 41599
rect 21453 41559 21511 41565
rect 21928 41568 22385 41596
rect 2041 41531 2099 41537
rect 2041 41497 2053 41531
rect 2087 41528 2099 41531
rect 4062 41528 4068 41540
rect 2087 41500 4068 41528
rect 2087 41497 2099 41500
rect 2041 41491 2099 41497
rect 4062 41488 4068 41500
rect 4120 41488 4126 41540
rect 21545 41463 21603 41469
rect 21545 41429 21557 41463
rect 21591 41460 21603 41463
rect 21726 41460 21732 41472
rect 21591 41432 21732 41460
rect 21591 41429 21603 41432
rect 21545 41423 21603 41429
rect 21726 41420 21732 41432
rect 21784 41420 21790 41472
rect 21928 41469 21956 41568
rect 22373 41565 22385 41568
rect 22419 41565 22431 41599
rect 22373 41559 22431 41565
rect 37461 41599 37519 41605
rect 37461 41565 37473 41599
rect 37507 41596 37519 41599
rect 38102 41596 38108 41608
rect 37507 41568 38108 41596
rect 37507 41565 37519 41568
rect 37461 41559 37519 41565
rect 38102 41556 38108 41568
rect 38160 41556 38166 41608
rect 21913 41463 21971 41469
rect 21913 41429 21925 41463
rect 21959 41429 21971 41463
rect 21913 41423 21971 41429
rect 1104 41370 38824 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 38824 41370
rect 1104 41296 38824 41318
rect 27154 41216 27160 41268
rect 27212 41256 27218 41268
rect 27525 41259 27583 41265
rect 27525 41256 27537 41259
rect 27212 41228 27537 41256
rect 27212 41216 27218 41228
rect 27525 41225 27537 41228
rect 27571 41225 27583 41259
rect 28721 41259 28779 41265
rect 28721 41256 28733 41259
rect 27525 41219 27583 41225
rect 27908 41228 28733 41256
rect 27338 41080 27344 41132
rect 27396 41120 27402 41132
rect 27908 41129 27936 41228
rect 28721 41225 28733 41228
rect 28767 41256 28779 41259
rect 35710 41256 35716 41268
rect 28767 41228 35716 41256
rect 28767 41225 28779 41228
rect 28721 41219 28779 41225
rect 35710 41216 35716 41228
rect 35768 41216 35774 41268
rect 27985 41191 28043 41197
rect 27985 41157 27997 41191
rect 28031 41188 28043 41191
rect 28031 41160 35894 41188
rect 28031 41157 28043 41160
rect 27985 41151 28043 41157
rect 27893 41123 27951 41129
rect 27893 41120 27905 41123
rect 27396 41092 27905 41120
rect 27396 41080 27402 41092
rect 27893 41089 27905 41092
rect 27939 41089 27951 41123
rect 27893 41083 27951 41089
rect 1949 41055 2007 41061
rect 1949 41021 1961 41055
rect 1995 41021 2007 41055
rect 2222 41052 2228 41064
rect 2183 41024 2228 41052
rect 1949 41015 2007 41021
rect 1964 40984 1992 41015
rect 2222 41012 2228 41024
rect 2280 41052 2286 41064
rect 2685 41055 2743 41061
rect 2685 41052 2697 41055
rect 2280 41024 2697 41052
rect 2280 41012 2286 41024
rect 2685 41021 2697 41024
rect 2731 41021 2743 41055
rect 2685 41015 2743 41021
rect 21634 41012 21640 41064
rect 21692 41052 21698 41064
rect 26973 41055 27031 41061
rect 26973 41052 26985 41055
rect 21692 41024 26985 41052
rect 21692 41012 21698 41024
rect 26973 41021 26985 41024
rect 27019 41052 27031 41055
rect 28077 41055 28135 41061
rect 28077 41052 28089 41055
rect 27019 41024 28089 41052
rect 27019 41021 27031 41024
rect 26973 41015 27031 41021
rect 28077 41021 28089 41024
rect 28123 41021 28135 41055
rect 28077 41015 28135 41021
rect 19242 40984 19248 40996
rect 1964 40956 19248 40984
rect 19242 40944 19248 40956
rect 19300 40944 19306 40996
rect 35866 40984 35894 41160
rect 37461 41123 37519 41129
rect 37461 41089 37473 41123
rect 37507 41120 37519 41123
rect 38102 41120 38108 41132
rect 37507 41092 38108 41120
rect 37507 41089 37519 41092
rect 37461 41083 37519 41089
rect 38102 41080 38108 41092
rect 38160 41080 38166 41132
rect 37921 40987 37979 40993
rect 37921 40984 37933 40987
rect 35866 40956 37933 40984
rect 37921 40953 37933 40956
rect 37967 40953 37979 40987
rect 37921 40947 37979 40953
rect 20898 40916 20904 40928
rect 20859 40888 20904 40916
rect 20898 40876 20904 40888
rect 20956 40916 20962 40928
rect 21726 40916 21732 40928
rect 20956 40888 21732 40916
rect 20956 40876 20962 40888
rect 21726 40876 21732 40888
rect 21784 40876 21790 40928
rect 1104 40826 38824 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 38824 40826
rect 1104 40752 38824 40774
rect 37461 40511 37519 40517
rect 37461 40477 37473 40511
rect 37507 40508 37519 40511
rect 38102 40508 38108 40520
rect 37507 40480 38108 40508
rect 37507 40477 37519 40480
rect 37461 40471 37519 40477
rect 38102 40468 38108 40480
rect 38160 40468 38166 40520
rect 1854 40440 1860 40452
rect 1815 40412 1860 40440
rect 1854 40400 1860 40412
rect 1912 40400 1918 40452
rect 2038 40440 2044 40452
rect 1999 40412 2044 40440
rect 2038 40400 2044 40412
rect 2096 40400 2102 40452
rect 22738 40400 22744 40452
rect 22796 40440 22802 40452
rect 22796 40412 37964 40440
rect 22796 40400 22802 40412
rect 1872 40372 1900 40400
rect 37936 40381 37964 40412
rect 2501 40375 2559 40381
rect 2501 40372 2513 40375
rect 1872 40344 2513 40372
rect 2501 40341 2513 40344
rect 2547 40341 2559 40375
rect 2501 40335 2559 40341
rect 37921 40375 37979 40381
rect 37921 40341 37933 40375
rect 37967 40341 37979 40375
rect 37921 40335 37979 40341
rect 1104 40282 38824 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 38824 40282
rect 1104 40208 38824 40230
rect 37369 40035 37427 40041
rect 37369 40001 37381 40035
rect 37415 40032 37427 40035
rect 37829 40035 37887 40041
rect 37829 40032 37841 40035
rect 37415 40004 37841 40032
rect 37415 40001 37427 40004
rect 37369 39995 37427 40001
rect 37829 40001 37841 40004
rect 37875 40032 37887 40035
rect 38286 40032 38292 40044
rect 37875 40004 38292 40032
rect 37875 40001 37887 40004
rect 37829 39995 37887 40001
rect 38286 39992 38292 40004
rect 38344 39992 38350 40044
rect 1394 39964 1400 39976
rect 1355 39936 1400 39964
rect 1394 39924 1400 39936
rect 1452 39924 1458 39976
rect 1578 39924 1584 39976
rect 1636 39964 1642 39976
rect 1673 39967 1731 39973
rect 1673 39964 1685 39967
rect 1636 39936 1685 39964
rect 1636 39924 1642 39936
rect 1673 39933 1685 39936
rect 1719 39933 1731 39967
rect 1673 39927 1731 39933
rect 38010 39828 38016 39840
rect 37971 39800 38016 39828
rect 38010 39788 38016 39800
rect 38068 39788 38074 39840
rect 1104 39738 38824 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 38824 39738
rect 1104 39664 38824 39686
rect 21910 39584 21916 39636
rect 21968 39624 21974 39636
rect 22649 39627 22707 39633
rect 22649 39624 22661 39627
rect 21968 39596 22661 39624
rect 21968 39584 21974 39596
rect 22649 39593 22661 39596
rect 22695 39624 22707 39627
rect 24854 39624 24860 39636
rect 22695 39596 24860 39624
rect 22695 39593 22707 39596
rect 22649 39587 22707 39593
rect 24854 39584 24860 39596
rect 24912 39584 24918 39636
rect 1394 39556 1400 39568
rect 1355 39528 1400 39556
rect 1394 39516 1400 39528
rect 1452 39516 1458 39568
rect 20257 39491 20315 39497
rect 20257 39457 20269 39491
rect 20303 39488 20315 39491
rect 20806 39488 20812 39500
rect 20303 39460 20812 39488
rect 20303 39457 20315 39460
rect 20257 39451 20315 39457
rect 20806 39448 20812 39460
rect 20864 39488 20870 39500
rect 21910 39488 21916 39500
rect 20864 39460 21916 39488
rect 20864 39448 20870 39460
rect 21910 39448 21916 39460
rect 21968 39448 21974 39500
rect 2682 39380 2688 39432
rect 2740 39420 2746 39432
rect 10318 39420 10324 39432
rect 2740 39392 10324 39420
rect 2740 39380 2746 39392
rect 10318 39380 10324 39392
rect 10376 39380 10382 39432
rect 19426 39380 19432 39432
rect 19484 39420 19490 39432
rect 19613 39423 19671 39429
rect 19613 39420 19625 39423
rect 19484 39392 19625 39420
rect 19484 39380 19490 39392
rect 19613 39389 19625 39392
rect 19659 39389 19671 39423
rect 20622 39420 20628 39432
rect 20583 39392 20628 39420
rect 19613 39383 19671 39389
rect 20622 39380 20628 39392
rect 20680 39380 20686 39432
rect 22002 39380 22008 39432
rect 22060 39429 22066 39432
rect 22060 39423 22109 39429
rect 22060 39389 22063 39423
rect 22097 39420 22109 39423
rect 22097 39392 22153 39420
rect 22097 39389 22109 39392
rect 22060 39383 22109 39389
rect 22060 39380 22066 39383
rect 1946 39312 1952 39364
rect 2004 39352 2010 39364
rect 12250 39352 12256 39364
rect 2004 39324 12256 39352
rect 2004 39312 2010 39324
rect 12250 39312 12256 39324
rect 12308 39312 12314 39364
rect 20990 39312 20996 39364
rect 21048 39312 21054 39364
rect 1104 39194 38824 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 38824 39194
rect 1104 39120 38824 39142
rect 20622 39040 20628 39092
rect 20680 39080 20686 39092
rect 21131 39083 21189 39089
rect 21131 39080 21143 39083
rect 20680 39052 21143 39080
rect 20680 39040 20686 39052
rect 21131 39049 21143 39052
rect 21177 39049 21189 39083
rect 21131 39043 21189 39049
rect 21913 39015 21971 39021
rect 21913 39012 21925 39015
rect 20746 38984 21925 39012
rect 21913 38981 21925 38984
rect 21959 38981 21971 39015
rect 21913 38975 21971 38981
rect 1673 38947 1731 38953
rect 1673 38913 1685 38947
rect 1719 38944 1731 38947
rect 2225 38947 2283 38953
rect 2225 38944 2237 38947
rect 1719 38916 2237 38944
rect 1719 38913 1731 38916
rect 1673 38907 1731 38913
rect 2225 38913 2237 38916
rect 2271 38944 2283 38947
rect 15470 38944 15476 38956
rect 2271 38916 15476 38944
rect 2271 38913 2283 38916
rect 2225 38907 2283 38913
rect 15470 38904 15476 38916
rect 15528 38904 15534 38956
rect 19426 38904 19432 38956
rect 19484 38944 19490 38956
rect 19705 38947 19763 38953
rect 19705 38944 19717 38947
rect 19484 38916 19717 38944
rect 19484 38904 19490 38916
rect 19705 38913 19717 38916
rect 19751 38913 19763 38947
rect 19705 38907 19763 38913
rect 21266 38904 21272 38956
rect 21324 38944 21330 38956
rect 22005 38947 22063 38953
rect 22005 38944 22017 38947
rect 21324 38916 22017 38944
rect 21324 38904 21330 38916
rect 22005 38913 22017 38916
rect 22051 38944 22063 38947
rect 22465 38947 22523 38953
rect 22465 38944 22477 38947
rect 22051 38916 22477 38944
rect 22051 38913 22063 38916
rect 22005 38907 22063 38913
rect 22465 38913 22477 38916
rect 22511 38913 22523 38947
rect 37829 38947 37887 38953
rect 37829 38944 37841 38947
rect 22465 38907 22523 38913
rect 37292 38916 37841 38944
rect 19337 38879 19395 38885
rect 19337 38845 19349 38879
rect 19383 38876 19395 38879
rect 20806 38876 20812 38888
rect 19383 38848 20812 38876
rect 19383 38845 19395 38848
rect 19337 38839 19395 38845
rect 20806 38836 20812 38848
rect 20864 38836 20870 38888
rect 1486 38808 1492 38820
rect 1447 38780 1492 38808
rect 1486 38768 1492 38780
rect 1544 38768 1550 38820
rect 27614 38700 27620 38752
rect 27672 38740 27678 38752
rect 37292 38749 37320 38916
rect 37829 38913 37841 38916
rect 37875 38913 37887 38947
rect 37829 38907 37887 38913
rect 38010 38808 38016 38820
rect 37971 38780 38016 38808
rect 38010 38768 38016 38780
rect 38068 38768 38074 38820
rect 37277 38743 37335 38749
rect 37277 38740 37289 38743
rect 27672 38712 37289 38740
rect 27672 38700 27678 38712
rect 37277 38709 37289 38712
rect 37323 38709 37335 38743
rect 37277 38703 37335 38709
rect 1104 38650 38824 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 38824 38650
rect 1104 38576 38824 38598
rect 20717 38539 20775 38545
rect 20717 38505 20729 38539
rect 20763 38536 20775 38539
rect 20990 38536 20996 38548
rect 20763 38508 20996 38536
rect 20763 38505 20775 38508
rect 20717 38499 20775 38505
rect 20990 38496 20996 38508
rect 21048 38496 21054 38548
rect 21910 38536 21916 38548
rect 21871 38508 21916 38536
rect 21910 38496 21916 38508
rect 21968 38496 21974 38548
rect 1949 38335 2007 38341
rect 1949 38301 1961 38335
rect 1995 38301 2007 38335
rect 2222 38332 2228 38344
rect 2183 38304 2228 38332
rect 1949 38295 2007 38301
rect 1964 38264 1992 38295
rect 2222 38292 2228 38304
rect 2280 38332 2286 38344
rect 2685 38335 2743 38341
rect 2685 38332 2697 38335
rect 2280 38304 2697 38332
rect 2280 38292 2286 38304
rect 2685 38301 2697 38304
rect 2731 38301 2743 38335
rect 2685 38295 2743 38301
rect 14458 38292 14464 38344
rect 14516 38332 14522 38344
rect 15010 38332 15016 38344
rect 14516 38304 15016 38332
rect 14516 38292 14522 38304
rect 15010 38292 15016 38304
rect 15068 38332 15074 38344
rect 20625 38335 20683 38341
rect 20625 38332 20637 38335
rect 15068 38304 20637 38332
rect 15068 38292 15074 38304
rect 20625 38301 20637 38304
rect 20671 38332 20683 38335
rect 21266 38332 21272 38344
rect 20671 38304 21272 38332
rect 20671 38301 20683 38304
rect 20625 38295 20683 38301
rect 21266 38292 21272 38304
rect 21324 38292 21330 38344
rect 37461 38335 37519 38341
rect 37461 38301 37473 38335
rect 37507 38332 37519 38335
rect 38102 38332 38108 38344
rect 37507 38304 38108 38332
rect 37507 38301 37519 38304
rect 37461 38295 37519 38301
rect 38102 38292 38108 38304
rect 38160 38292 38166 38344
rect 20990 38264 20996 38276
rect 1964 38236 20996 38264
rect 20990 38224 20996 38236
rect 21048 38224 21054 38276
rect 37734 38156 37740 38208
rect 37792 38196 37798 38208
rect 37921 38199 37979 38205
rect 37921 38196 37933 38199
rect 37792 38168 37933 38196
rect 37792 38156 37798 38168
rect 37921 38165 37933 38168
rect 37967 38165 37979 38199
rect 37921 38159 37979 38165
rect 1104 38106 38824 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 38824 38106
rect 1104 38032 38824 38054
rect 8386 37992 8392 38004
rect 8347 37964 8392 37992
rect 8386 37952 8392 37964
rect 8444 37952 8450 38004
rect 15470 37952 15476 38004
rect 15528 37992 15534 38004
rect 22278 37992 22284 38004
rect 15528 37964 22284 37992
rect 15528 37952 15534 37964
rect 22278 37952 22284 37964
rect 22336 37952 22342 38004
rect 4062 37884 4068 37936
rect 4120 37924 4126 37936
rect 24946 37924 24952 37936
rect 4120 37896 24952 37924
rect 4120 37884 4126 37896
rect 24946 37884 24952 37896
rect 25004 37884 25010 37936
rect 8570 37856 8576 37868
rect 8531 37828 8576 37856
rect 8570 37816 8576 37828
rect 8628 37816 8634 37868
rect 35342 37816 35348 37868
rect 35400 37856 35406 37868
rect 37829 37859 37887 37865
rect 37829 37856 37841 37859
rect 35400 37828 37841 37856
rect 35400 37816 35406 37828
rect 37829 37825 37841 37828
rect 37875 37825 37887 37859
rect 37829 37819 37887 37825
rect 1949 37791 2007 37797
rect 1949 37757 1961 37791
rect 1995 37757 2007 37791
rect 2222 37788 2228 37800
rect 2183 37760 2228 37788
rect 1949 37751 2007 37757
rect 1964 37720 1992 37751
rect 2222 37748 2228 37760
rect 2280 37788 2286 37800
rect 2685 37791 2743 37797
rect 2685 37788 2697 37791
rect 2280 37760 2697 37788
rect 2280 37748 2286 37760
rect 2685 37757 2697 37760
rect 2731 37757 2743 37791
rect 2685 37751 2743 37757
rect 22554 37720 22560 37732
rect 1964 37692 22560 37720
rect 22554 37680 22560 37692
rect 22612 37680 22618 37732
rect 38010 37652 38016 37664
rect 37971 37624 38016 37652
rect 38010 37612 38016 37624
rect 38068 37612 38074 37664
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 8570 37408 8576 37460
rect 8628 37448 8634 37460
rect 9033 37451 9091 37457
rect 9033 37448 9045 37451
rect 8628 37420 9045 37448
rect 8628 37408 8634 37420
rect 9033 37417 9045 37420
rect 9079 37417 9091 37451
rect 22738 37448 22744 37460
rect 22699 37420 22744 37448
rect 9033 37411 9091 37417
rect 22738 37408 22744 37420
rect 22796 37408 22802 37460
rect 9585 37315 9643 37321
rect 9585 37281 9597 37315
rect 9631 37312 9643 37315
rect 9950 37312 9956 37324
rect 9631 37284 9956 37312
rect 9631 37281 9643 37284
rect 9585 37275 9643 37281
rect 9950 37272 9956 37284
rect 10008 37272 10014 37324
rect 1673 37247 1731 37253
rect 1673 37213 1685 37247
rect 1719 37244 1731 37247
rect 9490 37244 9496 37256
rect 1719 37216 2176 37244
rect 9451 37216 9496 37244
rect 1719 37213 1731 37216
rect 1673 37207 1731 37213
rect 2148 37120 2176 37216
rect 9490 37204 9496 37216
rect 9548 37204 9554 37256
rect 22005 37247 22063 37253
rect 22005 37213 22017 37247
rect 22051 37244 22063 37247
rect 22094 37244 22100 37256
rect 22051 37216 22100 37244
rect 22051 37213 22063 37216
rect 22005 37207 22063 37213
rect 22094 37204 22100 37216
rect 22152 37204 22158 37256
rect 37829 37247 37887 37253
rect 37829 37244 37841 37247
rect 31726 37216 37841 37244
rect 9401 37179 9459 37185
rect 9401 37145 9413 37179
rect 9447 37176 9459 37179
rect 10321 37179 10379 37185
rect 10321 37176 10333 37179
rect 9447 37148 10333 37176
rect 9447 37145 9459 37148
rect 9401 37139 9459 37145
rect 10321 37145 10333 37148
rect 10367 37176 10379 37179
rect 31726 37176 31754 37216
rect 37829 37213 37841 37216
rect 37875 37213 37887 37247
rect 38102 37244 38108 37256
rect 38063 37216 38108 37244
rect 37829 37207 37887 37213
rect 38102 37204 38108 37216
rect 38160 37204 38166 37256
rect 10367 37148 31754 37176
rect 10367 37145 10379 37148
rect 10321 37139 10379 37145
rect 1486 37108 1492 37120
rect 1447 37080 1492 37108
rect 1486 37068 1492 37080
rect 1544 37068 1550 37120
rect 2130 37108 2136 37120
rect 2091 37080 2136 37108
rect 2130 37068 2136 37080
rect 2188 37068 2194 37120
rect 22189 37111 22247 37117
rect 22189 37077 22201 37111
rect 22235 37108 22247 37111
rect 31478 37108 31484 37120
rect 22235 37080 31484 37108
rect 22235 37077 22247 37080
rect 22189 37071 22247 37077
rect 31478 37068 31484 37080
rect 31536 37068 31542 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 22186 36904 22192 36916
rect 22147 36876 22192 36904
rect 22186 36864 22192 36876
rect 22244 36864 22250 36916
rect 22281 36907 22339 36913
rect 22281 36873 22293 36907
rect 22327 36904 22339 36907
rect 22738 36904 22744 36916
rect 22327 36876 22744 36904
rect 22327 36873 22339 36876
rect 22281 36867 22339 36873
rect 22738 36864 22744 36876
rect 22796 36864 22802 36916
rect 23474 36904 23480 36916
rect 23435 36876 23480 36904
rect 23474 36864 23480 36876
rect 23532 36864 23538 36916
rect 38102 36836 38108 36848
rect 38063 36808 38108 36836
rect 38102 36796 38108 36808
rect 38160 36796 38166 36848
rect 21726 36700 21732 36712
rect 21192 36672 21732 36700
rect 9950 36564 9956 36576
rect 9863 36536 9956 36564
rect 9950 36524 9956 36536
rect 10008 36564 10014 36576
rect 21192 36573 21220 36672
rect 21726 36660 21732 36672
rect 21784 36700 21790 36712
rect 22373 36703 22431 36709
rect 22373 36700 22385 36703
rect 21784 36672 22385 36700
rect 21784 36660 21790 36672
rect 22373 36669 22385 36672
rect 22419 36669 22431 36703
rect 22373 36663 22431 36669
rect 21177 36567 21235 36573
rect 21177 36564 21189 36567
rect 10008 36536 21189 36564
rect 10008 36524 10014 36536
rect 21177 36533 21189 36536
rect 21223 36533 21235 36567
rect 21818 36564 21824 36576
rect 21779 36536 21824 36564
rect 21177 36527 21235 36533
rect 21818 36524 21824 36536
rect 21876 36524 21882 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 22094 36320 22100 36372
rect 22152 36360 22158 36372
rect 23750 36360 23756 36372
rect 22152 36332 22197 36360
rect 23711 36332 23756 36360
rect 22152 36320 22158 36332
rect 23750 36320 23756 36332
rect 23808 36320 23814 36372
rect 24302 36320 24308 36372
rect 24360 36360 24366 36372
rect 24397 36363 24455 36369
rect 24397 36360 24409 36363
rect 24360 36332 24409 36360
rect 24360 36320 24366 36332
rect 24397 36329 24409 36332
rect 24443 36329 24455 36363
rect 24397 36323 24455 36329
rect 22002 36252 22008 36304
rect 22060 36292 22066 36304
rect 23109 36295 23167 36301
rect 23109 36292 23121 36295
rect 22060 36264 23121 36292
rect 22060 36252 22066 36264
rect 23109 36261 23121 36264
rect 23155 36261 23167 36295
rect 23109 36255 23167 36261
rect 21545 36227 21603 36233
rect 21545 36193 21557 36227
rect 21591 36224 21603 36227
rect 21591 36196 22692 36224
rect 21591 36193 21603 36196
rect 21545 36187 21603 36193
rect 1670 36156 1676 36168
rect 1631 36128 1676 36156
rect 1670 36116 1676 36128
rect 1728 36116 1734 36168
rect 21637 36159 21695 36165
rect 21637 36125 21649 36159
rect 21683 36156 21695 36159
rect 22002 36156 22008 36168
rect 21683 36128 22008 36156
rect 21683 36125 21695 36128
rect 21637 36119 21695 36125
rect 22002 36116 22008 36128
rect 22060 36116 22066 36168
rect 1486 36020 1492 36032
rect 1447 35992 1492 36020
rect 1486 35980 1492 35992
rect 1544 35980 1550 36032
rect 17218 35980 17224 36032
rect 17276 36020 17282 36032
rect 22664 36029 22692 36196
rect 35986 36116 35992 36168
rect 36044 36156 36050 36168
rect 37829 36159 37887 36165
rect 37829 36156 37841 36159
rect 36044 36128 37841 36156
rect 36044 36116 36050 36128
rect 37829 36125 37841 36128
rect 37875 36125 37887 36159
rect 37829 36119 37887 36125
rect 20809 36023 20867 36029
rect 20809 36020 20821 36023
rect 17276 35992 20821 36020
rect 17276 35980 17282 35992
rect 20809 35989 20821 35992
rect 20855 36020 20867 36023
rect 21729 36023 21787 36029
rect 21729 36020 21741 36023
rect 20855 35992 21741 36020
rect 20855 35989 20867 35992
rect 20809 35983 20867 35989
rect 21729 35989 21741 35992
rect 21775 35989 21787 36023
rect 21729 35983 21787 35989
rect 22649 36023 22707 36029
rect 22649 35989 22661 36023
rect 22695 36020 22707 36023
rect 23014 36020 23020 36032
rect 22695 35992 23020 36020
rect 22695 35989 22707 35992
rect 22649 35983 22707 35989
rect 23014 35980 23020 35992
rect 23072 35980 23078 36032
rect 38010 36020 38016 36032
rect 37971 35992 38016 36020
rect 38010 35980 38016 35992
rect 38068 35980 38074 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 6917 35819 6975 35825
rect 6917 35785 6929 35819
rect 6963 35785 6975 35819
rect 6917 35779 6975 35785
rect 7561 35819 7619 35825
rect 7561 35785 7573 35819
rect 7607 35785 7619 35819
rect 7561 35779 7619 35785
rect 22925 35819 22983 35825
rect 22925 35785 22937 35819
rect 22971 35816 22983 35819
rect 23474 35816 23480 35828
rect 22971 35788 23480 35816
rect 22971 35785 22983 35788
rect 22925 35779 22983 35785
rect 1673 35683 1731 35689
rect 1673 35649 1685 35683
rect 1719 35680 1731 35683
rect 6932 35680 6960 35779
rect 1719 35652 6960 35680
rect 7101 35683 7159 35689
rect 1719 35649 1731 35652
rect 1673 35643 1731 35649
rect 7101 35649 7113 35683
rect 7147 35680 7159 35683
rect 7576 35680 7604 35779
rect 23474 35776 23480 35788
rect 23532 35776 23538 35828
rect 24302 35776 24308 35828
rect 24360 35816 24366 35828
rect 24397 35819 24455 35825
rect 24397 35816 24409 35819
rect 24360 35788 24409 35816
rect 24360 35776 24366 35788
rect 24397 35785 24409 35788
rect 24443 35785 24455 35819
rect 24397 35779 24455 35785
rect 24489 35819 24547 35825
rect 24489 35785 24501 35819
rect 24535 35816 24547 35819
rect 28442 35816 28448 35828
rect 24535 35788 28448 35816
rect 24535 35785 24547 35788
rect 24489 35779 24547 35785
rect 28442 35776 28448 35788
rect 28500 35776 28506 35828
rect 22833 35751 22891 35757
rect 22833 35717 22845 35751
rect 22879 35748 22891 35751
rect 23750 35748 23756 35760
rect 22879 35720 23756 35748
rect 22879 35717 22891 35720
rect 22833 35711 22891 35717
rect 23750 35708 23756 35720
rect 23808 35708 23814 35760
rect 7147 35652 7604 35680
rect 7929 35683 7987 35689
rect 7147 35649 7159 35652
rect 7101 35643 7159 35649
rect 7929 35649 7941 35683
rect 7975 35680 7987 35683
rect 8754 35680 8760 35692
rect 7975 35652 8760 35680
rect 7975 35649 7987 35652
rect 7929 35643 7987 35649
rect 8754 35640 8760 35652
rect 8812 35640 8818 35692
rect 37461 35683 37519 35689
rect 37461 35649 37473 35683
rect 37507 35680 37519 35683
rect 38102 35680 38108 35692
rect 37507 35652 38108 35680
rect 37507 35649 37519 35652
rect 37461 35643 37519 35649
rect 38102 35640 38108 35652
rect 38160 35640 38166 35692
rect 6546 35572 6552 35624
rect 6604 35612 6610 35624
rect 8021 35615 8079 35621
rect 8021 35612 8033 35615
rect 6604 35584 8033 35612
rect 6604 35572 6610 35584
rect 8021 35581 8033 35584
rect 8067 35581 8079 35615
rect 8021 35575 8079 35581
rect 8205 35615 8263 35621
rect 8205 35581 8217 35615
rect 8251 35612 8263 35615
rect 8251 35584 9444 35612
rect 8251 35581 8263 35584
rect 8205 35575 8263 35581
rect 5442 35504 5448 35556
rect 5500 35544 5506 35556
rect 8220 35544 8248 35575
rect 5500 35516 8248 35544
rect 5500 35504 5506 35516
rect 1486 35476 1492 35488
rect 1447 35448 1492 35476
rect 1486 35436 1492 35448
rect 1544 35436 1550 35488
rect 2222 35476 2228 35488
rect 2183 35448 2228 35476
rect 2222 35436 2228 35448
rect 2280 35436 2286 35488
rect 8754 35476 8760 35488
rect 8715 35448 8760 35476
rect 8754 35436 8760 35448
rect 8812 35436 8818 35488
rect 9416 35485 9444 35584
rect 21634 35572 21640 35624
rect 21692 35612 21698 35624
rect 21913 35615 21971 35621
rect 21913 35612 21925 35615
rect 21692 35584 21925 35612
rect 21692 35572 21698 35584
rect 21913 35581 21925 35584
rect 21959 35612 21971 35615
rect 22002 35612 22008 35624
rect 21959 35584 22008 35612
rect 21959 35581 21971 35584
rect 21913 35575 21971 35581
rect 22002 35572 22008 35584
rect 22060 35612 22066 35624
rect 23017 35615 23075 35621
rect 23017 35612 23029 35615
rect 22060 35584 23029 35612
rect 22060 35572 22066 35584
rect 23017 35581 23029 35584
rect 23063 35581 23075 35615
rect 23017 35575 23075 35581
rect 23106 35572 23112 35624
rect 23164 35612 23170 35624
rect 24213 35615 24271 35621
rect 24213 35612 24225 35615
rect 23164 35584 24225 35612
rect 23164 35572 23170 35584
rect 24213 35581 24225 35584
rect 24259 35612 24271 35615
rect 25317 35615 25375 35621
rect 25317 35612 25329 35615
rect 24259 35584 25329 35612
rect 24259 35581 24271 35584
rect 24213 35575 24271 35581
rect 25317 35581 25329 35584
rect 25363 35581 25375 35615
rect 25317 35575 25375 35581
rect 9401 35479 9459 35485
rect 9401 35445 9413 35479
rect 9447 35476 9459 35479
rect 15194 35476 15200 35488
rect 9447 35448 15200 35476
rect 9447 35445 9459 35448
rect 9401 35439 9459 35445
rect 15194 35436 15200 35448
rect 15252 35436 15258 35488
rect 22370 35436 22376 35488
rect 22428 35476 22434 35488
rect 22465 35479 22523 35485
rect 22465 35476 22477 35479
rect 22428 35448 22477 35476
rect 22428 35436 22434 35448
rect 22465 35445 22477 35448
rect 22511 35445 22523 35479
rect 24854 35476 24860 35488
rect 24815 35448 24860 35476
rect 22465 35439 22523 35445
rect 24854 35436 24860 35448
rect 24912 35436 24918 35488
rect 37918 35476 37924 35488
rect 37879 35448 37924 35476
rect 37918 35436 37924 35448
rect 37976 35436 37982 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 1670 35232 1676 35284
rect 1728 35272 1734 35284
rect 2133 35275 2191 35281
rect 2133 35272 2145 35275
rect 1728 35244 2145 35272
rect 1728 35232 1734 35244
rect 2133 35241 2145 35244
rect 2179 35241 2191 35275
rect 2133 35235 2191 35241
rect 22649 35275 22707 35281
rect 22649 35241 22661 35275
rect 22695 35272 22707 35275
rect 23293 35275 23351 35281
rect 23293 35272 23305 35275
rect 22695 35244 23305 35272
rect 22695 35241 22707 35244
rect 22649 35235 22707 35241
rect 23293 35241 23305 35244
rect 23339 35272 23351 35275
rect 27338 35272 27344 35284
rect 23339 35244 27344 35272
rect 23339 35241 23351 35244
rect 23293 35235 23351 35241
rect 27338 35232 27344 35244
rect 27396 35232 27402 35284
rect 2222 35136 2228 35148
rect 1688 35108 2228 35136
rect 1688 35077 1716 35108
rect 2222 35096 2228 35108
rect 2280 35136 2286 35148
rect 22557 35139 22615 35145
rect 2280 35108 6914 35136
rect 2280 35096 2286 35108
rect 1673 35071 1731 35077
rect 1673 35037 1685 35071
rect 1719 35037 1731 35071
rect 2314 35068 2320 35080
rect 2275 35040 2320 35068
rect 1673 35031 1731 35037
rect 2314 35028 2320 35040
rect 2372 35028 2378 35080
rect 6886 35068 6914 35108
rect 22557 35105 22569 35139
rect 22603 35136 22615 35139
rect 23750 35136 23756 35148
rect 22603 35108 23756 35136
rect 22603 35105 22615 35108
rect 22557 35099 22615 35105
rect 23750 35096 23756 35108
rect 23808 35096 23814 35148
rect 20806 35068 20812 35080
rect 6886 35040 20812 35068
rect 20806 35028 20812 35040
rect 20864 35028 20870 35080
rect 20898 35028 20904 35080
rect 20956 35068 20962 35080
rect 21913 35071 21971 35077
rect 21913 35068 21925 35071
rect 20956 35040 21925 35068
rect 20956 35028 20962 35040
rect 21913 35037 21925 35040
rect 21959 35068 21971 35071
rect 22373 35071 22431 35077
rect 22373 35068 22385 35071
rect 21959 35040 22385 35068
rect 21959 35037 21971 35040
rect 21913 35031 21971 35037
rect 22373 35037 22385 35040
rect 22419 35037 22431 35071
rect 22373 35031 22431 35037
rect 22649 35071 22707 35077
rect 22649 35037 22661 35071
rect 22695 35037 22707 35071
rect 24854 35068 24860 35080
rect 24815 35040 24860 35068
rect 22649 35031 22707 35037
rect 21361 35003 21419 35009
rect 21361 34969 21373 35003
rect 21407 35000 21419 35003
rect 22094 35000 22100 35012
rect 21407 34972 22100 35000
rect 21407 34969 21419 34972
rect 21361 34963 21419 34969
rect 22094 34960 22100 34972
rect 22152 35000 22158 35012
rect 22664 35000 22692 35031
rect 24854 35028 24860 35040
rect 24912 35028 24918 35080
rect 22152 34972 22692 35000
rect 25041 35003 25099 35009
rect 22152 34960 22158 34972
rect 25041 34969 25053 35003
rect 25087 35000 25099 35003
rect 26878 35000 26884 35012
rect 25087 34972 26884 35000
rect 25087 34969 25099 34972
rect 25041 34963 25099 34969
rect 26878 34960 26884 34972
rect 26936 34960 26942 35012
rect 1486 34932 1492 34944
rect 1447 34904 1492 34932
rect 1486 34892 1492 34904
rect 1544 34892 1550 34944
rect 22830 34932 22836 34944
rect 22791 34904 22836 34932
rect 22830 34892 22836 34904
rect 22888 34892 22894 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 23201 34731 23259 34737
rect 6886 34700 22876 34728
rect 1949 34595 2007 34601
rect 1949 34561 1961 34595
rect 1995 34592 2007 34595
rect 6886 34592 6914 34700
rect 22370 34660 22376 34672
rect 22331 34632 22376 34660
rect 22370 34620 22376 34632
rect 22428 34620 22434 34672
rect 22848 34660 22876 34700
rect 23201 34697 23213 34731
rect 23247 34728 23259 34731
rect 23750 34728 23756 34740
rect 23247 34700 23756 34728
rect 23247 34697 23259 34700
rect 23201 34691 23259 34697
rect 23750 34688 23756 34700
rect 23808 34688 23814 34740
rect 27430 34688 27436 34740
rect 27488 34728 27494 34740
rect 27525 34731 27583 34737
rect 27525 34728 27537 34731
rect 27488 34700 27537 34728
rect 27488 34688 27494 34700
rect 27525 34697 27537 34700
rect 27571 34697 27583 34731
rect 27525 34691 27583 34697
rect 36906 34688 36912 34740
rect 36964 34728 36970 34740
rect 37921 34731 37979 34737
rect 37921 34728 37933 34731
rect 36964 34700 37933 34728
rect 36964 34688 36970 34700
rect 37921 34697 37933 34700
rect 37967 34697 37979 34731
rect 37921 34691 37979 34697
rect 23658 34660 23664 34672
rect 22848 34632 23664 34660
rect 23658 34620 23664 34632
rect 23716 34620 23722 34672
rect 22189 34595 22247 34601
rect 22189 34592 22201 34595
rect 1995 34564 6914 34592
rect 12406 34564 22201 34592
rect 1995 34561 2007 34564
rect 1949 34555 2007 34561
rect 2222 34524 2228 34536
rect 2183 34496 2228 34524
rect 2222 34484 2228 34496
rect 2280 34524 2286 34536
rect 2685 34527 2743 34533
rect 2685 34524 2697 34527
rect 2280 34496 2697 34524
rect 2280 34484 2286 34496
rect 2685 34493 2697 34496
rect 2731 34493 2743 34527
rect 2685 34487 2743 34493
rect 4798 34484 4804 34536
rect 4856 34524 4862 34536
rect 12406 34524 12434 34564
rect 22189 34561 22201 34564
rect 22235 34561 22247 34595
rect 27338 34592 27344 34604
rect 27299 34564 27344 34592
rect 22189 34555 22247 34561
rect 27338 34552 27344 34564
rect 27396 34552 27402 34604
rect 37461 34595 37519 34601
rect 37461 34561 37473 34595
rect 37507 34592 37519 34595
rect 38102 34592 38108 34604
rect 37507 34564 38108 34592
rect 37507 34561 37519 34564
rect 37461 34555 37519 34561
rect 38102 34552 38108 34564
rect 38160 34552 38166 34604
rect 4856 34496 12434 34524
rect 4856 34484 4862 34496
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 2314 34184 2320 34196
rect 2275 34156 2320 34184
rect 2314 34144 2320 34156
rect 2372 34144 2378 34196
rect 22373 34187 22431 34193
rect 22373 34153 22385 34187
rect 22419 34184 22431 34187
rect 22646 34184 22652 34196
rect 22419 34156 22652 34184
rect 22419 34153 22431 34156
rect 22373 34147 22431 34153
rect 22646 34144 22652 34156
rect 22704 34144 22710 34196
rect 27338 34184 27344 34196
rect 27299 34156 27344 34184
rect 27338 34144 27344 34156
rect 27396 34144 27402 34196
rect 22738 34076 22744 34128
rect 22796 34116 22802 34128
rect 23201 34119 23259 34125
rect 23201 34116 23213 34119
rect 22796 34088 23213 34116
rect 22796 34076 22802 34088
rect 23201 34085 23213 34088
rect 23247 34116 23259 34119
rect 23247 34088 35894 34116
rect 23247 34085 23259 34088
rect 23201 34079 23259 34085
rect 1673 34051 1731 34057
rect 1673 34017 1685 34051
rect 1719 34048 1731 34051
rect 21818 34048 21824 34060
rect 1719 34020 2912 34048
rect 21779 34020 21824 34048
rect 1719 34017 1731 34020
rect 1673 34011 1731 34017
rect 1762 33940 1768 33992
rect 1820 33980 1826 33992
rect 1949 33983 2007 33989
rect 1949 33980 1961 33983
rect 1820 33952 1961 33980
rect 1820 33940 1826 33952
rect 1949 33949 1961 33952
rect 1995 33949 2007 33983
rect 1949 33943 2007 33949
rect 1670 33804 1676 33856
rect 1728 33844 1734 33856
rect 2884 33853 2912 34020
rect 21818 34008 21824 34020
rect 21876 34008 21882 34060
rect 26697 34051 26755 34057
rect 26697 34048 26709 34051
rect 25516 34020 26709 34048
rect 21542 33980 21548 33992
rect 21503 33952 21548 33980
rect 21542 33940 21548 33952
rect 21600 33940 21606 33992
rect 22278 33940 22284 33992
rect 22336 33980 22342 33992
rect 22557 33983 22615 33989
rect 22557 33980 22569 33983
rect 22336 33952 22569 33980
rect 22336 33940 22342 33952
rect 22557 33949 22569 33952
rect 22603 33949 22615 33983
rect 22557 33943 22615 33949
rect 1857 33847 1915 33853
rect 1857 33844 1869 33847
rect 1728 33816 1869 33844
rect 1728 33804 1734 33816
rect 1857 33813 1869 33816
rect 1903 33813 1915 33847
rect 1857 33807 1915 33813
rect 2869 33847 2927 33853
rect 2869 33813 2881 33847
rect 2915 33844 2927 33847
rect 4614 33844 4620 33856
rect 2915 33816 4620 33844
rect 2915 33813 2927 33816
rect 2869 33807 2927 33813
rect 4614 33804 4620 33816
rect 4672 33804 4678 33856
rect 23750 33804 23756 33856
rect 23808 33844 23814 33856
rect 25516 33853 25544 34020
rect 26697 34017 26709 34020
rect 26743 34017 26755 34051
rect 26697 34011 26755 34017
rect 35866 33980 35894 34088
rect 37826 33980 37832 33992
rect 35866 33952 37832 33980
rect 37826 33940 37832 33952
rect 37884 33940 37890 33992
rect 26881 33915 26939 33921
rect 26881 33881 26893 33915
rect 26927 33912 26939 33915
rect 36906 33912 36912 33924
rect 26927 33884 31754 33912
rect 26927 33881 26939 33884
rect 26881 33875 26939 33881
rect 25501 33847 25559 33853
rect 25501 33844 25513 33847
rect 23808 33816 25513 33844
rect 23808 33804 23814 33816
rect 25501 33813 25513 33816
rect 25547 33813 25559 33847
rect 26142 33844 26148 33856
rect 26103 33816 26148 33844
rect 25501 33807 25559 33813
rect 26142 33804 26148 33816
rect 26200 33844 26206 33856
rect 26973 33847 27031 33853
rect 26973 33844 26985 33847
rect 26200 33816 26985 33844
rect 26200 33804 26206 33816
rect 26973 33813 26985 33816
rect 27019 33813 27031 33847
rect 31726 33844 31754 33884
rect 35866 33884 36912 33912
rect 35866 33844 35894 33884
rect 36906 33872 36912 33884
rect 36964 33872 36970 33924
rect 31726 33816 35894 33844
rect 26973 33807 27031 33813
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 1581 33643 1639 33649
rect 1581 33609 1593 33643
rect 1627 33640 1639 33643
rect 5445 33643 5503 33649
rect 5445 33640 5457 33643
rect 1627 33612 5457 33640
rect 1627 33609 1639 33612
rect 1581 33603 1639 33609
rect 5445 33609 5457 33612
rect 5491 33609 5503 33643
rect 17862 33640 17868 33652
rect 17823 33612 17868 33640
rect 5445 33603 5503 33609
rect 17862 33600 17868 33612
rect 17920 33600 17926 33652
rect 22278 33640 22284 33652
rect 22239 33612 22284 33640
rect 22278 33600 22284 33612
rect 22336 33600 22342 33652
rect 22738 33640 22744 33652
rect 22699 33612 22744 33640
rect 22738 33600 22744 33612
rect 22796 33600 22802 33652
rect 23290 33572 23296 33584
rect 12406 33544 23296 33572
rect 1394 33504 1400 33516
rect 1355 33476 1400 33504
rect 1394 33464 1400 33476
rect 1452 33504 1458 33516
rect 2041 33507 2099 33513
rect 2041 33504 2053 33507
rect 1452 33476 2053 33504
rect 1452 33464 1458 33476
rect 2041 33473 2053 33476
rect 2087 33473 2099 33507
rect 2041 33467 2099 33473
rect 5537 33507 5595 33513
rect 5537 33473 5549 33507
rect 5583 33504 5595 33507
rect 6365 33507 6423 33513
rect 6365 33504 6377 33507
rect 5583 33476 6377 33504
rect 5583 33473 5595 33476
rect 5537 33467 5595 33473
rect 6365 33473 6377 33476
rect 6411 33504 6423 33507
rect 12406 33504 12434 33544
rect 23290 33532 23296 33544
rect 23348 33532 23354 33584
rect 6411 33476 12434 33504
rect 6411 33473 6423 33476
rect 6365 33467 6423 33473
rect 17126 33464 17132 33516
rect 17184 33504 17190 33516
rect 17773 33507 17831 33513
rect 17773 33504 17785 33507
rect 17184 33476 17785 33504
rect 17184 33464 17190 33476
rect 17773 33473 17785 33476
rect 17819 33473 17831 33507
rect 22649 33507 22707 33513
rect 22649 33504 22661 33507
rect 17773 33467 17831 33473
rect 22066 33476 22661 33504
rect 5442 33396 5448 33448
rect 5500 33436 5506 33448
rect 5629 33439 5687 33445
rect 5629 33436 5641 33439
rect 5500 33408 5641 33436
rect 5500 33396 5506 33408
rect 5629 33405 5641 33408
rect 5675 33405 5687 33439
rect 5629 33399 5687 33405
rect 17037 33439 17095 33445
rect 17037 33405 17049 33439
rect 17083 33436 17095 33439
rect 17681 33439 17739 33445
rect 17681 33436 17693 33439
rect 17083 33408 17693 33436
rect 17083 33405 17095 33408
rect 17037 33399 17095 33405
rect 17681 33405 17693 33408
rect 17727 33436 17739 33439
rect 20254 33436 20260 33448
rect 17727 33408 20260 33436
rect 17727 33405 17739 33408
rect 17681 33399 17739 33405
rect 20254 33396 20260 33408
rect 20312 33396 20318 33448
rect 15102 33328 15108 33380
rect 15160 33368 15166 33380
rect 21177 33371 21235 33377
rect 21177 33368 21189 33371
rect 15160 33340 21189 33368
rect 15160 33328 15166 33340
rect 21177 33337 21189 33340
rect 21223 33368 21235 33371
rect 22066 33368 22094 33476
rect 22649 33473 22661 33476
rect 22695 33473 22707 33507
rect 22649 33467 22707 33473
rect 37461 33507 37519 33513
rect 37461 33473 37473 33507
rect 37507 33504 37519 33507
rect 38102 33504 38108 33516
rect 37507 33476 38108 33504
rect 37507 33473 37519 33476
rect 37461 33467 37519 33473
rect 38102 33464 38108 33476
rect 38160 33464 38166 33516
rect 22925 33439 22983 33445
rect 22925 33405 22937 33439
rect 22971 33436 22983 33439
rect 23477 33439 23535 33445
rect 23477 33436 23489 33439
rect 22971 33408 23489 33436
rect 22971 33405 22983 33408
rect 22925 33399 22983 33405
rect 23477 33405 23489 33408
rect 23523 33405 23535 33439
rect 23477 33399 23535 33405
rect 21223 33340 22094 33368
rect 21223 33337 21235 33340
rect 21177 33331 21235 33337
rect 5077 33303 5135 33309
rect 5077 33269 5089 33303
rect 5123 33300 5135 33303
rect 5166 33300 5172 33312
rect 5123 33272 5172 33300
rect 5123 33269 5135 33272
rect 5077 33263 5135 33269
rect 5166 33260 5172 33272
rect 5224 33260 5230 33312
rect 18230 33300 18236 33312
rect 18191 33272 18236 33300
rect 18230 33260 18236 33272
rect 18288 33260 18294 33312
rect 20254 33260 20260 33312
rect 20312 33300 20318 33312
rect 22940 33300 22968 33399
rect 23290 33328 23296 33380
rect 23348 33368 23354 33380
rect 37921 33371 37979 33377
rect 37921 33368 37933 33371
rect 23348 33340 37933 33368
rect 23348 33328 23354 33340
rect 37921 33337 37933 33340
rect 37967 33337 37979 33371
rect 37921 33331 37979 33337
rect 20312 33272 22968 33300
rect 20312 33260 20318 33272
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 5442 33056 5448 33108
rect 5500 33096 5506 33108
rect 5905 33099 5963 33105
rect 5905 33096 5917 33099
rect 5500 33068 5917 33096
rect 5500 33056 5506 33068
rect 5905 33065 5917 33068
rect 5951 33065 5963 33099
rect 17126 33096 17132 33108
rect 17087 33068 17132 33096
rect 5905 33059 5963 33065
rect 17126 33056 17132 33068
rect 17184 33056 17190 33108
rect 22189 33099 22247 33105
rect 22189 33065 22201 33099
rect 22235 33096 22247 33099
rect 27614 33096 27620 33108
rect 22235 33068 27620 33096
rect 22235 33065 22247 33068
rect 22189 33059 22247 33065
rect 27614 33056 27620 33068
rect 27672 33056 27678 33108
rect 29733 33099 29791 33105
rect 29733 33065 29745 33099
rect 29779 33096 29791 33099
rect 35986 33096 35992 33108
rect 29779 33068 35992 33096
rect 29779 33065 29791 33068
rect 29733 33059 29791 33065
rect 35986 33056 35992 33068
rect 36044 33056 36050 33108
rect 23017 33031 23075 33037
rect 23017 32997 23029 33031
rect 23063 33028 23075 33031
rect 23382 33028 23388 33040
rect 23063 33000 23388 33028
rect 23063 32997 23075 33000
rect 23017 32991 23075 32997
rect 23382 32988 23388 33000
rect 23440 32988 23446 33040
rect 22649 32963 22707 32969
rect 22649 32929 22661 32963
rect 22695 32960 22707 32963
rect 22830 32960 22836 32972
rect 22695 32932 22836 32960
rect 22695 32929 22707 32932
rect 22649 32923 22707 32929
rect 22830 32920 22836 32932
rect 22888 32920 22894 32972
rect 1394 32892 1400 32904
rect 1355 32864 1400 32892
rect 1394 32852 1400 32864
rect 1452 32892 1458 32904
rect 2041 32895 2099 32901
rect 2041 32892 2053 32895
rect 1452 32864 2053 32892
rect 1452 32852 1458 32864
rect 2041 32861 2053 32864
rect 2087 32861 2099 32895
rect 2041 32855 2099 32861
rect 22005 32895 22063 32901
rect 22005 32861 22017 32895
rect 22051 32892 22063 32895
rect 22554 32892 22560 32904
rect 22051 32864 22560 32892
rect 22051 32861 22063 32864
rect 22005 32855 22063 32861
rect 22554 32852 22560 32864
rect 22612 32852 22618 32904
rect 29362 32852 29368 32904
rect 29420 32892 29426 32904
rect 29549 32895 29607 32901
rect 29549 32892 29561 32895
rect 29420 32864 29561 32892
rect 29420 32852 29426 32864
rect 29549 32861 29561 32864
rect 29595 32861 29607 32895
rect 29549 32855 29607 32861
rect 37461 32895 37519 32901
rect 37461 32861 37473 32895
rect 37507 32892 37519 32895
rect 38102 32892 38108 32904
rect 37507 32864 38108 32892
rect 37507 32861 37519 32864
rect 37461 32855 37519 32861
rect 38102 32852 38108 32864
rect 38160 32852 38166 32904
rect 15102 32824 15108 32836
rect 1596 32796 15108 32824
rect 1596 32765 1624 32796
rect 15102 32784 15108 32796
rect 15160 32784 15166 32836
rect 21726 32784 21732 32836
rect 21784 32824 21790 32836
rect 23569 32827 23627 32833
rect 23569 32824 23581 32827
rect 21784 32796 23581 32824
rect 21784 32784 21790 32796
rect 23569 32793 23581 32796
rect 23615 32824 23627 32827
rect 23750 32824 23756 32836
rect 23615 32796 23756 32824
rect 23615 32793 23627 32796
rect 23569 32787 23627 32793
rect 23750 32784 23756 32796
rect 23808 32784 23814 32836
rect 1581 32759 1639 32765
rect 1581 32725 1593 32759
rect 1627 32725 1639 32759
rect 1581 32719 1639 32725
rect 20714 32716 20720 32768
rect 20772 32756 20778 32768
rect 21269 32759 21327 32765
rect 21269 32756 21281 32759
rect 20772 32728 21281 32756
rect 20772 32716 20778 32728
rect 21269 32725 21281 32728
rect 21315 32725 21327 32759
rect 21269 32719 21327 32725
rect 22646 32716 22652 32768
rect 22704 32756 22710 32768
rect 23109 32759 23167 32765
rect 23109 32756 23121 32759
rect 22704 32728 23121 32756
rect 22704 32716 22710 32728
rect 23109 32725 23121 32728
rect 23155 32725 23167 32759
rect 23109 32719 23167 32725
rect 36538 32716 36544 32768
rect 36596 32756 36602 32768
rect 37921 32759 37979 32765
rect 37921 32756 37933 32759
rect 36596 32728 37933 32756
rect 36596 32716 36602 32728
rect 37921 32725 37933 32728
rect 37967 32725 37979 32759
rect 37921 32719 37979 32725
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 19242 32512 19248 32564
rect 19300 32552 19306 32564
rect 20073 32555 20131 32561
rect 20073 32552 20085 32555
rect 19300 32524 20085 32552
rect 19300 32512 19306 32524
rect 20073 32521 20085 32524
rect 20119 32521 20131 32555
rect 20073 32515 20131 32521
rect 20990 32512 20996 32564
rect 21048 32552 21054 32564
rect 21910 32552 21916 32564
rect 21048 32524 21916 32552
rect 21048 32512 21054 32524
rect 21910 32512 21916 32524
rect 21968 32552 21974 32564
rect 22189 32555 22247 32561
rect 22189 32552 22201 32555
rect 21968 32524 22201 32552
rect 21968 32512 21974 32524
rect 22189 32521 22201 32524
rect 22235 32521 22247 32555
rect 22554 32552 22560 32564
rect 22515 32524 22560 32552
rect 22189 32515 22247 32521
rect 22554 32512 22560 32524
rect 22612 32512 22618 32564
rect 23661 32555 23719 32561
rect 23661 32521 23673 32555
rect 23707 32552 23719 32555
rect 24489 32555 24547 32561
rect 24489 32552 24501 32555
rect 23707 32524 24501 32552
rect 23707 32521 23719 32524
rect 23661 32515 23719 32521
rect 24489 32521 24501 32524
rect 24535 32552 24547 32555
rect 27062 32552 27068 32564
rect 24535 32524 27068 32552
rect 24535 32521 24547 32524
rect 24489 32515 24547 32521
rect 27062 32512 27068 32524
rect 27120 32512 27126 32564
rect 29362 32552 29368 32564
rect 29323 32524 29368 32552
rect 29362 32512 29368 32524
rect 29420 32512 29426 32564
rect 37921 32555 37979 32561
rect 37921 32552 37933 32555
rect 35866 32524 37933 32552
rect 20714 32444 20720 32496
rect 20772 32484 20778 32496
rect 22097 32487 22155 32493
rect 22097 32484 22109 32487
rect 20772 32456 22109 32484
rect 20772 32444 20778 32456
rect 22097 32453 22109 32456
rect 22143 32453 22155 32487
rect 23566 32484 23572 32496
rect 23479 32456 23572 32484
rect 22097 32447 22155 32453
rect 23566 32444 23572 32456
rect 23624 32484 23630 32496
rect 35866 32484 35894 32524
rect 37921 32521 37933 32524
rect 37967 32521 37979 32555
rect 37921 32515 37979 32521
rect 23624 32456 35894 32484
rect 23624 32444 23630 32456
rect 1673 32419 1731 32425
rect 1673 32385 1685 32419
rect 1719 32416 1731 32419
rect 2682 32416 2688 32428
rect 1719 32388 2688 32416
rect 1719 32385 1731 32388
rect 1673 32379 1731 32385
rect 2682 32376 2688 32388
rect 2740 32376 2746 32428
rect 21085 32419 21143 32425
rect 21085 32385 21097 32419
rect 21131 32416 21143 32419
rect 21358 32416 21364 32428
rect 21131 32388 21364 32416
rect 21131 32385 21143 32388
rect 21085 32379 21143 32385
rect 21358 32376 21364 32388
rect 21416 32376 21422 32428
rect 28997 32419 29055 32425
rect 28997 32416 29009 32419
rect 28092 32388 29009 32416
rect 21726 32308 21732 32360
rect 21784 32348 21790 32360
rect 21913 32351 21971 32357
rect 21913 32348 21925 32351
rect 21784 32320 21925 32348
rect 21784 32308 21790 32320
rect 21913 32317 21925 32320
rect 21959 32317 21971 32351
rect 23750 32348 23756 32360
rect 23711 32320 23756 32348
rect 21913 32311 21971 32317
rect 23750 32308 23756 32320
rect 23808 32308 23814 32360
rect 21269 32283 21327 32289
rect 21269 32249 21281 32283
rect 21315 32280 21327 32283
rect 21315 32252 23796 32280
rect 21315 32249 21327 32252
rect 21269 32243 21327 32249
rect 1486 32212 1492 32224
rect 1447 32184 1492 32212
rect 1486 32172 1492 32184
rect 1544 32172 1550 32224
rect 23198 32212 23204 32224
rect 23159 32184 23204 32212
rect 23198 32172 23204 32184
rect 23256 32172 23262 32224
rect 23768 32212 23796 32252
rect 23842 32240 23848 32292
rect 23900 32280 23906 32292
rect 28092 32289 28120 32388
rect 28997 32385 29009 32388
rect 29043 32385 29055 32419
rect 28997 32379 29055 32385
rect 37461 32419 37519 32425
rect 37461 32385 37473 32419
rect 37507 32416 37519 32419
rect 38102 32416 38108 32428
rect 37507 32388 38108 32416
rect 37507 32385 37519 32388
rect 37461 32379 37519 32385
rect 38102 32376 38108 32388
rect 38160 32376 38166 32428
rect 28718 32348 28724 32360
rect 28679 32320 28724 32348
rect 28718 32308 28724 32320
rect 28776 32308 28782 32360
rect 28905 32351 28963 32357
rect 28905 32317 28917 32351
rect 28951 32348 28963 32351
rect 29822 32348 29828 32360
rect 28951 32320 29828 32348
rect 28951 32317 28963 32320
rect 28905 32311 28963 32317
rect 29822 32308 29828 32320
rect 29880 32308 29886 32360
rect 28077 32283 28135 32289
rect 28077 32280 28089 32283
rect 23900 32252 28089 32280
rect 23900 32240 23906 32252
rect 28077 32249 28089 32252
rect 28123 32249 28135 32283
rect 28077 32243 28135 32249
rect 27890 32212 27896 32224
rect 23768 32184 27896 32212
rect 27890 32172 27896 32184
rect 27948 32172 27954 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 2682 32008 2688 32020
rect 2643 31980 2688 32008
rect 2682 31968 2688 31980
rect 2740 31968 2746 32020
rect 21358 32008 21364 32020
rect 6886 31980 21220 32008
rect 21319 31980 21364 32008
rect 5534 31900 5540 31952
rect 5592 31940 5598 31952
rect 6886 31940 6914 31980
rect 5592 31912 6914 31940
rect 5592 31900 5598 31912
rect 15010 31900 15016 31952
rect 15068 31940 15074 31952
rect 15657 31943 15715 31949
rect 15657 31940 15669 31943
rect 15068 31912 15669 31940
rect 15068 31900 15074 31912
rect 15657 31909 15669 31912
rect 15703 31940 15715 31943
rect 17313 31943 17371 31949
rect 17313 31940 17325 31943
rect 15703 31912 17325 31940
rect 15703 31909 15715 31912
rect 15657 31903 15715 31909
rect 1673 31875 1731 31881
rect 1673 31841 1685 31875
rect 1719 31872 1731 31875
rect 4062 31872 4068 31884
rect 1719 31844 4068 31872
rect 1719 31841 1731 31844
rect 1673 31835 1731 31841
rect 4062 31832 4068 31844
rect 4120 31832 4126 31884
rect 1394 31804 1400 31816
rect 1355 31776 1400 31804
rect 1394 31764 1400 31776
rect 1452 31764 1458 31816
rect 2866 31804 2872 31816
rect 2827 31776 2872 31804
rect 2866 31764 2872 31776
rect 2924 31764 2930 31816
rect 15028 31813 15056 31900
rect 15013 31807 15071 31813
rect 15013 31773 15025 31807
rect 15059 31773 15071 31807
rect 15013 31767 15071 31773
rect 15105 31807 15163 31813
rect 15105 31773 15117 31807
rect 15151 31804 15163 31807
rect 15286 31804 15292 31816
rect 15151 31776 15292 31804
rect 15151 31773 15163 31776
rect 15105 31767 15163 31773
rect 15286 31764 15292 31776
rect 15344 31764 15350 31816
rect 16868 31813 16896 31912
rect 17313 31909 17325 31912
rect 17359 31909 17371 31943
rect 17313 31903 17371 31909
rect 19242 31900 19248 31952
rect 19300 31940 19306 31952
rect 19300 31912 20944 31940
rect 19300 31900 19306 31912
rect 17865 31875 17923 31881
rect 17865 31841 17877 31875
rect 17911 31872 17923 31875
rect 18230 31872 18236 31884
rect 17911 31844 18236 31872
rect 17911 31841 17923 31844
rect 17865 31835 17923 31841
rect 18230 31832 18236 31844
rect 18288 31832 18294 31884
rect 20162 31872 20168 31884
rect 20075 31844 20168 31872
rect 20162 31832 20168 31844
rect 20220 31872 20226 31884
rect 20916 31881 20944 31912
rect 20717 31875 20775 31881
rect 20717 31872 20729 31875
rect 20220 31844 20729 31872
rect 20220 31832 20226 31844
rect 20717 31841 20729 31844
rect 20763 31841 20775 31875
rect 20717 31835 20775 31841
rect 20901 31875 20959 31881
rect 20901 31841 20913 31875
rect 20947 31841 20959 31875
rect 20901 31835 20959 31841
rect 16853 31807 16911 31813
rect 16853 31773 16865 31807
rect 16899 31773 16911 31807
rect 16853 31767 16911 31773
rect 18141 31807 18199 31813
rect 18141 31773 18153 31807
rect 18187 31804 18199 31807
rect 20990 31804 20996 31816
rect 18187 31776 20996 31804
rect 18187 31773 18199 31776
rect 18141 31767 18199 31773
rect 20990 31764 20996 31776
rect 21048 31764 21054 31816
rect 21192 31736 21220 31980
rect 21358 31968 21364 31980
rect 21416 31968 21422 32020
rect 21910 32008 21916 32020
rect 21823 31980 21916 32008
rect 21910 31968 21916 31980
rect 21968 32008 21974 32020
rect 23106 32008 23112 32020
rect 21968 31980 23112 32008
rect 21968 31968 21974 31980
rect 23106 31968 23112 31980
rect 23164 31968 23170 32020
rect 23382 32008 23388 32020
rect 23343 31980 23388 32008
rect 23382 31968 23388 31980
rect 23440 31968 23446 32020
rect 22480 31912 22968 31940
rect 21634 31832 21640 31884
rect 21692 31872 21698 31884
rect 21692 31844 22048 31872
rect 21692 31832 21698 31844
rect 22020 31816 22048 31844
rect 22002 31764 22008 31816
rect 22060 31804 22066 31816
rect 22480 31804 22508 31912
rect 22060 31776 22508 31804
rect 22741 31807 22799 31813
rect 22060 31764 22066 31776
rect 22741 31773 22753 31807
rect 22787 31773 22799 31807
rect 22940 31804 22968 31912
rect 23106 31872 23112 31884
rect 23067 31844 23112 31872
rect 23106 31832 23112 31844
rect 23164 31832 23170 31884
rect 23226 31875 23284 31881
rect 23226 31841 23238 31875
rect 23272 31872 23284 31875
rect 23566 31872 23572 31884
rect 23272 31844 23572 31872
rect 23272 31841 23284 31844
rect 23226 31835 23284 31841
rect 23566 31832 23572 31844
rect 23624 31832 23630 31884
rect 37829 31875 37887 31881
rect 37829 31841 37841 31875
rect 37875 31872 37887 31875
rect 38378 31872 38384 31884
rect 37875 31844 38384 31872
rect 37875 31841 37887 31844
rect 37829 31835 37887 31841
rect 38378 31832 38384 31844
rect 38436 31832 38442 31884
rect 28445 31807 28503 31813
rect 28445 31804 28457 31807
rect 22940 31776 28457 31804
rect 22741 31767 22799 31773
rect 28445 31773 28457 31776
rect 28491 31804 28503 31807
rect 28718 31804 28724 31816
rect 28491 31776 28724 31804
rect 28491 31773 28503 31776
rect 28445 31767 28503 31773
rect 22756 31736 22784 31767
rect 28718 31764 28724 31776
rect 28776 31764 28782 31816
rect 37369 31807 37427 31813
rect 37369 31773 37381 31807
rect 37415 31804 37427 31807
rect 38010 31804 38016 31816
rect 37415 31776 38016 31804
rect 37415 31773 37427 31776
rect 37369 31767 37427 31773
rect 38010 31764 38016 31776
rect 38068 31764 38074 31816
rect 21192 31708 22784 31736
rect 16758 31668 16764 31680
rect 16719 31640 16764 31668
rect 16758 31628 16764 31640
rect 16816 31628 16822 31680
rect 20990 31668 20996 31680
rect 20951 31640 20996 31668
rect 20990 31628 20996 31640
rect 21048 31628 21054 31680
rect 22756 31668 22784 31708
rect 23017 31739 23075 31745
rect 23017 31705 23029 31739
rect 23063 31736 23075 31739
rect 23063 31708 24348 31736
rect 23063 31705 23075 31708
rect 23017 31699 23075 31705
rect 24320 31680 24348 31708
rect 23842 31668 23848 31680
rect 22756 31640 23848 31668
rect 23842 31628 23848 31640
rect 23900 31628 23906 31680
rect 24302 31628 24308 31680
rect 24360 31668 24366 31680
rect 24397 31671 24455 31677
rect 24397 31668 24409 31671
rect 24360 31640 24409 31668
rect 24360 31628 24366 31640
rect 24397 31637 24409 31640
rect 24443 31637 24455 31671
rect 24397 31631 24455 31637
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 2317 31467 2375 31473
rect 2317 31433 2329 31467
rect 2363 31464 2375 31467
rect 2866 31464 2872 31476
rect 2363 31436 2872 31464
rect 2363 31433 2375 31436
rect 2317 31427 2375 31433
rect 2866 31424 2872 31436
rect 2924 31424 2930 31476
rect 3970 31424 3976 31476
rect 4028 31464 4034 31476
rect 20257 31467 20315 31473
rect 20257 31464 20269 31467
rect 4028 31436 20269 31464
rect 4028 31424 4034 31436
rect 20257 31433 20269 31436
rect 20303 31464 20315 31467
rect 20990 31464 20996 31476
rect 20303 31436 20996 31464
rect 20303 31433 20315 31436
rect 20257 31427 20315 31433
rect 20990 31424 20996 31436
rect 21048 31424 21054 31476
rect 21726 31424 21732 31476
rect 21784 31464 21790 31476
rect 21821 31467 21879 31473
rect 21821 31464 21833 31467
rect 21784 31436 21833 31464
rect 21784 31424 21790 31436
rect 21821 31433 21833 31436
rect 21867 31433 21879 31467
rect 21821 31427 21879 31433
rect 23106 31424 23112 31476
rect 23164 31464 23170 31476
rect 23293 31467 23351 31473
rect 23293 31464 23305 31467
rect 23164 31436 23305 31464
rect 23164 31424 23170 31436
rect 23293 31433 23305 31436
rect 23339 31433 23351 31467
rect 23842 31464 23848 31476
rect 23803 31436 23848 31464
rect 23293 31427 23351 31433
rect 23842 31424 23848 31436
rect 23900 31424 23906 31476
rect 1949 31399 2007 31405
rect 1949 31365 1961 31399
rect 1995 31396 2007 31399
rect 2590 31396 2596 31408
rect 1995 31368 2596 31396
rect 1995 31365 2007 31368
rect 1949 31359 2007 31365
rect 2590 31356 2596 31368
rect 2648 31356 2654 31408
rect 2777 31399 2835 31405
rect 2777 31365 2789 31399
rect 2823 31396 2835 31399
rect 5442 31396 5448 31408
rect 2823 31368 5448 31396
rect 2823 31365 2835 31368
rect 2777 31359 2835 31365
rect 2792 31328 2820 31359
rect 5442 31356 5448 31368
rect 5500 31356 5506 31408
rect 15286 31356 15292 31408
rect 15344 31356 15350 31408
rect 22741 31399 22799 31405
rect 22741 31365 22753 31399
rect 22787 31396 22799 31399
rect 23198 31396 23204 31408
rect 22787 31368 23204 31396
rect 22787 31365 22799 31368
rect 22741 31359 22799 31365
rect 23198 31356 23204 31368
rect 23256 31356 23262 31408
rect 5166 31328 5172 31340
rect 1688 31300 2820 31328
rect 5127 31300 5172 31328
rect 1688 31269 1716 31300
rect 5166 31288 5172 31300
rect 5224 31288 5230 31340
rect 14185 31331 14243 31337
rect 14185 31297 14197 31331
rect 14231 31328 14243 31331
rect 14274 31328 14280 31340
rect 14231 31300 14280 31328
rect 14231 31297 14243 31300
rect 14185 31291 14243 31297
rect 14274 31288 14280 31300
rect 14332 31288 14338 31340
rect 20806 31288 20812 31340
rect 20864 31328 20870 31340
rect 22922 31328 22928 31340
rect 20864 31300 22928 31328
rect 20864 31288 20870 31300
rect 22922 31288 22928 31300
rect 22980 31288 22986 31340
rect 1673 31263 1731 31269
rect 1673 31229 1685 31263
rect 1719 31229 1731 31263
rect 1854 31260 1860 31272
rect 1815 31232 1860 31260
rect 1673 31223 1731 31229
rect 1854 31220 1860 31232
rect 1912 31220 1918 31272
rect 14550 31260 14556 31272
rect 14511 31232 14556 31260
rect 14550 31220 14556 31232
rect 14608 31220 14614 31272
rect 15979 31263 16037 31269
rect 15979 31229 15991 31263
rect 16025 31260 16037 31263
rect 17221 31263 17279 31269
rect 17221 31260 17233 31263
rect 16025 31232 17233 31260
rect 16025 31229 16037 31232
rect 15979 31223 16037 31229
rect 17221 31229 17233 31232
rect 17267 31229 17279 31263
rect 17221 31223 17279 31229
rect 18046 31220 18052 31272
rect 18104 31260 18110 31272
rect 22557 31263 22615 31269
rect 22557 31260 22569 31263
rect 18104 31232 22569 31260
rect 18104 31220 18110 31232
rect 22557 31229 22569 31232
rect 22603 31229 22615 31263
rect 22557 31223 22615 31229
rect 20898 31152 20904 31204
rect 20956 31192 20962 31204
rect 37366 31192 37372 31204
rect 20956 31164 37372 31192
rect 20956 31152 20962 31164
rect 37366 31152 37372 31164
rect 37424 31152 37430 31204
rect 1578 31084 1584 31136
rect 1636 31124 1642 31136
rect 1762 31124 1768 31136
rect 1636 31096 1768 31124
rect 1636 31084 1642 31096
rect 1762 31084 1768 31096
rect 1820 31084 1826 31136
rect 4982 31124 4988 31136
rect 4943 31096 4988 31124
rect 4982 31084 4988 31096
rect 5040 31084 5046 31136
rect 15746 31084 15752 31136
rect 15804 31124 15810 31136
rect 16669 31127 16727 31133
rect 16669 31124 16681 31127
rect 15804 31096 16681 31124
rect 15804 31084 15810 31096
rect 16669 31093 16681 31096
rect 16715 31093 16727 31127
rect 16669 31087 16727 31093
rect 18230 31084 18236 31136
rect 18288 31124 18294 31136
rect 21726 31124 21732 31136
rect 18288 31096 21732 31124
rect 18288 31084 18294 31096
rect 21726 31084 21732 31096
rect 21784 31084 21790 31136
rect 24486 31124 24492 31136
rect 24399 31096 24492 31124
rect 24486 31084 24492 31096
rect 24544 31124 24550 31136
rect 37458 31124 37464 31136
rect 24544 31096 37464 31124
rect 24544 31084 24550 31096
rect 37458 31084 37464 31096
rect 37516 31084 37522 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 1394 30920 1400 30932
rect 1355 30892 1400 30920
rect 1394 30880 1400 30892
rect 1452 30880 1458 30932
rect 14550 30920 14556 30932
rect 14511 30892 14556 30920
rect 14550 30880 14556 30892
rect 14608 30880 14614 30932
rect 17218 30861 17224 30864
rect 17175 30855 17224 30861
rect 17175 30821 17187 30855
rect 17221 30821 17224 30855
rect 17175 30815 17224 30821
rect 17218 30812 17224 30815
rect 17276 30812 17282 30864
rect 24486 30852 24492 30864
rect 23492 30824 24492 30852
rect 14274 30744 14280 30796
rect 14332 30784 14338 30796
rect 15381 30787 15439 30793
rect 15381 30784 15393 30787
rect 14332 30756 15393 30784
rect 14332 30744 14338 30756
rect 15381 30753 15393 30756
rect 15427 30753 15439 30787
rect 15746 30784 15752 30796
rect 15707 30756 15752 30784
rect 15381 30747 15439 30753
rect 15746 30744 15752 30756
rect 15804 30744 15810 30796
rect 23492 30793 23520 30824
rect 24486 30812 24492 30824
rect 24544 30812 24550 30864
rect 23477 30787 23535 30793
rect 23477 30753 23489 30787
rect 23523 30753 23535 30787
rect 23477 30747 23535 30753
rect 23569 30787 23627 30793
rect 23569 30753 23581 30787
rect 23615 30753 23627 30787
rect 23569 30747 23627 30753
rect 23584 30716 23612 30747
rect 22480 30688 23612 30716
rect 16758 30608 16764 30660
rect 16816 30608 16822 30660
rect 22480 30592 22508 30688
rect 22462 30580 22468 30592
rect 22423 30552 22468 30580
rect 22462 30540 22468 30552
rect 22520 30540 22526 30592
rect 23014 30580 23020 30592
rect 22975 30552 23020 30580
rect 23014 30540 23020 30552
rect 23072 30540 23078 30592
rect 23385 30583 23443 30589
rect 23385 30549 23397 30583
rect 23431 30580 23443 30583
rect 24302 30580 24308 30592
rect 23431 30552 24308 30580
rect 23431 30549 23443 30552
rect 23385 30543 23443 30549
rect 24302 30540 24308 30552
rect 24360 30580 24366 30592
rect 24397 30583 24455 30589
rect 24397 30580 24409 30583
rect 24360 30552 24409 30580
rect 24360 30540 24366 30552
rect 24397 30549 24409 30552
rect 24443 30549 24455 30583
rect 24397 30543 24455 30549
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 22557 30311 22615 30317
rect 22557 30277 22569 30311
rect 22603 30308 22615 30311
rect 23014 30308 23020 30320
rect 22603 30280 23020 30308
rect 22603 30277 22615 30280
rect 22557 30271 22615 30277
rect 23014 30268 23020 30280
rect 23072 30268 23078 30320
rect 23658 30268 23664 30320
rect 23716 30308 23722 30320
rect 24305 30311 24363 30317
rect 24305 30308 24317 30311
rect 23716 30280 24317 30308
rect 23716 30268 23722 30280
rect 24305 30277 24317 30280
rect 24351 30277 24363 30311
rect 24305 30271 24363 30277
rect 1673 30243 1731 30249
rect 1673 30209 1685 30243
rect 1719 30240 1731 30243
rect 2225 30243 2283 30249
rect 2225 30240 2237 30243
rect 1719 30212 2237 30240
rect 1719 30209 1731 30212
rect 1673 30203 1731 30209
rect 2225 30209 2237 30212
rect 2271 30240 2283 30243
rect 17218 30240 17224 30252
rect 2271 30212 17224 30240
rect 2271 30209 2283 30212
rect 2225 30203 2283 30209
rect 17218 30200 17224 30212
rect 17276 30200 17282 30252
rect 23385 30243 23443 30249
rect 23385 30209 23397 30243
rect 23431 30240 23443 30243
rect 24397 30243 24455 30249
rect 23431 30212 23980 30240
rect 23431 30209 23443 30212
rect 23385 30203 23443 30209
rect 22738 30132 22744 30184
rect 22796 30172 22802 30184
rect 23014 30172 23020 30184
rect 22796 30144 23020 30172
rect 22796 30132 22802 30144
rect 23014 30132 23020 30144
rect 23072 30132 23078 30184
rect 21174 30064 21180 30116
rect 21232 30104 21238 30116
rect 23952 30113 23980 30212
rect 24397 30209 24409 30243
rect 24443 30240 24455 30243
rect 25133 30243 25191 30249
rect 25133 30240 25145 30243
rect 24443 30212 25145 30240
rect 24443 30209 24455 30212
rect 24397 30203 24455 30209
rect 25133 30209 25145 30212
rect 25179 30240 25191 30243
rect 27522 30240 27528 30252
rect 25179 30212 26234 30240
rect 27483 30212 27528 30240
rect 25179 30209 25191 30212
rect 25133 30203 25191 30209
rect 24581 30175 24639 30181
rect 24581 30141 24593 30175
rect 24627 30172 24639 30175
rect 24854 30172 24860 30184
rect 24627 30144 24860 30172
rect 24627 30141 24639 30144
rect 24581 30135 24639 30141
rect 24854 30132 24860 30144
rect 24912 30172 24918 30184
rect 24912 30144 25820 30172
rect 24912 30132 24918 30144
rect 22373 30107 22431 30113
rect 22373 30104 22385 30107
rect 21232 30076 22385 30104
rect 21232 30064 21238 30076
rect 22373 30073 22385 30076
rect 22419 30073 22431 30107
rect 22373 30067 22431 30073
rect 23937 30107 23995 30113
rect 23937 30073 23949 30107
rect 23983 30073 23995 30107
rect 23937 30067 23995 30073
rect 1486 30036 1492 30048
rect 1447 30008 1492 30036
rect 1486 29996 1492 30008
rect 1544 29996 1550 30048
rect 23293 30039 23351 30045
rect 23293 30005 23305 30039
rect 23339 30036 23351 30039
rect 23842 30036 23848 30048
rect 23339 30008 23848 30036
rect 23339 30005 23351 30008
rect 23293 29999 23351 30005
rect 23842 29996 23848 30008
rect 23900 29996 23906 30048
rect 25792 30045 25820 30144
rect 26206 30104 26234 30212
rect 27522 30200 27528 30212
rect 27580 30200 27586 30252
rect 30374 30200 30380 30252
rect 30432 30240 30438 30252
rect 37829 30243 37887 30249
rect 37829 30240 37841 30243
rect 30432 30212 37841 30240
rect 30432 30200 30438 30212
rect 37829 30209 37841 30212
rect 37875 30209 37887 30243
rect 37829 30203 37887 30209
rect 37918 30104 37924 30116
rect 26206 30076 37924 30104
rect 37918 30064 37924 30076
rect 37976 30064 37982 30116
rect 25777 30039 25835 30045
rect 25777 30005 25789 30039
rect 25823 30036 25835 30039
rect 26050 30036 26056 30048
rect 25823 30008 26056 30036
rect 25823 30005 25835 30008
rect 25777 29999 25835 30005
rect 26050 29996 26056 30008
rect 26108 29996 26114 30048
rect 26970 30036 26976 30048
rect 26931 30008 26976 30036
rect 26970 29996 26976 30008
rect 27028 29996 27034 30048
rect 27709 30039 27767 30045
rect 27709 30005 27721 30039
rect 27755 30036 27767 30039
rect 30926 30036 30932 30048
rect 27755 30008 30932 30036
rect 27755 30005 27767 30008
rect 27709 29999 27767 30005
rect 30926 29996 30932 30008
rect 30984 29996 30990 30048
rect 38010 30036 38016 30048
rect 37971 30008 38016 30036
rect 38010 29996 38016 30008
rect 38068 29996 38074 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 20625 29835 20683 29841
rect 20625 29801 20637 29835
rect 20671 29832 20683 29835
rect 21082 29832 21088 29844
rect 20671 29804 21088 29832
rect 20671 29801 20683 29804
rect 20625 29795 20683 29801
rect 21082 29792 21088 29804
rect 21140 29792 21146 29844
rect 23382 29832 23388 29844
rect 21192 29804 23388 29832
rect 16942 29724 16948 29776
rect 17000 29764 17006 29776
rect 21192 29764 21220 29804
rect 23382 29792 23388 29804
rect 23440 29792 23446 29844
rect 23658 29792 23664 29844
rect 23716 29832 23722 29844
rect 23753 29835 23811 29841
rect 23753 29832 23765 29835
rect 23716 29804 23765 29832
rect 23716 29792 23722 29804
rect 23753 29801 23765 29804
rect 23799 29801 23811 29835
rect 27522 29832 27528 29844
rect 27483 29804 27528 29832
rect 23753 29795 23811 29801
rect 27522 29792 27528 29804
rect 27580 29792 27586 29844
rect 34606 29792 34612 29844
rect 34664 29832 34670 29844
rect 34885 29835 34943 29841
rect 34885 29832 34897 29835
rect 34664 29804 34897 29832
rect 34664 29792 34670 29804
rect 34885 29801 34897 29804
rect 34931 29801 34943 29835
rect 34885 29795 34943 29801
rect 22186 29764 22192 29776
rect 17000 29736 21220 29764
rect 22112 29736 22192 29764
rect 17000 29724 17006 29736
rect 22112 29705 22140 29736
rect 22186 29724 22192 29736
rect 22244 29724 22250 29776
rect 22278 29724 22284 29776
rect 22336 29764 22342 29776
rect 23106 29764 23112 29776
rect 22336 29736 23112 29764
rect 22336 29724 22342 29736
rect 23106 29724 23112 29736
rect 23164 29724 23170 29776
rect 22097 29699 22155 29705
rect 22097 29665 22109 29699
rect 22143 29665 22155 29699
rect 26970 29696 26976 29708
rect 22097 29659 22155 29665
rect 22848 29668 26976 29696
rect 1673 29631 1731 29637
rect 1673 29597 1685 29631
rect 1719 29628 1731 29631
rect 4982 29628 4988 29640
rect 1719 29600 4988 29628
rect 1719 29597 1731 29600
rect 1673 29591 1731 29597
rect 4982 29588 4988 29600
rect 5040 29588 5046 29640
rect 20438 29628 20444 29640
rect 20399 29600 20444 29628
rect 20438 29588 20444 29600
rect 20496 29588 20502 29640
rect 22186 29588 22192 29640
rect 22244 29628 22250 29640
rect 22373 29631 22431 29637
rect 22373 29628 22385 29631
rect 22244 29600 22385 29628
rect 22244 29588 22250 29600
rect 22373 29597 22385 29600
rect 22419 29597 22431 29631
rect 22373 29591 22431 29597
rect 9030 29520 9036 29572
rect 9088 29560 9094 29572
rect 20530 29560 20536 29572
rect 9088 29532 20536 29560
rect 9088 29520 9094 29532
rect 20530 29520 20536 29532
rect 20588 29520 20594 29572
rect 1486 29492 1492 29504
rect 1447 29464 1492 29492
rect 1486 29452 1492 29464
rect 1544 29452 1550 29504
rect 22554 29452 22560 29504
rect 22612 29492 22618 29504
rect 22848 29501 22876 29668
rect 26970 29656 26976 29668
rect 27028 29656 27034 29708
rect 36722 29696 36728 29708
rect 31036 29668 36728 29696
rect 23842 29588 23848 29640
rect 23900 29628 23906 29640
rect 31036 29628 31064 29668
rect 36722 29656 36728 29668
rect 36780 29656 36786 29708
rect 23900 29600 31064 29628
rect 23900 29588 23906 29600
rect 34238 29588 34244 29640
rect 34296 29628 34302 29640
rect 34701 29631 34759 29637
rect 34701 29628 34713 29631
rect 34296 29600 34713 29628
rect 34296 29588 34302 29600
rect 34701 29597 34713 29600
rect 34747 29597 34759 29631
rect 34701 29591 34759 29597
rect 37461 29631 37519 29637
rect 37461 29597 37473 29631
rect 37507 29628 37519 29631
rect 38102 29628 38108 29640
rect 37507 29600 38108 29628
rect 37507 29597 37519 29600
rect 37461 29591 37519 29597
rect 38102 29588 38108 29600
rect 38160 29588 38166 29640
rect 23106 29520 23112 29572
rect 23164 29520 23170 29572
rect 24762 29520 24768 29572
rect 24820 29560 24826 29572
rect 25501 29563 25559 29569
rect 24820 29532 24865 29560
rect 24820 29520 24826 29532
rect 25501 29529 25513 29563
rect 25547 29529 25559 29563
rect 25501 29523 25559 29529
rect 22833 29495 22891 29501
rect 22833 29492 22845 29495
rect 22612 29464 22845 29492
rect 22612 29452 22618 29464
rect 22833 29461 22845 29464
rect 22879 29461 22891 29495
rect 23124 29492 23152 29520
rect 25516 29492 25544 29523
rect 23124 29464 25544 29492
rect 22833 29455 22891 29461
rect 26050 29452 26056 29504
rect 26108 29492 26114 29504
rect 26145 29495 26203 29501
rect 26145 29492 26157 29495
rect 26108 29464 26157 29492
rect 26108 29452 26114 29464
rect 26145 29461 26157 29464
rect 26191 29461 26203 29495
rect 27062 29492 27068 29504
rect 27023 29464 27068 29492
rect 26145 29455 26203 29461
rect 27062 29452 27068 29464
rect 27120 29452 27126 29504
rect 27157 29495 27215 29501
rect 27157 29461 27169 29495
rect 27203 29492 27215 29495
rect 27982 29492 27988 29504
rect 27203 29464 27988 29492
rect 27203 29461 27215 29464
rect 27157 29455 27215 29461
rect 27982 29452 27988 29464
rect 28040 29452 28046 29504
rect 37918 29492 37924 29504
rect 37879 29464 37924 29492
rect 37918 29452 37924 29464
rect 37976 29452 37982 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 19334 29288 19340 29300
rect 2746 29260 19340 29288
rect 1394 29152 1400 29164
rect 1355 29124 1400 29152
rect 1394 29112 1400 29124
rect 1452 29152 1458 29164
rect 2041 29155 2099 29161
rect 2041 29152 2053 29155
rect 1452 29124 2053 29152
rect 1452 29112 1458 29124
rect 2041 29121 2053 29124
rect 2087 29121 2099 29155
rect 2041 29115 2099 29121
rect 1581 29019 1639 29025
rect 1581 28985 1593 29019
rect 1627 29016 1639 29019
rect 2746 29016 2774 29260
rect 19334 29248 19340 29260
rect 19392 29248 19398 29300
rect 19797 29291 19855 29297
rect 19797 29257 19809 29291
rect 19843 29288 19855 29291
rect 20346 29288 20352 29300
rect 19843 29260 20352 29288
rect 19843 29257 19855 29260
rect 19797 29251 19855 29257
rect 20346 29248 20352 29260
rect 20404 29248 20410 29300
rect 22186 29288 22192 29300
rect 22147 29260 22192 29288
rect 22186 29248 22192 29260
rect 22244 29248 22250 29300
rect 23290 29288 23296 29300
rect 22480 29260 23296 29288
rect 22480 29232 22508 29260
rect 23290 29248 23296 29260
rect 23348 29248 23354 29300
rect 23382 29248 23388 29300
rect 23440 29288 23446 29300
rect 27062 29288 27068 29300
rect 23440 29260 27068 29288
rect 23440 29248 23446 29260
rect 27062 29248 27068 29260
rect 27120 29248 27126 29300
rect 34238 29288 34244 29300
rect 34199 29260 34244 29288
rect 34238 29248 34244 29260
rect 34296 29248 34302 29300
rect 15194 29180 15200 29232
rect 15252 29220 15258 29232
rect 16025 29223 16083 29229
rect 16025 29220 16037 29223
rect 15252 29192 16037 29220
rect 15252 29180 15258 29192
rect 16025 29189 16037 29192
rect 16071 29220 16083 29223
rect 22462 29220 22468 29232
rect 16071 29192 22468 29220
rect 16071 29189 16083 29192
rect 16025 29183 16083 29189
rect 22462 29180 22468 29192
rect 22520 29180 22526 29232
rect 22649 29223 22707 29229
rect 22649 29189 22661 29223
rect 22695 29220 22707 29223
rect 24029 29223 24087 29229
rect 24029 29220 24041 29223
rect 22695 29192 24041 29220
rect 22695 29189 22707 29192
rect 22649 29183 22707 29189
rect 24029 29189 24041 29192
rect 24075 29220 24087 29223
rect 33873 29223 33931 29229
rect 24075 29192 26234 29220
rect 24075 29189 24087 29192
rect 24029 29183 24087 29189
rect 15473 29155 15531 29161
rect 15473 29121 15485 29155
rect 15519 29121 15531 29155
rect 15473 29115 15531 29121
rect 20257 29155 20315 29161
rect 20257 29121 20269 29155
rect 20303 29152 20315 29155
rect 20806 29152 20812 29164
rect 20303 29124 20812 29152
rect 20303 29121 20315 29124
rect 20257 29115 20315 29121
rect 4614 29044 4620 29096
rect 4672 29084 4678 29096
rect 5258 29084 5264 29096
rect 4672 29056 5264 29084
rect 4672 29044 4678 29056
rect 5258 29044 5264 29056
rect 5316 29084 5322 29096
rect 15488 29084 15516 29115
rect 20806 29112 20812 29124
rect 20864 29112 20870 29164
rect 22557 29155 22615 29161
rect 22557 29121 22569 29155
rect 22603 29152 22615 29155
rect 26206 29152 26234 29192
rect 33873 29189 33885 29223
rect 33919 29220 33931 29223
rect 37918 29220 37924 29232
rect 33919 29192 37924 29220
rect 33919 29189 33931 29192
rect 33873 29183 33931 29189
rect 37918 29180 37924 29192
rect 37976 29180 37982 29232
rect 37461 29155 37519 29161
rect 22603 29124 23244 29152
rect 26206 29124 35894 29152
rect 22603 29121 22615 29124
rect 22557 29115 22615 29121
rect 16669 29087 16727 29093
rect 16669 29084 16681 29087
rect 5316 29056 16681 29084
rect 5316 29044 5322 29056
rect 16669 29053 16681 29056
rect 16715 29084 16727 29087
rect 18598 29084 18604 29096
rect 16715 29056 18604 29084
rect 16715 29053 16727 29056
rect 16669 29047 16727 29053
rect 18598 29044 18604 29056
rect 18656 29044 18662 29096
rect 20530 29084 20536 29096
rect 20491 29056 20536 29084
rect 20530 29044 20536 29056
rect 20588 29044 20594 29096
rect 22741 29087 22799 29093
rect 22741 29053 22753 29087
rect 22787 29053 22799 29087
rect 22741 29047 22799 29053
rect 1627 28988 2774 29016
rect 1627 28985 1639 28988
rect 1581 28979 1639 28985
rect 22554 28976 22560 29028
rect 22612 29016 22618 29028
rect 22756 29016 22784 29047
rect 23216 29028 23244 29124
rect 23290 29044 23296 29096
rect 23348 29084 23354 29096
rect 26970 29084 26976 29096
rect 23348 29056 26976 29084
rect 23348 29044 23354 29056
rect 26970 29044 26976 29056
rect 27028 29044 27034 29096
rect 33594 29084 33600 29096
rect 33555 29056 33600 29084
rect 33594 29044 33600 29056
rect 33652 29044 33658 29096
rect 33781 29087 33839 29093
rect 33781 29053 33793 29087
rect 33827 29053 33839 29087
rect 35866 29084 35894 29124
rect 37461 29121 37473 29155
rect 37507 29152 37519 29155
rect 38102 29152 38108 29164
rect 37507 29124 38108 29152
rect 37507 29121 37519 29124
rect 37461 29115 37519 29121
rect 38102 29112 38108 29124
rect 38160 29112 38166 29164
rect 37550 29084 37556 29096
rect 35866 29056 37556 29084
rect 33781 29047 33839 29053
rect 22612 28988 22784 29016
rect 22612 28976 22618 28988
rect 23198 28976 23204 29028
rect 23256 29016 23262 29028
rect 23385 29019 23443 29025
rect 23385 29016 23397 29019
rect 23256 28988 23397 29016
rect 23256 28976 23262 28988
rect 23385 28985 23397 28988
rect 23431 28985 23443 29019
rect 32950 29016 32956 29028
rect 32911 28988 32956 29016
rect 23385 28979 23443 28985
rect 32950 28976 32956 28988
rect 33008 29016 33014 29028
rect 33796 29016 33824 29047
rect 37550 29044 37556 29056
rect 37608 29044 37614 29096
rect 33008 28988 33824 29016
rect 33008 28976 33014 28988
rect 36630 28976 36636 29028
rect 36688 29016 36694 29028
rect 37921 29019 37979 29025
rect 37921 29016 37933 29019
rect 36688 28988 37933 29016
rect 36688 28976 36694 28988
rect 37921 28985 37933 28988
rect 37967 28985 37979 29019
rect 37921 28979 37979 28985
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 20806 28744 20812 28756
rect 20767 28716 20812 28744
rect 20806 28704 20812 28716
rect 20864 28704 20870 28756
rect 33410 28744 33416 28756
rect 33323 28716 33416 28744
rect 33410 28704 33416 28716
rect 33468 28744 33474 28756
rect 33594 28744 33600 28756
rect 33468 28716 33600 28744
rect 33468 28704 33474 28716
rect 33594 28704 33600 28716
rect 33652 28704 33658 28756
rect 4706 28636 4712 28688
rect 4764 28676 4770 28688
rect 25958 28676 25964 28688
rect 4764 28648 25964 28676
rect 4764 28636 4770 28648
rect 25958 28636 25964 28648
rect 26016 28636 26022 28688
rect 19426 28568 19432 28620
rect 19484 28608 19490 28620
rect 20162 28608 20168 28620
rect 19484 28580 20168 28608
rect 19484 28568 19490 28580
rect 20162 28568 20168 28580
rect 20220 28608 20226 28620
rect 21361 28611 21419 28617
rect 21361 28608 21373 28611
rect 20220 28580 21373 28608
rect 20220 28568 20226 28580
rect 21361 28577 21373 28580
rect 21407 28608 21419 28611
rect 22462 28608 22468 28620
rect 21407 28580 22468 28608
rect 21407 28577 21419 28580
rect 21361 28571 21419 28577
rect 22462 28568 22468 28580
rect 22520 28568 22526 28620
rect 3234 28500 3240 28552
rect 3292 28540 3298 28552
rect 22005 28543 22063 28549
rect 22005 28540 22017 28543
rect 3292 28512 22017 28540
rect 3292 28500 3298 28512
rect 22005 28509 22017 28512
rect 22051 28509 22063 28543
rect 22005 28503 22063 28509
rect 20346 28432 20352 28484
rect 20404 28472 20410 28484
rect 21177 28475 21235 28481
rect 21177 28472 21189 28475
rect 20404 28444 21189 28472
rect 20404 28432 20410 28444
rect 21177 28441 21189 28444
rect 21223 28441 21235 28475
rect 21177 28435 21235 28441
rect 21910 28432 21916 28484
rect 21968 28472 21974 28484
rect 22189 28475 22247 28481
rect 22189 28472 22201 28475
rect 21968 28444 22201 28472
rect 21968 28432 21974 28444
rect 22189 28441 22201 28444
rect 22235 28441 22247 28475
rect 22189 28435 22247 28441
rect 4614 28364 4620 28416
rect 4672 28404 4678 28416
rect 4985 28407 5043 28413
rect 4985 28404 4997 28407
rect 4672 28376 4997 28404
rect 4672 28364 4678 28376
rect 4985 28373 4997 28376
rect 5031 28373 5043 28407
rect 4985 28367 5043 28373
rect 19426 28364 19432 28416
rect 19484 28404 19490 28416
rect 19613 28407 19671 28413
rect 19613 28404 19625 28407
rect 19484 28376 19625 28404
rect 19484 28364 19490 28376
rect 19613 28373 19625 28376
rect 19659 28373 19671 28407
rect 20162 28404 20168 28416
rect 20123 28376 20168 28404
rect 19613 28367 19671 28373
rect 20162 28364 20168 28376
rect 20220 28364 20226 28416
rect 21269 28407 21327 28413
rect 21269 28373 21281 28407
rect 21315 28404 21327 28407
rect 22094 28404 22100 28416
rect 21315 28376 22100 28404
rect 21315 28373 21327 28376
rect 21269 28367 21327 28373
rect 22094 28364 22100 28376
rect 22152 28404 22158 28416
rect 22741 28407 22799 28413
rect 22741 28404 22753 28407
rect 22152 28376 22753 28404
rect 22152 28364 22158 28376
rect 22741 28373 22753 28376
rect 22787 28373 22799 28407
rect 22741 28367 22799 28373
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 1581 28203 1639 28209
rect 1581 28169 1593 28203
rect 1627 28200 1639 28203
rect 4433 28203 4491 28209
rect 4433 28200 4445 28203
rect 1627 28172 4445 28200
rect 1627 28169 1639 28172
rect 1581 28163 1639 28169
rect 4433 28169 4445 28172
rect 4479 28169 4491 28203
rect 4433 28163 4491 28169
rect 4525 28203 4583 28209
rect 4525 28169 4537 28203
rect 4571 28200 4583 28203
rect 5350 28200 5356 28212
rect 4571 28172 5356 28200
rect 4571 28169 4583 28172
rect 4525 28163 4583 28169
rect 5350 28160 5356 28172
rect 5408 28160 5414 28212
rect 19334 28200 19340 28212
rect 19295 28172 19340 28200
rect 19334 28160 19340 28172
rect 19392 28160 19398 28212
rect 20349 28203 20407 28209
rect 20349 28169 20361 28203
rect 20395 28200 20407 28203
rect 20438 28200 20444 28212
rect 20395 28172 20444 28200
rect 20395 28169 20407 28172
rect 20349 28163 20407 28169
rect 20438 28160 20444 28172
rect 20496 28160 20502 28212
rect 21910 28200 21916 28212
rect 21871 28172 21916 28200
rect 21910 28160 21916 28172
rect 21968 28160 21974 28212
rect 22281 28203 22339 28209
rect 22281 28169 22293 28203
rect 22327 28200 22339 28203
rect 23106 28200 23112 28212
rect 22327 28172 23112 28200
rect 22327 28169 22339 28172
rect 22281 28163 22339 28169
rect 23106 28160 23112 28172
rect 23164 28160 23170 28212
rect 19352 28132 19380 28160
rect 20717 28135 20775 28141
rect 20717 28132 20729 28135
rect 19352 28104 20729 28132
rect 20717 28101 20729 28104
rect 20763 28101 20775 28135
rect 20717 28095 20775 28101
rect 22002 28092 22008 28144
rect 22060 28132 22066 28144
rect 22060 28104 35894 28132
rect 22060 28092 22066 28104
rect 1394 28064 1400 28076
rect 1355 28036 1400 28064
rect 1394 28024 1400 28036
rect 1452 28064 1458 28076
rect 2041 28067 2099 28073
rect 2041 28064 2053 28067
rect 1452 28036 2053 28064
rect 1452 28024 1458 28036
rect 2041 28033 2053 28036
rect 2087 28033 2099 28067
rect 2041 28027 2099 28033
rect 19889 28067 19947 28073
rect 19889 28033 19901 28067
rect 19935 28064 19947 28067
rect 20809 28067 20867 28073
rect 20809 28064 20821 28067
rect 19935 28036 20821 28064
rect 19935 28033 19947 28036
rect 19889 28027 19947 28033
rect 20809 28033 20821 28036
rect 20855 28064 20867 28067
rect 21266 28064 21272 28076
rect 20855 28036 21272 28064
rect 20855 28033 20867 28036
rect 20809 28027 20867 28033
rect 21266 28024 21272 28036
rect 21324 28024 21330 28076
rect 25314 28064 25320 28076
rect 22066 28036 25320 28064
rect 4341 27999 4399 28005
rect 4341 27965 4353 27999
rect 4387 27996 4399 27999
rect 4614 27996 4620 28008
rect 4387 27968 4620 27996
rect 4387 27965 4399 27968
rect 4341 27959 4399 27965
rect 4614 27956 4620 27968
rect 4672 27956 4678 28008
rect 20162 27956 20168 28008
rect 20220 27996 20226 28008
rect 20901 27999 20959 28005
rect 20901 27996 20913 27999
rect 20220 27968 20913 27996
rect 20220 27956 20226 27968
rect 20901 27965 20913 27968
rect 20947 27996 20959 27999
rect 22066 27996 22094 28036
rect 25314 28024 25320 28036
rect 25372 28024 25378 28076
rect 25593 28067 25651 28073
rect 25593 28033 25605 28067
rect 25639 28064 25651 28067
rect 26050 28064 26056 28076
rect 25639 28036 26056 28064
rect 25639 28033 25651 28036
rect 25593 28027 25651 28033
rect 26050 28024 26056 28036
rect 26108 28064 26114 28076
rect 26108 28036 27108 28064
rect 26108 28024 26114 28036
rect 20947 27968 22094 27996
rect 22373 27999 22431 28005
rect 20947 27965 20959 27968
rect 20901 27959 20959 27965
rect 22373 27965 22385 27999
rect 22419 27965 22431 27999
rect 22373 27959 22431 27965
rect 22388 27928 22416 27959
rect 22462 27956 22468 28008
rect 22520 27996 22526 28008
rect 23109 27999 23167 28005
rect 23109 27996 23121 27999
rect 22520 27968 23121 27996
rect 22520 27956 22526 27968
rect 23109 27965 23121 27968
rect 23155 27965 23167 27999
rect 25958 27996 25964 28008
rect 25919 27968 25964 27996
rect 23109 27959 23167 27965
rect 25958 27956 25964 27968
rect 26016 27956 26022 28008
rect 22388 27900 23520 27928
rect 23492 27872 23520 27900
rect 4890 27860 4896 27872
rect 4851 27832 4896 27860
rect 4890 27820 4896 27832
rect 4948 27820 4954 27872
rect 23474 27820 23480 27872
rect 23532 27860 23538 27872
rect 23661 27863 23719 27869
rect 23661 27860 23673 27863
rect 23532 27832 23673 27860
rect 23532 27820 23538 27832
rect 23661 27829 23673 27832
rect 23707 27829 23719 27863
rect 25976 27860 26004 27956
rect 26142 27860 26148 27872
rect 25976 27832 26148 27860
rect 23661 27823 23719 27829
rect 26142 27820 26148 27832
rect 26200 27820 26206 27872
rect 27080 27869 27108 28036
rect 35866 27928 35894 28104
rect 37829 28067 37887 28073
rect 37829 28064 37841 28067
rect 37292 28036 37841 28064
rect 37292 27937 37320 28036
rect 37829 28033 37841 28036
rect 37875 28033 37887 28067
rect 37829 28027 37887 28033
rect 37277 27931 37335 27937
rect 37277 27928 37289 27931
rect 35866 27900 37289 27928
rect 37277 27897 37289 27900
rect 37323 27897 37335 27931
rect 38010 27928 38016 27940
rect 37971 27900 38016 27928
rect 37277 27891 37335 27897
rect 38010 27888 38016 27900
rect 38068 27888 38074 27940
rect 27065 27863 27123 27869
rect 27065 27829 27077 27863
rect 27111 27860 27123 27863
rect 37550 27860 37556 27872
rect 27111 27832 37556 27860
rect 27111 27829 27123 27832
rect 27065 27823 27123 27829
rect 37550 27820 37556 27832
rect 37608 27820 37614 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 20346 27616 20352 27668
rect 20404 27656 20410 27668
rect 21453 27659 21511 27665
rect 21453 27656 21465 27659
rect 20404 27628 21465 27656
rect 20404 27616 20410 27628
rect 21453 27625 21465 27628
rect 21499 27656 21511 27659
rect 23017 27659 23075 27665
rect 21499 27628 22416 27656
rect 21499 27625 21511 27628
rect 21453 27619 21511 27625
rect 1581 27591 1639 27597
rect 1581 27557 1593 27591
rect 1627 27588 1639 27591
rect 1854 27588 1860 27600
rect 1627 27560 1860 27588
rect 1627 27557 1639 27560
rect 1581 27551 1639 27557
rect 1854 27548 1860 27560
rect 1912 27548 1918 27600
rect 20990 27588 20996 27600
rect 20951 27560 20996 27588
rect 20990 27548 20996 27560
rect 21048 27588 21054 27600
rect 22388 27597 22416 27628
rect 23017 27625 23029 27659
rect 23063 27656 23075 27659
rect 23106 27656 23112 27668
rect 23063 27628 23112 27656
rect 23063 27625 23075 27628
rect 23017 27619 23075 27625
rect 23106 27616 23112 27628
rect 23164 27616 23170 27668
rect 22373 27591 22431 27597
rect 21048 27560 21588 27588
rect 21048 27548 21054 27560
rect 19426 27480 19432 27532
rect 19484 27520 19490 27532
rect 21560 27529 21588 27560
rect 22373 27557 22385 27591
rect 22419 27557 22431 27591
rect 22373 27551 22431 27557
rect 19797 27523 19855 27529
rect 19797 27520 19809 27523
rect 19484 27492 19809 27520
rect 19484 27480 19490 27492
rect 19797 27489 19809 27492
rect 19843 27489 19855 27523
rect 19797 27483 19855 27489
rect 21545 27523 21603 27529
rect 21545 27489 21557 27523
rect 21591 27489 21603 27523
rect 21545 27483 21603 27489
rect 1394 27452 1400 27464
rect 1355 27424 1400 27452
rect 1394 27412 1400 27424
rect 1452 27452 1458 27464
rect 2041 27455 2099 27461
rect 2041 27452 2053 27455
rect 1452 27424 2053 27452
rect 1452 27412 1458 27424
rect 2041 27421 2053 27424
rect 2087 27421 2099 27455
rect 2041 27415 2099 27421
rect 4890 27412 4896 27464
rect 4948 27452 4954 27464
rect 5261 27455 5319 27461
rect 5261 27452 5273 27455
rect 4948 27424 5273 27452
rect 4948 27412 4954 27424
rect 5261 27421 5273 27424
rect 5307 27421 5319 27455
rect 20898 27452 20904 27464
rect 5261 27415 5319 27421
rect 12406 27424 20904 27452
rect 5442 27384 5448 27396
rect 5403 27356 5448 27384
rect 5442 27344 5448 27356
rect 5500 27344 5506 27396
rect 3234 27276 3240 27328
rect 3292 27316 3298 27328
rect 12406 27316 12434 27424
rect 20898 27412 20904 27424
rect 20956 27452 20962 27464
rect 21453 27455 21511 27461
rect 21453 27452 21465 27455
rect 20956 27424 21465 27452
rect 20956 27412 20962 27424
rect 21453 27421 21465 27424
rect 21499 27421 21511 27455
rect 21453 27415 21511 27421
rect 21729 27455 21787 27461
rect 21729 27421 21741 27455
rect 21775 27452 21787 27455
rect 23106 27452 23112 27464
rect 21775 27424 23112 27452
rect 21775 27421 21787 27424
rect 21729 27415 21787 27421
rect 23106 27412 23112 27424
rect 23164 27412 23170 27464
rect 37829 27455 37887 27461
rect 37829 27452 37841 27455
rect 37292 27424 37841 27452
rect 17954 27344 17960 27396
rect 18012 27384 18018 27396
rect 18693 27387 18751 27393
rect 18693 27384 18705 27387
rect 18012 27356 18705 27384
rect 18012 27344 18018 27356
rect 18693 27353 18705 27356
rect 18739 27384 18751 27387
rect 20073 27387 20131 27393
rect 20073 27384 20085 27387
rect 18739 27356 20085 27384
rect 18739 27353 18751 27356
rect 18693 27347 18751 27353
rect 20073 27353 20085 27356
rect 20119 27353 20131 27387
rect 20073 27347 20131 27353
rect 37292 27328 37320 27424
rect 37829 27421 37841 27424
rect 37875 27421 37887 27455
rect 37829 27415 37887 27421
rect 19978 27316 19984 27328
rect 3292 27288 12434 27316
rect 19939 27288 19984 27316
rect 3292 27276 3298 27288
rect 19978 27276 19984 27288
rect 20036 27276 20042 27328
rect 20438 27316 20444 27328
rect 20399 27288 20444 27316
rect 20438 27276 20444 27288
rect 20496 27276 20502 27328
rect 21910 27316 21916 27328
rect 21871 27288 21916 27316
rect 21910 27276 21916 27288
rect 21968 27276 21974 27328
rect 37274 27316 37280 27328
rect 37235 27288 37280 27316
rect 37274 27276 37280 27288
rect 37332 27276 37338 27328
rect 38010 27316 38016 27328
rect 37971 27288 38016 27316
rect 38010 27276 38016 27288
rect 38068 27276 38074 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 14642 27072 14648 27124
rect 14700 27112 14706 27124
rect 18969 27115 19027 27121
rect 18969 27112 18981 27115
rect 14700 27084 18981 27112
rect 14700 27072 14706 27084
rect 18969 27081 18981 27084
rect 19015 27112 19027 27115
rect 19978 27112 19984 27124
rect 19015 27084 19984 27112
rect 19015 27081 19027 27084
rect 18969 27075 19027 27081
rect 19978 27072 19984 27084
rect 20036 27072 20042 27124
rect 22278 27112 22284 27124
rect 22066 27084 22284 27112
rect 5626 27004 5632 27056
rect 5684 27044 5690 27056
rect 21174 27044 21180 27056
rect 5684 27016 21180 27044
rect 5684 27004 5690 27016
rect 21174 27004 21180 27016
rect 21232 27004 21238 27056
rect 1673 26979 1731 26985
rect 1673 26945 1685 26979
rect 1719 26976 1731 26979
rect 2225 26979 2283 26985
rect 2225 26976 2237 26979
rect 1719 26948 2237 26976
rect 1719 26945 1731 26948
rect 1673 26939 1731 26945
rect 2225 26945 2237 26948
rect 2271 26976 2283 26979
rect 14826 26976 14832 26988
rect 2271 26948 14832 26976
rect 2271 26945 2283 26948
rect 2225 26939 2283 26945
rect 14826 26936 14832 26948
rect 14884 26936 14890 26988
rect 20073 26979 20131 26985
rect 20073 26945 20085 26979
rect 20119 26976 20131 26979
rect 20438 26976 20444 26988
rect 20119 26948 20444 26976
rect 20119 26945 20131 26948
rect 20073 26939 20131 26945
rect 20438 26936 20444 26948
rect 20496 26936 20502 26988
rect 20717 26979 20775 26985
rect 20717 26945 20729 26979
rect 20763 26976 20775 26979
rect 21821 26979 21879 26985
rect 21821 26976 21833 26979
rect 20763 26948 21833 26976
rect 20763 26945 20775 26948
rect 20717 26939 20775 26945
rect 21821 26945 21833 26948
rect 21867 26976 21879 26979
rect 22066 26976 22094 27084
rect 22278 27072 22284 27084
rect 22336 27072 22342 27124
rect 22465 27115 22523 27121
rect 22465 27081 22477 27115
rect 22511 27112 22523 27115
rect 23106 27112 23112 27124
rect 22511 27084 23112 27112
rect 22511 27081 22523 27084
rect 22465 27075 22523 27081
rect 23106 27072 23112 27084
rect 23164 27072 23170 27124
rect 21867 26948 22094 26976
rect 37461 26979 37519 26985
rect 21867 26945 21879 26948
rect 21821 26939 21879 26945
rect 37461 26945 37473 26979
rect 37507 26976 37519 26979
rect 38102 26976 38108 26988
rect 37507 26948 38108 26976
rect 37507 26945 37519 26948
rect 37461 26939 37519 26945
rect 4062 26868 4068 26920
rect 4120 26908 4126 26920
rect 6362 26908 6368 26920
rect 4120 26880 6368 26908
rect 4120 26868 4126 26880
rect 6362 26868 6368 26880
rect 6420 26868 6426 26920
rect 18598 26868 18604 26920
rect 18656 26908 18662 26920
rect 20732 26908 20760 26939
rect 38102 26936 38108 26948
rect 38160 26936 38166 26988
rect 20990 26908 20996 26920
rect 18656 26880 20760 26908
rect 20903 26880 20996 26908
rect 18656 26868 18662 26880
rect 20990 26868 20996 26880
rect 21048 26908 21054 26920
rect 21634 26908 21640 26920
rect 21048 26880 21640 26908
rect 21048 26868 21054 26880
rect 21634 26868 21640 26880
rect 21692 26868 21698 26920
rect 20257 26843 20315 26849
rect 20257 26809 20269 26843
rect 20303 26840 20315 26843
rect 20303 26812 26234 26840
rect 20303 26809 20315 26812
rect 20257 26803 20315 26809
rect 1486 26772 1492 26784
rect 1447 26744 1492 26772
rect 1486 26732 1492 26744
rect 1544 26732 1550 26784
rect 19426 26732 19432 26784
rect 19484 26772 19490 26784
rect 19521 26775 19579 26781
rect 19521 26772 19533 26775
rect 19484 26744 19533 26772
rect 19484 26732 19490 26744
rect 19521 26741 19533 26744
rect 19567 26741 19579 26775
rect 23198 26772 23204 26784
rect 23159 26744 23204 26772
rect 19521 26735 19579 26741
rect 23198 26732 23204 26744
rect 23256 26732 23262 26784
rect 26206 26772 26234 26812
rect 37274 26772 37280 26784
rect 26206 26744 37280 26772
rect 37274 26732 37280 26744
rect 37332 26732 37338 26784
rect 37918 26772 37924 26784
rect 37879 26744 37924 26772
rect 37918 26732 37924 26744
rect 37976 26732 37982 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 18598 26568 18604 26580
rect 18559 26540 18604 26568
rect 18598 26528 18604 26540
rect 18656 26528 18662 26580
rect 20898 26568 20904 26580
rect 20859 26540 20904 26568
rect 20898 26528 20904 26540
rect 20956 26568 20962 26580
rect 22741 26571 22799 26577
rect 20956 26540 22416 26568
rect 20956 26528 20962 26540
rect 21450 26460 21456 26512
rect 21508 26500 21514 26512
rect 22281 26503 22339 26509
rect 22281 26500 22293 26503
rect 21508 26472 22293 26500
rect 21508 26460 21514 26472
rect 22281 26469 22293 26472
rect 22327 26469 22339 26503
rect 22388 26500 22416 26540
rect 22741 26537 22753 26571
rect 22787 26568 22799 26571
rect 23382 26568 23388 26580
rect 22787 26540 23388 26568
rect 22787 26537 22799 26540
rect 22741 26531 22799 26537
rect 23382 26528 23388 26540
rect 23440 26528 23446 26580
rect 26418 26500 26424 26512
rect 22388 26472 26424 26500
rect 22281 26463 22339 26469
rect 26418 26460 26424 26472
rect 26476 26460 26482 26512
rect 38010 26500 38016 26512
rect 37971 26472 38016 26500
rect 38010 26460 38016 26472
rect 38068 26460 38074 26512
rect 23198 26392 23204 26444
rect 23256 26432 23262 26444
rect 37918 26432 37924 26444
rect 23256 26404 37924 26432
rect 23256 26392 23262 26404
rect 37918 26392 37924 26404
rect 37976 26392 37982 26444
rect 1673 26367 1731 26373
rect 1673 26333 1685 26367
rect 1719 26364 1731 26367
rect 3326 26364 3332 26376
rect 1719 26336 3332 26364
rect 1719 26333 1731 26336
rect 1673 26327 1731 26333
rect 3326 26324 3332 26336
rect 3384 26324 3390 26376
rect 21726 26324 21732 26376
rect 21784 26364 21790 26376
rect 21821 26367 21879 26373
rect 21821 26364 21833 26367
rect 21784 26336 21833 26364
rect 21784 26324 21790 26336
rect 21821 26333 21833 26336
rect 21867 26364 21879 26367
rect 22465 26367 22523 26373
rect 22465 26364 22477 26367
rect 21867 26336 22477 26364
rect 21867 26333 21879 26336
rect 21821 26327 21879 26333
rect 22465 26333 22477 26336
rect 22511 26333 22523 26367
rect 22465 26327 22523 26333
rect 22833 26367 22891 26373
rect 22833 26333 22845 26367
rect 22879 26364 22891 26367
rect 23216 26364 23244 26392
rect 22879 26336 23244 26364
rect 27249 26367 27307 26373
rect 22879 26333 22891 26336
rect 22833 26327 22891 26333
rect 27249 26333 27261 26367
rect 27295 26364 27307 26367
rect 27706 26364 27712 26376
rect 27295 26336 27712 26364
rect 27295 26333 27307 26336
rect 27249 26327 27307 26333
rect 27706 26324 27712 26336
rect 27764 26324 27770 26376
rect 37369 26367 37427 26373
rect 37369 26333 37381 26367
rect 37415 26364 37427 26367
rect 37829 26367 37887 26373
rect 37829 26364 37841 26367
rect 37415 26336 37841 26364
rect 37415 26333 37427 26336
rect 37369 26327 37427 26333
rect 37829 26333 37841 26336
rect 37875 26364 37887 26367
rect 38562 26364 38568 26376
rect 37875 26336 38568 26364
rect 37875 26333 37887 26336
rect 37829 26327 37887 26333
rect 38562 26324 38568 26336
rect 38620 26324 38626 26376
rect 30374 26296 30380 26308
rect 27448 26268 30380 26296
rect 1486 26228 1492 26240
rect 1447 26200 1492 26228
rect 1486 26188 1492 26200
rect 1544 26188 1550 26240
rect 23382 26228 23388 26240
rect 23343 26200 23388 26228
rect 23382 26188 23388 26200
rect 23440 26188 23446 26240
rect 27448 26237 27476 26268
rect 30374 26256 30380 26268
rect 30432 26256 30438 26308
rect 27433 26231 27491 26237
rect 27433 26197 27445 26231
rect 27479 26228 27491 26231
rect 27479 26200 27513 26228
rect 27479 26197 27491 26200
rect 27433 26191 27491 26197
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 18966 25984 18972 26036
rect 19024 26024 19030 26036
rect 19613 26027 19671 26033
rect 19613 26024 19625 26027
rect 19024 25996 19625 26024
rect 19024 25984 19030 25996
rect 19613 25993 19625 25996
rect 19659 25993 19671 26027
rect 19613 25987 19671 25993
rect 20901 26027 20959 26033
rect 20901 25993 20913 26027
rect 20947 26024 20959 26027
rect 20990 26024 20996 26036
rect 20947 25996 20996 26024
rect 20947 25993 20959 25996
rect 20901 25987 20959 25993
rect 20990 25984 20996 25996
rect 21048 25984 21054 26036
rect 23842 26024 23848 26036
rect 23803 25996 23848 26024
rect 23842 25984 23848 25996
rect 23900 25984 23906 26036
rect 26418 26024 26424 26036
rect 26379 25996 26424 26024
rect 26418 25984 26424 25996
rect 26476 26024 26482 26036
rect 27341 26027 27399 26033
rect 27341 26024 27353 26027
rect 26476 25996 27353 26024
rect 26476 25984 26482 25996
rect 27341 25993 27353 25996
rect 27387 25993 27399 26027
rect 27706 26024 27712 26036
rect 27667 25996 27712 26024
rect 27341 25987 27399 25993
rect 27706 25984 27712 25996
rect 27764 25984 27770 26036
rect 18138 25888 18144 25900
rect 18051 25860 18144 25888
rect 18138 25848 18144 25860
rect 18196 25888 18202 25900
rect 18598 25888 18604 25900
rect 18196 25860 18604 25888
rect 18196 25848 18202 25860
rect 18598 25848 18604 25860
rect 18656 25888 18662 25900
rect 19061 25891 19119 25897
rect 19061 25888 19073 25891
rect 18656 25860 19073 25888
rect 18656 25848 18662 25860
rect 19061 25857 19073 25860
rect 19107 25857 19119 25891
rect 19061 25851 19119 25857
rect 22370 25848 22376 25900
rect 22428 25888 22434 25900
rect 22649 25891 22707 25897
rect 22649 25888 22661 25891
rect 22428 25860 22661 25888
rect 22428 25848 22434 25860
rect 22649 25857 22661 25860
rect 22695 25857 22707 25891
rect 22649 25851 22707 25857
rect 22741 25891 22799 25897
rect 22741 25857 22753 25891
rect 22787 25888 22799 25891
rect 23860 25888 23888 25984
rect 22787 25860 23888 25888
rect 22787 25857 22799 25860
rect 22741 25851 22799 25857
rect 18417 25823 18475 25829
rect 18417 25789 18429 25823
rect 18463 25820 18475 25823
rect 19426 25820 19432 25832
rect 18463 25792 19432 25820
rect 18463 25789 18475 25792
rect 18417 25783 18475 25789
rect 19426 25780 19432 25792
rect 19484 25820 19490 25832
rect 20622 25820 20628 25832
rect 19484 25792 20628 25820
rect 19484 25780 19490 25792
rect 20622 25780 20628 25792
rect 20680 25780 20686 25832
rect 22462 25820 22468 25832
rect 22423 25792 22468 25820
rect 22462 25780 22468 25792
rect 22520 25780 22526 25832
rect 22554 25780 22560 25832
rect 22612 25820 22618 25832
rect 27062 25820 27068 25832
rect 22612 25792 22657 25820
rect 27023 25792 27068 25820
rect 22612 25780 22618 25792
rect 27062 25780 27068 25792
rect 27120 25780 27126 25832
rect 27249 25823 27307 25829
rect 27249 25789 27261 25823
rect 27295 25820 27307 25823
rect 37918 25820 37924 25832
rect 27295 25792 37924 25820
rect 27295 25789 27307 25792
rect 27249 25783 27307 25789
rect 37918 25780 37924 25792
rect 37976 25780 37982 25832
rect 21634 25712 21640 25764
rect 21692 25752 21698 25764
rect 23385 25755 23443 25761
rect 23385 25752 23397 25755
rect 21692 25724 23397 25752
rect 21692 25712 21698 25724
rect 23385 25721 23397 25724
rect 23431 25752 23443 25755
rect 36630 25752 36636 25764
rect 23431 25724 36636 25752
rect 23431 25721 23443 25724
rect 23385 25715 23443 25721
rect 36630 25712 36636 25724
rect 36688 25712 36694 25764
rect 1673 25687 1731 25693
rect 1673 25653 1685 25687
rect 1719 25684 1731 25687
rect 1854 25684 1860 25696
rect 1719 25656 1860 25684
rect 1719 25653 1731 25656
rect 1673 25647 1731 25653
rect 1854 25644 1860 25656
rect 1912 25644 1918 25696
rect 2314 25644 2320 25696
rect 2372 25684 2378 25696
rect 18046 25684 18052 25696
rect 2372 25656 18052 25684
rect 2372 25644 2378 25656
rect 18046 25644 18052 25656
rect 18104 25644 18110 25696
rect 20346 25684 20352 25696
rect 20307 25656 20352 25684
rect 20346 25644 20352 25656
rect 20404 25644 20410 25696
rect 22281 25687 22339 25693
rect 22281 25653 22293 25687
rect 22327 25684 22339 25687
rect 22646 25684 22652 25696
rect 22327 25656 22652 25684
rect 22327 25653 22339 25656
rect 22281 25647 22339 25653
rect 22646 25644 22652 25656
rect 22704 25644 22710 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 25314 25440 25320 25492
rect 25372 25480 25378 25492
rect 25501 25483 25559 25489
rect 25501 25480 25513 25483
rect 25372 25452 25513 25480
rect 25372 25440 25378 25452
rect 25501 25449 25513 25452
rect 25547 25449 25559 25483
rect 37918 25480 37924 25492
rect 37879 25452 37924 25480
rect 25501 25443 25559 25449
rect 37918 25440 37924 25452
rect 37976 25440 37982 25492
rect 20622 25372 20628 25424
rect 20680 25412 20686 25424
rect 20680 25384 21772 25412
rect 20680 25372 20686 25384
rect 18966 25304 18972 25356
rect 19024 25344 19030 25356
rect 19705 25347 19763 25353
rect 19705 25344 19717 25347
rect 19024 25316 19717 25344
rect 19024 25304 19030 25316
rect 19705 25313 19717 25316
rect 19751 25313 19763 25347
rect 19705 25307 19763 25313
rect 19889 25347 19947 25353
rect 19889 25313 19901 25347
rect 19935 25344 19947 25347
rect 20990 25344 20996 25356
rect 19935 25316 20996 25344
rect 19935 25313 19947 25316
rect 19889 25307 19947 25313
rect 20990 25304 20996 25316
rect 21048 25304 21054 25356
rect 21634 25344 21640 25356
rect 21595 25316 21640 25344
rect 21634 25304 21640 25316
rect 21692 25304 21698 25356
rect 21744 25353 21772 25384
rect 22278 25372 22284 25424
rect 22336 25412 22342 25424
rect 24394 25412 24400 25424
rect 22336 25384 24400 25412
rect 22336 25372 22342 25384
rect 24394 25372 24400 25384
rect 24452 25372 24458 25424
rect 21729 25347 21787 25353
rect 21729 25313 21741 25347
rect 21775 25313 21787 25347
rect 22922 25344 22928 25356
rect 22883 25316 22928 25344
rect 21729 25307 21787 25313
rect 22922 25304 22928 25316
rect 22980 25304 22986 25356
rect 1854 25276 1860 25288
rect 1815 25248 1860 25276
rect 1854 25236 1860 25248
rect 1912 25236 1918 25288
rect 17865 25279 17923 25285
rect 17865 25245 17877 25279
rect 17911 25276 17923 25279
rect 18138 25276 18144 25288
rect 17911 25248 18144 25276
rect 17911 25245 17923 25248
rect 17865 25239 17923 25245
rect 18138 25236 18144 25248
rect 18196 25236 18202 25288
rect 19613 25279 19671 25285
rect 19613 25245 19625 25279
rect 19659 25276 19671 25279
rect 20346 25276 20352 25288
rect 19659 25248 20352 25276
rect 19659 25245 19671 25248
rect 19613 25239 19671 25245
rect 20346 25236 20352 25248
rect 20404 25276 20410 25288
rect 23106 25276 23112 25288
rect 20404 25248 23112 25276
rect 20404 25236 20410 25248
rect 23106 25236 23112 25248
rect 23164 25236 23170 25288
rect 23201 25279 23259 25285
rect 23201 25245 23213 25279
rect 23247 25276 23259 25279
rect 23658 25276 23664 25288
rect 23247 25248 23664 25276
rect 23247 25245 23259 25248
rect 23201 25239 23259 25245
rect 23658 25236 23664 25248
rect 23716 25236 23722 25288
rect 23753 25279 23811 25285
rect 23753 25245 23765 25279
rect 23799 25276 23811 25279
rect 35434 25276 35440 25288
rect 23799 25248 35440 25276
rect 23799 25245 23811 25248
rect 23753 25239 23811 25245
rect 2041 25211 2099 25217
rect 2041 25177 2053 25211
rect 2087 25208 2099 25211
rect 2590 25208 2596 25220
rect 2087 25180 2596 25208
rect 2087 25177 2099 25180
rect 2041 25171 2099 25177
rect 2590 25168 2596 25180
rect 2648 25168 2654 25220
rect 18230 25208 18236 25220
rect 18191 25180 18236 25208
rect 18230 25168 18236 25180
rect 18288 25168 18294 25220
rect 19334 25168 19340 25220
rect 19392 25208 19398 25220
rect 19392 25180 21588 25208
rect 19392 25168 19398 25180
rect 19242 25140 19248 25152
rect 19203 25112 19248 25140
rect 19242 25100 19248 25112
rect 19300 25100 19306 25152
rect 20622 25100 20628 25152
rect 20680 25140 20686 25152
rect 20717 25143 20775 25149
rect 20717 25140 20729 25143
rect 20680 25112 20729 25140
rect 20680 25100 20686 25112
rect 20717 25109 20729 25112
rect 20763 25109 20775 25143
rect 21174 25140 21180 25152
rect 21135 25112 21180 25140
rect 20717 25103 20775 25109
rect 21174 25100 21180 25112
rect 21232 25100 21238 25152
rect 21560 25149 21588 25180
rect 21545 25143 21603 25149
rect 21545 25109 21557 25143
rect 21591 25140 21603 25143
rect 23768 25140 23796 25239
rect 35434 25236 35440 25248
rect 35492 25236 35498 25288
rect 37461 25279 37519 25285
rect 37461 25245 37473 25279
rect 37507 25276 37519 25279
rect 38102 25276 38108 25288
rect 37507 25248 38108 25276
rect 37507 25245 37519 25248
rect 37461 25239 37519 25245
rect 38102 25236 38108 25248
rect 38160 25236 38166 25288
rect 25038 25208 25044 25220
rect 24951 25180 25044 25208
rect 25038 25168 25044 25180
rect 25096 25208 25102 25220
rect 25096 25180 35894 25208
rect 25096 25168 25102 25180
rect 21591 25112 23796 25140
rect 21591 25109 21603 25112
rect 21545 25103 21603 25109
rect 24394 25100 24400 25152
rect 24452 25140 24458 25152
rect 26234 25140 26240 25152
rect 24452 25112 26240 25140
rect 24452 25100 24458 25112
rect 26234 25100 26240 25112
rect 26292 25140 26298 25152
rect 26789 25143 26847 25149
rect 26789 25140 26801 25143
rect 26292 25112 26801 25140
rect 26292 25100 26298 25112
rect 26789 25109 26801 25112
rect 26835 25140 26847 25143
rect 27062 25140 27068 25152
rect 26835 25112 27068 25140
rect 26835 25109 26847 25112
rect 26789 25103 26847 25109
rect 27062 25100 27068 25112
rect 27120 25100 27126 25152
rect 35866 25140 35894 25180
rect 37826 25140 37832 25152
rect 35866 25112 37832 25140
rect 37826 25100 37832 25112
rect 37884 25100 37890 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 22002 24936 22008 24948
rect 21963 24908 22008 24936
rect 22002 24896 22008 24908
rect 22060 24896 22066 24948
rect 22833 24939 22891 24945
rect 22833 24905 22845 24939
rect 22879 24905 22891 24939
rect 23658 24936 23664 24948
rect 23619 24908 23664 24936
rect 22833 24899 22891 24905
rect 22848 24868 22876 24899
rect 23658 24896 23664 24908
rect 23716 24896 23722 24948
rect 23382 24868 23388 24880
rect 22848 24840 23388 24868
rect 23382 24828 23388 24840
rect 23440 24868 23446 24880
rect 25038 24868 25044 24880
rect 23440 24840 25044 24868
rect 23440 24828 23446 24840
rect 25038 24828 25044 24840
rect 25096 24828 25102 24880
rect 1394 24800 1400 24812
rect 1355 24772 1400 24800
rect 1394 24760 1400 24772
rect 1452 24800 1458 24812
rect 2041 24803 2099 24809
rect 2041 24800 2053 24803
rect 1452 24772 2053 24800
rect 1452 24760 1458 24772
rect 2041 24769 2053 24772
rect 2087 24769 2099 24803
rect 17954 24800 17960 24812
rect 17915 24772 17960 24800
rect 2041 24763 2099 24769
rect 17954 24760 17960 24772
rect 18012 24760 18018 24812
rect 19242 24800 19248 24812
rect 19203 24772 19248 24800
rect 19242 24760 19248 24772
rect 19300 24760 19306 24812
rect 21174 24760 21180 24812
rect 21232 24800 21238 24812
rect 21269 24803 21327 24809
rect 21269 24800 21281 24803
rect 21232 24772 21281 24800
rect 21232 24760 21238 24772
rect 21269 24769 21281 24772
rect 21315 24769 21327 24803
rect 21818 24800 21824 24812
rect 21779 24772 21824 24800
rect 21269 24763 21327 24769
rect 21818 24760 21824 24772
rect 21876 24760 21882 24812
rect 24029 24803 24087 24809
rect 22066 24772 23336 24800
rect 18966 24732 18972 24744
rect 18927 24704 18972 24732
rect 18966 24692 18972 24704
rect 19024 24692 19030 24744
rect 20990 24732 20996 24744
rect 20951 24704 20996 24732
rect 20990 24692 20996 24704
rect 21048 24692 21054 24744
rect 21082 24692 21088 24744
rect 21140 24732 21146 24744
rect 22066 24732 22094 24772
rect 21140 24704 22094 24732
rect 21140 24692 21146 24704
rect 22278 24692 22284 24744
rect 22336 24732 22342 24744
rect 22557 24735 22615 24741
rect 22557 24732 22569 24735
rect 22336 24704 22569 24732
rect 22336 24692 22342 24704
rect 22557 24701 22569 24704
rect 22603 24701 22615 24735
rect 22557 24695 22615 24701
rect 22741 24735 22799 24741
rect 22741 24701 22753 24735
rect 22787 24701 22799 24735
rect 22741 24695 22799 24701
rect 1581 24667 1639 24673
rect 1581 24633 1593 24667
rect 1627 24664 1639 24667
rect 19889 24667 19947 24673
rect 19889 24664 19901 24667
rect 1627 24636 19901 24664
rect 1627 24633 1639 24636
rect 1581 24627 1639 24633
rect 19889 24633 19901 24636
rect 19935 24664 19947 24667
rect 19935 24636 22094 24664
rect 19935 24633 19947 24636
rect 19889 24627 19947 24633
rect 22066 24596 22094 24636
rect 22756 24596 22784 24695
rect 22066 24568 22784 24596
rect 23106 24556 23112 24608
rect 23164 24596 23170 24608
rect 23201 24599 23259 24605
rect 23201 24596 23213 24599
rect 23164 24568 23213 24596
rect 23164 24556 23170 24568
rect 23201 24565 23213 24568
rect 23247 24565 23259 24599
rect 23308 24596 23336 24772
rect 24029 24769 24041 24803
rect 24075 24800 24087 24803
rect 25314 24800 25320 24812
rect 24075 24772 24808 24800
rect 25275 24772 25320 24800
rect 24075 24769 24087 24772
rect 24029 24763 24087 24769
rect 24780 24744 24808 24772
rect 25314 24760 25320 24772
rect 25372 24760 25378 24812
rect 37461 24803 37519 24809
rect 25424 24772 35894 24800
rect 24121 24735 24179 24741
rect 24121 24701 24133 24735
rect 24167 24701 24179 24735
rect 24121 24695 24179 24701
rect 24136 24664 24164 24695
rect 24210 24692 24216 24744
rect 24268 24732 24274 24744
rect 24268 24704 24313 24732
rect 24268 24692 24274 24704
rect 24762 24692 24768 24744
rect 24820 24732 24826 24744
rect 25424 24732 25452 24772
rect 24820 24704 25452 24732
rect 25869 24735 25927 24741
rect 24820 24692 24826 24704
rect 25869 24701 25881 24735
rect 25915 24732 25927 24735
rect 33410 24732 33416 24744
rect 25915 24704 33416 24732
rect 25915 24701 25927 24704
rect 25869 24695 25927 24701
rect 25222 24664 25228 24676
rect 24136 24636 25228 24664
rect 25222 24624 25228 24636
rect 25280 24624 25286 24676
rect 25884 24596 25912 24695
rect 33410 24692 33416 24704
rect 33468 24692 33474 24744
rect 35866 24664 35894 24772
rect 37461 24769 37473 24803
rect 37507 24800 37519 24803
rect 38102 24800 38108 24812
rect 37507 24772 38108 24800
rect 37507 24769 37519 24772
rect 37461 24763 37519 24769
rect 38102 24760 38108 24772
rect 38160 24760 38166 24812
rect 37921 24667 37979 24673
rect 37921 24664 37933 24667
rect 35866 24636 37933 24664
rect 37921 24633 37933 24636
rect 37967 24633 37979 24667
rect 37921 24627 37979 24633
rect 27890 24596 27896 24608
rect 23308 24568 25912 24596
rect 27851 24568 27896 24596
rect 23201 24559 23259 24565
rect 27890 24556 27896 24568
rect 27948 24556 27954 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 18509 24395 18567 24401
rect 18509 24361 18521 24395
rect 18555 24392 18567 24395
rect 19334 24392 19340 24404
rect 18555 24364 19340 24392
rect 18555 24361 18567 24364
rect 18509 24355 18567 24361
rect 19334 24352 19340 24364
rect 19392 24352 19398 24404
rect 22554 24352 22560 24404
rect 22612 24392 22618 24404
rect 23661 24395 23719 24401
rect 23661 24392 23673 24395
rect 22612 24364 23673 24392
rect 22612 24352 22618 24364
rect 23661 24361 23673 24364
rect 23707 24361 23719 24395
rect 24762 24392 24768 24404
rect 24723 24364 24768 24392
rect 23661 24355 23719 24361
rect 24762 24352 24768 24364
rect 24820 24352 24826 24404
rect 29641 24395 29699 24401
rect 29641 24392 29653 24395
rect 28276 24364 29653 24392
rect 16206 24284 16212 24336
rect 16264 24324 16270 24336
rect 21637 24327 21695 24333
rect 16264 24296 20208 24324
rect 16264 24284 16270 24296
rect 20180 24265 20208 24296
rect 21637 24293 21649 24327
rect 21683 24324 21695 24327
rect 21910 24324 21916 24336
rect 21683 24296 21916 24324
rect 21683 24293 21695 24296
rect 21637 24287 21695 24293
rect 21910 24284 21916 24296
rect 21968 24284 21974 24336
rect 23477 24327 23535 24333
rect 23477 24324 23489 24327
rect 23032 24296 23489 24324
rect 17589 24259 17647 24265
rect 17589 24225 17601 24259
rect 17635 24256 17647 24259
rect 20165 24259 20223 24265
rect 17635 24228 18552 24256
rect 17635 24225 17647 24228
rect 17589 24219 17647 24225
rect 13541 24191 13599 24197
rect 13541 24157 13553 24191
rect 13587 24188 13599 24191
rect 13630 24188 13636 24200
rect 13587 24160 13636 24188
rect 13587 24157 13599 24160
rect 13541 24151 13599 24157
rect 13630 24148 13636 24160
rect 13688 24148 13694 24200
rect 17037 24191 17095 24197
rect 17037 24157 17049 24191
rect 17083 24188 17095 24191
rect 18322 24188 18328 24200
rect 17083 24160 18328 24188
rect 17083 24157 17095 24160
rect 17037 24151 17095 24157
rect 18322 24148 18328 24160
rect 18380 24148 18386 24200
rect 18524 24197 18552 24228
rect 20165 24225 20177 24259
rect 20211 24225 20223 24259
rect 21450 24256 21456 24268
rect 21411 24228 21456 24256
rect 20165 24219 20223 24225
rect 21450 24216 21456 24228
rect 21508 24216 21514 24268
rect 23032 24265 23060 24296
rect 23477 24293 23489 24296
rect 23523 24293 23535 24327
rect 23477 24287 23535 24293
rect 23017 24259 23075 24265
rect 23017 24225 23029 24259
rect 23063 24225 23075 24259
rect 23017 24219 23075 24225
rect 23198 24216 23204 24268
rect 23256 24256 23262 24268
rect 24673 24259 24731 24265
rect 24673 24256 24685 24259
rect 23256 24228 24685 24256
rect 23256 24216 23262 24228
rect 24673 24225 24685 24228
rect 24719 24256 24731 24259
rect 25869 24259 25927 24265
rect 25869 24256 25881 24259
rect 24719 24228 25881 24256
rect 24719 24225 24731 24228
rect 24673 24219 24731 24225
rect 25869 24225 25881 24228
rect 25915 24256 25927 24259
rect 25915 24228 26234 24256
rect 25915 24225 25927 24228
rect 25869 24219 25927 24225
rect 18509 24191 18567 24197
rect 18509 24157 18521 24191
rect 18555 24188 18567 24191
rect 19426 24188 19432 24200
rect 18555 24160 19432 24188
rect 18555 24157 18567 24160
rect 18509 24151 18567 24157
rect 19426 24148 19432 24160
rect 19484 24148 19490 24200
rect 19889 24191 19947 24197
rect 19889 24157 19901 24191
rect 19935 24188 19947 24191
rect 20070 24188 20076 24200
rect 19935 24160 20076 24188
rect 19935 24157 19947 24160
rect 19889 24151 19947 24157
rect 20070 24148 20076 24160
rect 20128 24148 20134 24200
rect 21729 24191 21787 24197
rect 21729 24157 21741 24191
rect 21775 24188 21787 24191
rect 22462 24188 22468 24200
rect 21775 24160 22468 24188
rect 21775 24157 21787 24160
rect 21729 24151 21787 24157
rect 22462 24148 22468 24160
rect 22520 24148 22526 24200
rect 22738 24188 22744 24200
rect 22699 24160 22744 24188
rect 22738 24148 22744 24160
rect 22796 24148 22802 24200
rect 24486 24148 24492 24200
rect 24544 24188 24550 24200
rect 24581 24191 24639 24197
rect 24581 24188 24593 24191
rect 24544 24160 24593 24188
rect 24544 24148 24550 24160
rect 24581 24157 24593 24160
rect 24627 24157 24639 24191
rect 24854 24188 24860 24200
rect 24815 24160 24860 24188
rect 24581 24151 24639 24157
rect 1854 24120 1860 24132
rect 1815 24092 1860 24120
rect 1854 24080 1860 24092
rect 1912 24080 1918 24132
rect 2038 24120 2044 24132
rect 1999 24092 2044 24120
rect 2038 24080 2044 24092
rect 2096 24080 2102 24132
rect 2222 24080 2228 24132
rect 2280 24120 2286 24132
rect 2280 24092 2774 24120
rect 2280 24080 2286 24092
rect 1872 24052 1900 24080
rect 2501 24055 2559 24061
rect 2501 24052 2513 24055
rect 1872 24024 2513 24052
rect 2501 24021 2513 24024
rect 2547 24021 2559 24055
rect 2746 24052 2774 24092
rect 17954 24080 17960 24132
rect 18012 24120 18018 24132
rect 18049 24123 18107 24129
rect 18049 24120 18061 24123
rect 18012 24092 18061 24120
rect 18012 24080 18018 24092
rect 18049 24089 18061 24092
rect 18095 24089 18107 24123
rect 18049 24083 18107 24089
rect 20898 24080 20904 24132
rect 20956 24120 20962 24132
rect 21910 24120 21916 24132
rect 20956 24092 21916 24120
rect 20956 24080 20962 24092
rect 21910 24080 21916 24092
rect 21968 24080 21974 24132
rect 22370 24120 22376 24132
rect 22066 24092 22376 24120
rect 13357 24055 13415 24061
rect 13357 24052 13369 24055
rect 2746 24024 13369 24052
rect 2501 24015 2559 24021
rect 13357 24021 13369 24024
rect 13403 24021 13415 24055
rect 18690 24052 18696 24064
rect 18651 24024 18696 24052
rect 13357 24015 13415 24021
rect 18690 24012 18696 24024
rect 18748 24012 18754 24064
rect 21729 24055 21787 24061
rect 21729 24021 21741 24055
rect 21775 24052 21787 24055
rect 22066 24052 22094 24092
rect 22370 24080 22376 24092
rect 22428 24120 22434 24132
rect 23845 24123 23903 24129
rect 23845 24120 23857 24123
rect 22428 24092 23857 24120
rect 22428 24080 22434 24092
rect 23845 24089 23857 24092
rect 23891 24089 23903 24123
rect 24596 24120 24624 24151
rect 24854 24148 24860 24160
rect 24912 24148 24918 24200
rect 26206 24188 26234 24228
rect 27890 24216 27896 24268
rect 27948 24256 27954 24268
rect 28276 24265 28304 24364
rect 29641 24361 29653 24364
rect 29687 24392 29699 24395
rect 36538 24392 36544 24404
rect 29687 24364 36544 24392
rect 29687 24361 29699 24364
rect 29641 24355 29699 24361
rect 36538 24352 36544 24364
rect 36596 24352 36602 24404
rect 28077 24259 28135 24265
rect 28077 24256 28089 24259
rect 27948 24228 28089 24256
rect 27948 24216 27954 24228
rect 28077 24225 28089 24228
rect 28123 24225 28135 24259
rect 28077 24219 28135 24225
rect 28261 24259 28319 24265
rect 28261 24225 28273 24259
rect 28307 24225 28319 24259
rect 37642 24256 37648 24268
rect 28261 24219 28319 24225
rect 28460 24228 37648 24256
rect 28460 24188 28488 24228
rect 37642 24216 37648 24228
rect 37700 24216 37706 24268
rect 26206 24160 28488 24188
rect 29454 24148 29460 24200
rect 29512 24188 29518 24200
rect 37829 24191 37887 24197
rect 37829 24188 37841 24191
rect 29512 24160 37841 24188
rect 29512 24148 29518 24160
rect 37829 24157 37841 24160
rect 37875 24157 37887 24191
rect 37829 24151 37887 24157
rect 27433 24123 27491 24129
rect 27433 24120 27445 24123
rect 24596 24092 27445 24120
rect 23845 24083 23903 24089
rect 27433 24089 27445 24092
rect 27479 24120 27491 24123
rect 28353 24123 28411 24129
rect 28353 24120 28365 24123
rect 27479 24092 28365 24120
rect 27479 24089 27491 24092
rect 27433 24083 27491 24089
rect 28353 24089 28365 24092
rect 28399 24089 28411 24123
rect 28353 24083 28411 24089
rect 21775 24024 22094 24052
rect 21775 24021 21787 24024
rect 21729 24015 21787 24021
rect 23290 24012 23296 24064
rect 23348 24052 23354 24064
rect 23635 24055 23693 24061
rect 23635 24052 23647 24055
rect 23348 24024 23647 24052
rect 23348 24012 23354 24024
rect 23635 24021 23647 24024
rect 23681 24021 23693 24055
rect 24394 24052 24400 24064
rect 24355 24024 24400 24052
rect 23635 24015 23693 24021
rect 24394 24012 24400 24024
rect 24452 24012 24458 24064
rect 25222 24012 25228 24064
rect 25280 24052 25286 24064
rect 25317 24055 25375 24061
rect 25317 24052 25329 24055
rect 25280 24024 25329 24052
rect 25280 24012 25286 24024
rect 25317 24021 25329 24024
rect 25363 24021 25375 24055
rect 25317 24015 25375 24021
rect 28534 24012 28540 24064
rect 28592 24052 28598 24064
rect 28721 24055 28779 24061
rect 28721 24052 28733 24055
rect 28592 24024 28733 24052
rect 28592 24012 28598 24024
rect 28721 24021 28733 24024
rect 28767 24021 28779 24055
rect 38010 24052 38016 24064
rect 37971 24024 38016 24052
rect 28721 24015 28779 24021
rect 38010 24012 38016 24024
rect 38068 24012 38074 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 13630 23848 13636 23860
rect 13591 23820 13636 23848
rect 13630 23808 13636 23820
rect 13688 23808 13694 23860
rect 21542 23848 21548 23860
rect 16960 23820 21548 23848
rect 2225 23783 2283 23789
rect 2225 23780 2237 23783
rect 1688 23752 2237 23780
rect 1688 23721 1716 23752
rect 2225 23749 2237 23752
rect 2271 23780 2283 23783
rect 16960 23780 16988 23820
rect 21542 23808 21548 23820
rect 21600 23808 21606 23860
rect 21818 23848 21824 23860
rect 21779 23820 21824 23848
rect 21818 23808 21824 23820
rect 21876 23808 21882 23860
rect 21910 23808 21916 23860
rect 21968 23848 21974 23860
rect 24210 23848 24216 23860
rect 21968 23820 24216 23848
rect 21968 23808 21974 23820
rect 24210 23808 24216 23820
rect 24268 23848 24274 23860
rect 24489 23851 24547 23857
rect 24489 23848 24501 23851
rect 24268 23820 24501 23848
rect 24268 23808 24274 23820
rect 24489 23817 24501 23820
rect 24535 23817 24547 23851
rect 24489 23811 24547 23817
rect 2271 23752 16988 23780
rect 17589 23783 17647 23789
rect 2271 23749 2283 23752
rect 2225 23743 2283 23749
rect 17589 23749 17601 23783
rect 17635 23780 17647 23783
rect 18049 23783 18107 23789
rect 18049 23780 18061 23783
rect 17635 23752 18061 23780
rect 17635 23749 17647 23752
rect 17589 23743 17647 23749
rect 18049 23749 18061 23752
rect 18095 23780 18107 23783
rect 18138 23780 18144 23792
rect 18095 23752 18144 23780
rect 18095 23749 18107 23752
rect 18049 23743 18107 23749
rect 18138 23740 18144 23752
rect 18196 23740 18202 23792
rect 24394 23780 24400 23792
rect 21284 23752 24400 23780
rect 1673 23715 1731 23721
rect 1673 23681 1685 23715
rect 1719 23681 1731 23715
rect 1673 23675 1731 23681
rect 14001 23715 14059 23721
rect 14001 23681 14013 23715
rect 14047 23712 14059 23715
rect 14047 23684 14964 23712
rect 14047 23681 14059 23684
rect 14001 23675 14059 23681
rect 8202 23604 8208 23656
rect 8260 23644 8266 23656
rect 13173 23647 13231 23653
rect 13173 23644 13185 23647
rect 8260 23616 13185 23644
rect 8260 23604 8266 23616
rect 13173 23613 13185 23616
rect 13219 23644 13231 23647
rect 14093 23647 14151 23653
rect 14093 23644 14105 23647
rect 13219 23616 14105 23644
rect 13219 23613 13231 23616
rect 13173 23607 13231 23613
rect 14093 23613 14105 23616
rect 14139 23613 14151 23647
rect 14093 23607 14151 23613
rect 14277 23647 14335 23653
rect 14277 23613 14289 23647
rect 14323 23644 14335 23647
rect 14550 23644 14556 23656
rect 14323 23616 14556 23644
rect 14323 23613 14335 23616
rect 14277 23607 14335 23613
rect 14550 23604 14556 23616
rect 14608 23604 14614 23656
rect 1486 23508 1492 23520
rect 1447 23480 1492 23508
rect 1486 23468 1492 23480
rect 1544 23468 1550 23520
rect 14936 23517 14964 23684
rect 17954 23672 17960 23724
rect 18012 23712 18018 23724
rect 18230 23712 18236 23724
rect 18012 23684 18236 23712
rect 18012 23672 18018 23684
rect 18230 23672 18236 23684
rect 18288 23672 18294 23724
rect 18690 23672 18696 23724
rect 18748 23712 18754 23724
rect 21284 23721 21312 23752
rect 24394 23740 24400 23752
rect 24452 23740 24458 23792
rect 21085 23715 21143 23721
rect 21085 23712 21097 23715
rect 18748 23684 21097 23712
rect 18748 23672 18754 23684
rect 21085 23681 21097 23684
rect 21131 23681 21143 23715
rect 21085 23675 21143 23681
rect 21269 23715 21327 23721
rect 21269 23681 21281 23715
rect 21315 23681 21327 23715
rect 21269 23675 21327 23681
rect 21726 23672 21732 23724
rect 21784 23712 21790 23724
rect 22189 23715 22247 23721
rect 22189 23712 22201 23715
rect 21784 23684 22201 23712
rect 21784 23672 21790 23684
rect 22189 23681 22201 23684
rect 22235 23681 22247 23715
rect 23106 23712 23112 23724
rect 23067 23684 23112 23712
rect 22189 23675 22247 23681
rect 23106 23672 23112 23684
rect 23164 23672 23170 23724
rect 18877 23647 18935 23653
rect 18877 23613 18889 23647
rect 18923 23613 18935 23647
rect 19426 23644 19432 23656
rect 19387 23616 19432 23644
rect 18877 23607 18935 23613
rect 14921 23511 14979 23517
rect 14921 23477 14933 23511
rect 14967 23508 14979 23511
rect 15194 23508 15200 23520
rect 14967 23480 15200 23508
rect 14967 23477 14979 23480
rect 14921 23471 14979 23477
rect 15194 23468 15200 23480
rect 15252 23468 15258 23520
rect 18892 23508 18920 23607
rect 19426 23604 19432 23616
rect 19484 23604 19490 23656
rect 19705 23647 19763 23653
rect 19705 23613 19717 23647
rect 19751 23613 19763 23647
rect 22278 23644 22284 23656
rect 22239 23616 22284 23644
rect 19705 23607 19763 23613
rect 19334 23536 19340 23588
rect 19392 23576 19398 23588
rect 19720 23576 19748 23607
rect 22278 23604 22284 23616
rect 22336 23604 22342 23656
rect 22370 23604 22376 23656
rect 22428 23644 22434 23656
rect 23382 23644 23388 23656
rect 22428 23616 22473 23644
rect 23343 23616 23388 23644
rect 22428 23604 22434 23616
rect 23382 23604 23388 23616
rect 23440 23604 23446 23656
rect 19392 23548 19748 23576
rect 21269 23579 21327 23585
rect 19392 23536 19398 23548
rect 21269 23545 21281 23579
rect 21315 23576 21327 23579
rect 22554 23576 22560 23588
rect 21315 23548 22560 23576
rect 21315 23545 21327 23548
rect 21269 23539 21327 23545
rect 22554 23536 22560 23548
rect 22612 23576 22618 23588
rect 23290 23576 23296 23588
rect 22612 23548 23296 23576
rect 22612 23536 22618 23548
rect 23290 23536 23296 23548
rect 23348 23536 23354 23588
rect 24504 23576 24532 23811
rect 24854 23808 24860 23860
rect 24912 23848 24918 23860
rect 27617 23851 27675 23857
rect 27617 23848 27629 23851
rect 24912 23820 27629 23848
rect 24912 23808 24918 23820
rect 27617 23817 27629 23820
rect 27663 23848 27675 23851
rect 28445 23851 28503 23857
rect 28445 23848 28457 23851
rect 27663 23820 28457 23848
rect 27663 23817 27675 23820
rect 27617 23811 27675 23817
rect 28445 23817 28457 23820
rect 28491 23817 28503 23851
rect 29454 23848 29460 23860
rect 29415 23820 29460 23848
rect 28445 23811 28503 23817
rect 29454 23808 29460 23820
rect 29512 23808 29518 23860
rect 37366 23848 37372 23860
rect 37327 23820 37372 23848
rect 37366 23808 37372 23820
rect 37424 23808 37430 23860
rect 29273 23715 29331 23721
rect 29273 23712 29285 23715
rect 28828 23684 29285 23712
rect 27890 23644 27896 23656
rect 26206 23616 27896 23644
rect 26206 23576 26234 23616
rect 27890 23604 27896 23616
rect 27948 23644 27954 23656
rect 28169 23647 28227 23653
rect 28169 23644 28181 23647
rect 27948 23616 28181 23644
rect 27948 23604 27954 23616
rect 28169 23613 28181 23616
rect 28215 23613 28227 23647
rect 28169 23607 28227 23613
rect 28353 23647 28411 23653
rect 28353 23613 28365 23647
rect 28399 23613 28411 23647
rect 28353 23607 28411 23613
rect 24504 23548 26234 23576
rect 22370 23508 22376 23520
rect 18892 23480 22376 23508
rect 22370 23468 22376 23480
rect 22428 23468 22434 23520
rect 24486 23468 24492 23520
rect 24544 23508 24550 23520
rect 24949 23511 25007 23517
rect 24949 23508 24961 23511
rect 24544 23480 24961 23508
rect 24544 23468 24550 23480
rect 24949 23477 24961 23480
rect 24995 23477 25007 23511
rect 28368 23508 28396 23607
rect 28828 23585 28856 23684
rect 29273 23681 29285 23684
rect 29319 23681 29331 23715
rect 37384 23712 37412 23808
rect 37829 23715 37887 23721
rect 37829 23712 37841 23715
rect 37384 23684 37841 23712
rect 29273 23675 29331 23681
rect 37829 23681 37841 23684
rect 37875 23681 37887 23715
rect 37829 23675 37887 23681
rect 28813 23579 28871 23585
rect 28813 23545 28825 23579
rect 28859 23545 28871 23579
rect 28813 23539 28871 23545
rect 29914 23508 29920 23520
rect 28368 23480 29920 23508
rect 24949 23471 25007 23477
rect 29914 23468 29920 23480
rect 29972 23468 29978 23520
rect 38010 23508 38016 23520
rect 37971 23480 38016 23508
rect 38010 23468 38016 23480
rect 38068 23468 38074 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 18322 23264 18328 23316
rect 18380 23304 18386 23316
rect 18598 23304 18604 23316
rect 18380 23276 18604 23304
rect 18380 23264 18386 23276
rect 18598 23264 18604 23276
rect 18656 23264 18662 23316
rect 19245 23307 19303 23313
rect 19245 23273 19257 23307
rect 19291 23304 19303 23307
rect 19426 23304 19432 23316
rect 19291 23276 19432 23304
rect 19291 23273 19303 23276
rect 19245 23267 19303 23273
rect 19426 23264 19432 23276
rect 19484 23264 19490 23316
rect 20070 23264 20076 23316
rect 20128 23304 20134 23316
rect 20441 23307 20499 23313
rect 20441 23304 20453 23307
rect 20128 23276 20453 23304
rect 20128 23264 20134 23276
rect 20441 23273 20453 23276
rect 20487 23273 20499 23307
rect 20441 23267 20499 23273
rect 24489 23307 24547 23313
rect 24489 23273 24501 23307
rect 24535 23304 24547 23307
rect 24854 23304 24860 23316
rect 24535 23276 24860 23304
rect 24535 23273 24547 23276
rect 24489 23267 24547 23273
rect 24854 23264 24860 23276
rect 24912 23264 24918 23316
rect 27890 23304 27896 23316
rect 27851 23276 27896 23304
rect 27890 23264 27896 23276
rect 27948 23264 27954 23316
rect 5074 23196 5080 23248
rect 5132 23236 5138 23248
rect 5132 23208 12434 23236
rect 5132 23196 5138 23208
rect 10318 23168 10324 23180
rect 10279 23140 10324 23168
rect 10318 23128 10324 23140
rect 10376 23128 10382 23180
rect 10045 23103 10103 23109
rect 10045 23069 10057 23103
rect 10091 23100 10103 23103
rect 10226 23100 10232 23112
rect 10091 23072 10232 23100
rect 10091 23069 10103 23072
rect 10045 23063 10103 23069
rect 10226 23060 10232 23072
rect 10284 23060 10290 23112
rect 12406 23100 12434 23208
rect 20622 23196 20628 23248
rect 20680 23236 20686 23248
rect 22554 23236 22560 23248
rect 20680 23208 21036 23236
rect 20680 23196 20686 23208
rect 15194 23128 15200 23180
rect 15252 23168 15258 23180
rect 15252 23140 16804 23168
rect 15252 23128 15258 23140
rect 16301 23103 16359 23109
rect 16301 23100 16313 23103
rect 12406 23072 16313 23100
rect 16301 23069 16313 23072
rect 16347 23069 16359 23103
rect 16301 23063 16359 23069
rect 16577 23103 16635 23109
rect 16577 23069 16589 23103
rect 16623 23100 16635 23103
rect 16666 23100 16672 23112
rect 16623 23072 16672 23100
rect 16623 23069 16635 23072
rect 16577 23063 16635 23069
rect 16666 23060 16672 23072
rect 16724 23060 16730 23112
rect 16776 23100 16804 23140
rect 18506 23128 18512 23180
rect 18564 23168 18570 23180
rect 19705 23171 19763 23177
rect 19705 23168 19717 23171
rect 18564 23140 19717 23168
rect 18564 23128 18570 23140
rect 19705 23137 19717 23140
rect 19751 23137 19763 23171
rect 19705 23131 19763 23137
rect 19889 23171 19947 23177
rect 19889 23137 19901 23171
rect 19935 23168 19947 23171
rect 19978 23168 19984 23180
rect 19935 23140 19984 23168
rect 19935 23137 19947 23140
rect 19889 23131 19947 23137
rect 19978 23128 19984 23140
rect 20036 23168 20042 23180
rect 20898 23168 20904 23180
rect 20036 23140 20904 23168
rect 20036 23128 20042 23140
rect 20898 23128 20904 23140
rect 20956 23128 20962 23180
rect 21008 23177 21036 23208
rect 22296 23208 22560 23236
rect 22296 23177 22324 23208
rect 22554 23196 22560 23208
rect 22612 23196 22618 23248
rect 23477 23239 23535 23245
rect 23477 23205 23489 23239
rect 23523 23236 23535 23239
rect 26234 23236 26240 23248
rect 23523 23208 26240 23236
rect 23523 23205 23535 23208
rect 23477 23199 23535 23205
rect 26234 23196 26240 23208
rect 26292 23236 26298 23248
rect 26786 23236 26792 23248
rect 26292 23208 26792 23236
rect 26292 23196 26298 23208
rect 26786 23196 26792 23208
rect 26844 23196 26850 23248
rect 20993 23171 21051 23177
rect 20993 23137 21005 23171
rect 21039 23168 21051 23171
rect 22281 23171 22339 23177
rect 22281 23168 22293 23171
rect 21039 23140 22293 23168
rect 21039 23137 21051 23140
rect 20993 23131 21051 23137
rect 22281 23137 22293 23140
rect 22327 23137 22339 23171
rect 22281 23131 22339 23137
rect 22370 23128 22376 23180
rect 22428 23168 22434 23180
rect 22465 23171 22523 23177
rect 22465 23168 22477 23171
rect 22428 23140 22477 23168
rect 22428 23128 22434 23140
rect 22465 23137 22477 23140
rect 22511 23168 22523 23171
rect 23014 23168 23020 23180
rect 22511 23140 23020 23168
rect 22511 23137 22523 23140
rect 22465 23131 22523 23137
rect 23014 23128 23020 23140
rect 23072 23128 23078 23180
rect 22922 23100 22928 23112
rect 16776 23072 22928 23100
rect 22922 23060 22928 23072
rect 22980 23060 22986 23112
rect 28534 23100 28540 23112
rect 28495 23072 28540 23100
rect 28534 23060 28540 23072
rect 28592 23060 28598 23112
rect 19518 22992 19524 23044
rect 19576 23032 19582 23044
rect 19613 23035 19671 23041
rect 19613 23032 19625 23035
rect 19576 23004 19625 23032
rect 19576 22992 19582 23004
rect 19613 23001 19625 23004
rect 19659 23032 19671 23035
rect 20254 23032 20260 23044
rect 19659 23004 20260 23032
rect 19659 23001 19671 23004
rect 19613 22995 19671 23001
rect 20254 22992 20260 23004
rect 20312 22992 20318 23044
rect 22557 23035 22615 23041
rect 22557 23001 22569 23035
rect 22603 23032 22615 23035
rect 23658 23032 23664 23044
rect 22603 23004 23664 23032
rect 22603 23001 22615 23004
rect 22557 22995 22615 23001
rect 23658 22992 23664 23004
rect 23716 22992 23722 23044
rect 14550 22964 14556 22976
rect 14511 22936 14556 22964
rect 14550 22924 14556 22936
rect 14608 22924 14614 22976
rect 18598 22924 18604 22976
rect 18656 22964 18662 22976
rect 20809 22967 20867 22973
rect 20809 22964 20821 22967
rect 18656 22936 20821 22964
rect 18656 22924 18662 22936
rect 20809 22933 20821 22936
rect 20855 22933 20867 22967
rect 20809 22927 20867 22933
rect 20898 22924 20904 22976
rect 20956 22964 20962 22976
rect 20956 22936 21001 22964
rect 20956 22924 20962 22936
rect 21634 22924 21640 22976
rect 21692 22964 21698 22976
rect 21729 22967 21787 22973
rect 21729 22964 21741 22967
rect 21692 22936 21741 22964
rect 21692 22924 21698 22936
rect 21729 22933 21741 22936
rect 21775 22964 21787 22967
rect 22278 22964 22284 22976
rect 21775 22936 22284 22964
rect 21775 22933 21787 22936
rect 21729 22927 21787 22933
rect 22278 22924 22284 22936
rect 22336 22924 22342 22976
rect 22925 22967 22983 22973
rect 22925 22933 22937 22967
rect 22971 22964 22983 22967
rect 23290 22964 23296 22976
rect 22971 22936 23296 22964
rect 22971 22933 22983 22936
rect 22925 22927 22983 22933
rect 23290 22924 23296 22936
rect 23348 22924 23354 22976
rect 28721 22967 28779 22973
rect 28721 22933 28733 22967
rect 28767 22964 28779 22967
rect 30834 22964 30840 22976
rect 28767 22936 30840 22964
rect 28767 22933 28779 22936
rect 28721 22927 28779 22933
rect 30834 22924 30840 22936
rect 30892 22924 30898 22976
rect 38102 22964 38108 22976
rect 38063 22936 38108 22964
rect 38102 22924 38108 22936
rect 38160 22924 38166 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 10226 22760 10232 22772
rect 10187 22732 10232 22760
rect 10226 22720 10232 22732
rect 10284 22720 10290 22772
rect 16666 22760 16672 22772
rect 16627 22732 16672 22760
rect 16666 22720 16672 22732
rect 16724 22720 16730 22772
rect 18506 22720 18512 22772
rect 18564 22760 18570 22772
rect 18601 22763 18659 22769
rect 18601 22760 18613 22763
rect 18564 22732 18613 22760
rect 18564 22720 18570 22732
rect 18601 22729 18613 22732
rect 18647 22729 18659 22763
rect 18601 22723 18659 22729
rect 19245 22763 19303 22769
rect 19245 22729 19257 22763
rect 19291 22760 19303 22763
rect 19978 22760 19984 22772
rect 19291 22732 19984 22760
rect 19291 22729 19303 22732
rect 19245 22723 19303 22729
rect 19978 22720 19984 22732
rect 20036 22720 20042 22772
rect 20070 22720 20076 22772
rect 20128 22760 20134 22772
rect 20254 22760 20260 22772
rect 20128 22732 20260 22760
rect 20128 22720 20134 22732
rect 20254 22720 20260 22732
rect 20312 22720 20318 22772
rect 20898 22720 20904 22772
rect 20956 22760 20962 22772
rect 21177 22763 21235 22769
rect 21177 22760 21189 22763
rect 20956 22732 21189 22760
rect 20956 22720 20962 22732
rect 21177 22729 21189 22732
rect 21223 22760 21235 22763
rect 21266 22760 21272 22772
rect 21223 22732 21272 22760
rect 21223 22729 21235 22732
rect 21177 22723 21235 22729
rect 21266 22720 21272 22732
rect 21324 22720 21330 22772
rect 21726 22720 21732 22772
rect 21784 22760 21790 22772
rect 21821 22763 21879 22769
rect 21821 22760 21833 22763
rect 21784 22732 21833 22760
rect 21784 22720 21790 22732
rect 21821 22729 21833 22732
rect 21867 22729 21879 22763
rect 22462 22760 22468 22772
rect 22423 22732 22468 22760
rect 21821 22723 21879 22729
rect 22462 22720 22468 22732
rect 22520 22720 22526 22772
rect 23566 22760 23572 22772
rect 23527 22732 23572 22760
rect 23566 22720 23572 22732
rect 23624 22720 23630 22772
rect 14550 22652 14556 22704
rect 14608 22692 14614 22704
rect 19705 22695 19763 22701
rect 19705 22692 19717 22695
rect 14608 22664 19717 22692
rect 14608 22652 14614 22664
rect 19705 22661 19717 22664
rect 19751 22692 19763 22695
rect 20622 22692 20628 22704
rect 19751 22664 20628 22692
rect 19751 22661 19763 22664
rect 19705 22655 19763 22661
rect 20622 22652 20628 22664
rect 20680 22652 20686 22704
rect 24578 22692 24584 22704
rect 22756 22664 24584 22692
rect 1394 22624 1400 22636
rect 1355 22596 1400 22624
rect 1394 22584 1400 22596
rect 1452 22624 1458 22636
rect 2041 22627 2099 22633
rect 2041 22624 2053 22627
rect 1452 22596 2053 22624
rect 1452 22584 1458 22596
rect 2041 22593 2053 22596
rect 2087 22593 2099 22627
rect 2041 22587 2099 22593
rect 9769 22627 9827 22633
rect 9769 22593 9781 22627
rect 9815 22624 9827 22627
rect 10502 22624 10508 22636
rect 9815 22596 10508 22624
rect 9815 22593 9827 22596
rect 9769 22587 9827 22593
rect 10502 22584 10508 22596
rect 10560 22624 10566 22636
rect 22756 22633 22784 22664
rect 24578 22652 24584 22664
rect 24636 22692 24642 22704
rect 24673 22695 24731 22701
rect 24673 22692 24685 22695
rect 24636 22664 24685 22692
rect 24636 22652 24642 22664
rect 24673 22661 24685 22664
rect 24719 22661 24731 22695
rect 24673 22655 24731 22661
rect 10597 22627 10655 22633
rect 10597 22624 10609 22627
rect 10560 22596 10609 22624
rect 10560 22584 10566 22596
rect 10597 22593 10609 22596
rect 10643 22593 10655 22627
rect 10597 22587 10655 22593
rect 10689 22627 10747 22633
rect 10689 22593 10701 22627
rect 10735 22624 10747 22627
rect 11517 22627 11575 22633
rect 11517 22624 11529 22627
rect 10735 22596 11529 22624
rect 10735 22593 10747 22596
rect 10689 22587 10747 22593
rect 11517 22593 11529 22596
rect 11563 22624 11575 22627
rect 17037 22627 17095 22633
rect 11563 22596 12434 22624
rect 11563 22593 11575 22596
rect 11517 22587 11575 22593
rect 10873 22559 10931 22565
rect 10873 22525 10885 22559
rect 10919 22556 10931 22559
rect 11146 22556 11152 22568
rect 10919 22528 11152 22556
rect 10919 22525 10931 22528
rect 10873 22519 10931 22525
rect 11146 22516 11152 22528
rect 11204 22516 11210 22568
rect 12406 22488 12434 22596
rect 17037 22593 17049 22627
rect 17083 22624 17095 22627
rect 22649 22627 22707 22633
rect 17083 22596 18000 22624
rect 17083 22593 17095 22596
rect 17037 22587 17095 22593
rect 17126 22556 17132 22568
rect 17087 22528 17132 22556
rect 17126 22516 17132 22528
rect 17184 22516 17190 22568
rect 17310 22556 17316 22568
rect 17271 22528 17316 22556
rect 17310 22516 17316 22528
rect 17368 22516 17374 22568
rect 17972 22565 18000 22596
rect 22649 22593 22661 22627
rect 22695 22593 22707 22627
rect 22649 22587 22707 22593
rect 22741 22627 22799 22633
rect 22741 22593 22753 22627
rect 22787 22593 22799 22627
rect 22922 22624 22928 22636
rect 22883 22596 22928 22624
rect 22741 22587 22799 22593
rect 17957 22559 18015 22565
rect 17957 22525 17969 22559
rect 18003 22556 18015 22559
rect 21450 22556 21456 22568
rect 18003 22528 21456 22556
rect 18003 22525 18015 22528
rect 17957 22519 18015 22525
rect 21450 22516 21456 22528
rect 21508 22516 21514 22568
rect 22664 22556 22692 22587
rect 22922 22584 22928 22596
rect 22980 22584 22986 22636
rect 23290 22584 23296 22636
rect 23348 22624 23354 22636
rect 23385 22627 23443 22633
rect 23385 22624 23397 22627
rect 23348 22596 23397 22624
rect 23348 22584 23354 22596
rect 23385 22593 23397 22596
rect 23431 22593 23443 22627
rect 23385 22587 23443 22593
rect 22830 22556 22836 22568
rect 22664 22528 22836 22556
rect 22830 22516 22836 22528
rect 22888 22516 22894 22568
rect 22940 22556 22968 22584
rect 24670 22556 24676 22568
rect 22940 22528 24676 22556
rect 24670 22516 24676 22528
rect 24728 22556 24734 22568
rect 25133 22559 25191 22565
rect 25133 22556 25145 22559
rect 24728 22528 25145 22556
rect 24728 22516 24734 22528
rect 25133 22525 25145 22528
rect 25179 22525 25191 22559
rect 37829 22559 37887 22565
rect 37829 22556 37841 22559
rect 25133 22519 25191 22525
rect 26206 22528 37841 22556
rect 26206 22488 26234 22528
rect 37829 22525 37841 22528
rect 37875 22525 37887 22559
rect 38102 22556 38108 22568
rect 38063 22528 38108 22556
rect 37829 22519 37887 22525
rect 38102 22516 38108 22528
rect 38160 22516 38166 22568
rect 12406 22460 26234 22488
rect 1578 22420 1584 22432
rect 1539 22392 1584 22420
rect 1578 22380 1584 22392
rect 1636 22380 1642 22432
rect 22925 22423 22983 22429
rect 22925 22389 22937 22423
rect 22971 22420 22983 22423
rect 23658 22420 23664 22432
rect 22971 22392 23664 22420
rect 22971 22389 22983 22392
rect 22925 22383 22983 22389
rect 23658 22380 23664 22392
rect 23716 22420 23722 22432
rect 24121 22423 24179 22429
rect 24121 22420 24133 22423
rect 23716 22392 24133 22420
rect 23716 22380 23722 22392
rect 24121 22389 24133 22392
rect 24167 22420 24179 22423
rect 24762 22420 24768 22432
rect 24167 22392 24768 22420
rect 24167 22389 24179 22392
rect 24121 22383 24179 22389
rect 24762 22380 24768 22392
rect 24820 22380 24826 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 1578 22176 1584 22228
rect 1636 22216 1642 22228
rect 17126 22216 17132 22228
rect 1636 22188 17132 22216
rect 1636 22176 1642 22188
rect 17126 22176 17132 22188
rect 17184 22176 17190 22228
rect 23566 22176 23572 22228
rect 23624 22216 23630 22228
rect 37366 22216 37372 22228
rect 23624 22188 37372 22216
rect 23624 22176 23630 22188
rect 37366 22176 37372 22188
rect 37424 22176 37430 22228
rect 37921 22151 37979 22157
rect 37921 22148 37933 22151
rect 20824 22120 37933 22148
rect 11146 22080 11152 22092
rect 11059 22052 11152 22080
rect 11146 22040 11152 22052
rect 11204 22080 11210 22092
rect 17954 22080 17960 22092
rect 11204 22052 17960 22080
rect 11204 22040 11210 22052
rect 17954 22040 17960 22052
rect 18012 22040 18018 22092
rect 20824 22089 20852 22120
rect 37921 22117 37933 22120
rect 37967 22117 37979 22151
rect 37921 22111 37979 22117
rect 20809 22083 20867 22089
rect 20809 22049 20821 22083
rect 20855 22080 20867 22083
rect 20993 22083 21051 22089
rect 20855 22052 20889 22080
rect 20855 22049 20867 22052
rect 20809 22043 20867 22049
rect 20993 22049 21005 22083
rect 21039 22080 21051 22083
rect 21082 22080 21088 22092
rect 21039 22052 21088 22080
rect 21039 22049 21051 22052
rect 20993 22043 21051 22049
rect 21082 22040 21088 22052
rect 21140 22040 21146 22092
rect 21913 22083 21971 22089
rect 21913 22049 21925 22083
rect 21959 22080 21971 22083
rect 22370 22080 22376 22092
rect 21959 22052 22376 22080
rect 21959 22049 21971 22052
rect 21913 22043 21971 22049
rect 22370 22040 22376 22052
rect 22428 22040 22434 22092
rect 22462 22040 22468 22092
rect 22520 22080 22526 22092
rect 22520 22052 22565 22080
rect 22520 22040 22526 22052
rect 1394 22012 1400 22024
rect 1355 21984 1400 22012
rect 1394 21972 1400 21984
rect 1452 22012 1458 22024
rect 2041 22015 2099 22021
rect 2041 22012 2053 22015
rect 1452 21984 2053 22012
rect 1452 21972 1458 21984
rect 2041 21981 2053 21984
rect 2087 21981 2099 22015
rect 2041 21975 2099 21981
rect 37461 22015 37519 22021
rect 37461 21981 37473 22015
rect 37507 22012 37519 22015
rect 38102 22012 38108 22024
rect 37507 21984 38108 22012
rect 37507 21981 37519 21984
rect 37461 21975 37519 21981
rect 38102 21972 38108 21984
rect 38160 21972 38166 22024
rect 19797 21947 19855 21953
rect 19797 21944 19809 21947
rect 6886 21916 19809 21944
rect 1581 21879 1639 21885
rect 1581 21845 1593 21879
rect 1627 21876 1639 21879
rect 1670 21876 1676 21888
rect 1627 21848 1676 21876
rect 1627 21845 1639 21848
rect 1581 21839 1639 21845
rect 1670 21836 1676 21848
rect 1728 21836 1734 21888
rect 3050 21836 3056 21888
rect 3108 21876 3114 21888
rect 6886 21876 6914 21916
rect 19797 21913 19809 21916
rect 19843 21944 19855 21947
rect 20717 21947 20775 21953
rect 20717 21944 20729 21947
rect 19843 21916 20729 21944
rect 19843 21913 19855 21916
rect 19797 21907 19855 21913
rect 20717 21913 20729 21916
rect 20763 21913 20775 21947
rect 20717 21907 20775 21913
rect 3108 21848 6914 21876
rect 3108 21836 3114 21848
rect 17310 21836 17316 21888
rect 17368 21876 17374 21888
rect 17586 21876 17592 21888
rect 17368 21848 17592 21876
rect 17368 21836 17374 21848
rect 17586 21836 17592 21848
rect 17644 21836 17650 21888
rect 20346 21876 20352 21888
rect 20307 21848 20352 21876
rect 20346 21836 20352 21848
rect 20404 21836 20410 21888
rect 22922 21876 22928 21888
rect 22883 21848 22928 21876
rect 22922 21836 22928 21848
rect 22980 21836 22986 21888
rect 23569 21879 23627 21885
rect 23569 21845 23581 21879
rect 23615 21876 23627 21879
rect 24762 21876 24768 21888
rect 23615 21848 24768 21876
rect 23615 21845 23627 21848
rect 23569 21839 23627 21845
rect 24762 21836 24768 21848
rect 24820 21836 24826 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 5350 21632 5356 21684
rect 5408 21672 5414 21684
rect 6917 21675 6975 21681
rect 6917 21672 6929 21675
rect 5408 21644 6929 21672
rect 5408 21632 5414 21644
rect 6917 21641 6929 21644
rect 6963 21641 6975 21675
rect 6917 21635 6975 21641
rect 1949 21539 2007 21545
rect 1949 21505 1961 21539
rect 1995 21536 2007 21539
rect 4062 21536 4068 21548
rect 1995 21508 4068 21536
rect 1995 21505 2007 21508
rect 1949 21499 2007 21505
rect 4062 21496 4068 21508
rect 4120 21496 4126 21548
rect 20346 21496 20352 21548
rect 20404 21536 20410 21548
rect 20441 21539 20499 21545
rect 20441 21536 20453 21539
rect 20404 21508 20453 21536
rect 20404 21496 20410 21508
rect 20441 21505 20453 21508
rect 20487 21505 20499 21539
rect 20441 21499 20499 21505
rect 37829 21539 37887 21545
rect 37829 21505 37841 21539
rect 37875 21536 37887 21539
rect 37918 21536 37924 21548
rect 37875 21508 37924 21536
rect 37875 21505 37887 21508
rect 37829 21499 37887 21505
rect 37918 21496 37924 21508
rect 37976 21496 37982 21548
rect 2038 21428 2044 21480
rect 2096 21468 2102 21480
rect 2225 21471 2283 21477
rect 2225 21468 2237 21471
rect 2096 21440 2237 21468
rect 2096 21428 2102 21440
rect 2225 21437 2237 21440
rect 2271 21437 2283 21471
rect 2225 21431 2283 21437
rect 17586 21360 17592 21412
rect 17644 21400 17650 21412
rect 21082 21400 21088 21412
rect 17644 21372 21088 21400
rect 17644 21360 17650 21372
rect 21082 21360 21088 21372
rect 21140 21400 21146 21412
rect 21140 21372 21312 21400
rect 21140 21360 21146 21372
rect 20530 21292 20536 21344
rect 20588 21332 20594 21344
rect 21284 21341 21312 21372
rect 24302 21360 24308 21412
rect 24360 21400 24366 21412
rect 37274 21400 37280 21412
rect 24360 21372 37280 21400
rect 24360 21360 24366 21372
rect 37274 21360 37280 21372
rect 37332 21360 37338 21412
rect 20625 21335 20683 21341
rect 20625 21332 20637 21335
rect 20588 21304 20637 21332
rect 20588 21292 20594 21304
rect 20625 21301 20637 21304
rect 20671 21301 20683 21335
rect 20625 21295 20683 21301
rect 21269 21335 21327 21341
rect 21269 21301 21281 21335
rect 21315 21332 21327 21335
rect 21726 21332 21732 21344
rect 21315 21304 21732 21332
rect 21315 21301 21327 21304
rect 21269 21295 21327 21301
rect 21726 21292 21732 21304
rect 21784 21292 21790 21344
rect 38010 21332 38016 21344
rect 37971 21304 38016 21332
rect 38010 21292 38016 21304
rect 38068 21292 38074 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 2038 21128 2044 21140
rect 1999 21100 2044 21128
rect 2038 21088 2044 21100
rect 2096 21088 2102 21140
rect 37826 21088 37832 21140
rect 37884 21128 37890 21140
rect 37921 21131 37979 21137
rect 37921 21128 37933 21131
rect 37884 21100 37933 21128
rect 37884 21088 37890 21100
rect 37921 21097 37933 21100
rect 37967 21097 37979 21131
rect 37921 21091 37979 21097
rect 5350 20952 5356 21004
rect 5408 20992 5414 21004
rect 6181 20995 6239 21001
rect 6181 20992 6193 20995
rect 5408 20964 6193 20992
rect 5408 20952 5414 20964
rect 6181 20961 6193 20964
rect 6227 20961 6239 20995
rect 6181 20955 6239 20961
rect 37274 20952 37280 21004
rect 37332 20992 37338 21004
rect 37826 20992 37832 21004
rect 37332 20964 37832 20992
rect 37332 20952 37338 20964
rect 37826 20952 37832 20964
rect 37884 20952 37890 21004
rect 1394 20924 1400 20936
rect 1355 20896 1400 20924
rect 1394 20884 1400 20896
rect 1452 20884 1458 20936
rect 6454 20924 6460 20936
rect 6415 20896 6460 20924
rect 6454 20884 6460 20896
rect 6512 20884 6518 20936
rect 37461 20927 37519 20933
rect 37461 20893 37473 20927
rect 37507 20924 37519 20927
rect 38102 20924 38108 20936
rect 37507 20896 38108 20924
rect 37507 20893 37519 20896
rect 37461 20887 37519 20893
rect 38102 20884 38108 20896
rect 38160 20884 38166 20936
rect 6365 20859 6423 20865
rect 6365 20856 6377 20859
rect 1596 20828 6377 20856
rect 1596 20797 1624 20828
rect 6365 20825 6377 20828
rect 6411 20825 6423 20859
rect 7377 20859 7435 20865
rect 7377 20856 7389 20859
rect 6365 20819 6423 20825
rect 6840 20828 7389 20856
rect 6840 20797 6868 20828
rect 7377 20825 7389 20828
rect 7423 20825 7435 20859
rect 7377 20819 7435 20825
rect 1581 20791 1639 20797
rect 1581 20757 1593 20791
rect 1627 20757 1639 20791
rect 1581 20751 1639 20757
rect 6825 20791 6883 20797
rect 6825 20757 6837 20791
rect 6871 20757 6883 20791
rect 7466 20788 7472 20800
rect 7427 20760 7472 20788
rect 6825 20751 6883 20757
rect 7466 20748 7472 20760
rect 7524 20748 7530 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 6454 20544 6460 20596
rect 6512 20584 6518 20596
rect 7101 20587 7159 20593
rect 7101 20584 7113 20587
rect 6512 20556 7113 20584
rect 6512 20544 6518 20556
rect 7101 20553 7113 20556
rect 7147 20553 7159 20587
rect 7101 20547 7159 20553
rect 32953 20587 33011 20593
rect 32953 20553 32965 20587
rect 32999 20584 33011 20587
rect 33410 20584 33416 20596
rect 32999 20556 33416 20584
rect 32999 20553 33011 20556
rect 32953 20547 33011 20553
rect 33410 20544 33416 20556
rect 33468 20544 33474 20596
rect 1394 20516 1400 20528
rect 1355 20488 1400 20516
rect 1394 20476 1400 20488
rect 1452 20476 1458 20528
rect 1578 20408 1584 20460
rect 1636 20448 1642 20460
rect 3237 20451 3295 20457
rect 3237 20448 3249 20451
rect 1636 20420 3249 20448
rect 1636 20408 1642 20420
rect 3237 20417 3249 20420
rect 3283 20417 3295 20451
rect 3237 20411 3295 20417
rect 33873 20451 33931 20457
rect 33873 20417 33885 20451
rect 33919 20448 33931 20451
rect 36262 20448 36268 20460
rect 33919 20420 36268 20448
rect 33919 20417 33931 20420
rect 33873 20411 33931 20417
rect 36262 20408 36268 20420
rect 36320 20408 36326 20460
rect 3329 20383 3387 20389
rect 3329 20349 3341 20383
rect 3375 20349 3387 20383
rect 3510 20380 3516 20392
rect 3471 20352 3516 20380
rect 3329 20343 3387 20349
rect 3344 20312 3372 20343
rect 3510 20340 3516 20352
rect 3568 20340 3574 20392
rect 33597 20383 33655 20389
rect 33597 20349 33609 20383
rect 33643 20380 33655 20383
rect 33778 20380 33784 20392
rect 33643 20352 33784 20380
rect 33643 20349 33655 20352
rect 33597 20343 33655 20349
rect 33778 20340 33784 20352
rect 33836 20340 33842 20392
rect 4157 20315 4215 20321
rect 4157 20312 4169 20315
rect 3344 20284 4169 20312
rect 4157 20281 4169 20284
rect 4203 20312 4215 20315
rect 32582 20312 32588 20324
rect 4203 20284 32588 20312
rect 4203 20281 4215 20284
rect 4157 20275 4215 20281
rect 32582 20272 32588 20284
rect 32640 20272 32646 20324
rect 2041 20247 2099 20253
rect 2041 20213 2053 20247
rect 2087 20244 2099 20247
rect 2222 20244 2228 20256
rect 2087 20216 2228 20244
rect 2087 20213 2099 20216
rect 2041 20207 2099 20213
rect 2222 20204 2228 20216
rect 2280 20204 2286 20256
rect 2866 20244 2872 20256
rect 2827 20216 2872 20244
rect 2866 20204 2872 20216
rect 2924 20204 2930 20256
rect 12529 20247 12587 20253
rect 12529 20213 12541 20247
rect 12575 20244 12587 20247
rect 12802 20244 12808 20256
rect 12575 20216 12808 20244
rect 12575 20213 12587 20216
rect 12529 20207 12587 20213
rect 12802 20204 12808 20216
rect 12860 20204 12866 20256
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 3510 20000 3516 20052
rect 3568 20040 3574 20052
rect 3881 20043 3939 20049
rect 3881 20040 3893 20043
rect 3568 20012 3893 20040
rect 3568 20000 3574 20012
rect 3881 20009 3893 20012
rect 3927 20040 3939 20043
rect 5350 20040 5356 20052
rect 3927 20012 5356 20040
rect 3927 20009 3939 20012
rect 3881 20003 3939 20009
rect 5350 20000 5356 20012
rect 5408 20000 5414 20052
rect 12250 20040 12256 20052
rect 12211 20012 12256 20040
rect 12250 20000 12256 20012
rect 12308 20040 12314 20052
rect 13170 20040 13176 20052
rect 12308 20012 13176 20040
rect 12308 20000 12314 20012
rect 13170 20000 13176 20012
rect 13228 20000 13234 20052
rect 14185 20043 14243 20049
rect 14185 20009 14197 20043
rect 14231 20040 14243 20043
rect 14550 20040 14556 20052
rect 14231 20012 14556 20040
rect 14231 20009 14243 20012
rect 14185 20003 14243 20009
rect 14550 20000 14556 20012
rect 14608 20000 14614 20052
rect 21821 20043 21879 20049
rect 21821 20009 21833 20043
rect 21867 20040 21879 20043
rect 21910 20040 21916 20052
rect 21867 20012 21916 20040
rect 21867 20009 21879 20012
rect 21821 20003 21879 20009
rect 21910 20000 21916 20012
rect 21968 20000 21974 20052
rect 5442 19932 5448 19984
rect 5500 19972 5506 19984
rect 37277 19975 37335 19981
rect 37277 19972 37289 19975
rect 5500 19944 37289 19972
rect 5500 19932 5506 19944
rect 37277 19941 37289 19944
rect 37323 19941 37335 19975
rect 37277 19935 37335 19941
rect 13449 19907 13507 19913
rect 13449 19873 13461 19907
rect 13495 19904 13507 19907
rect 14550 19904 14556 19916
rect 13495 19876 14556 19904
rect 13495 19873 13507 19876
rect 13449 19867 13507 19873
rect 14550 19864 14556 19876
rect 14608 19864 14614 19916
rect 15764 19876 31754 19904
rect 1946 19836 1952 19848
rect 1907 19808 1952 19836
rect 1946 19796 1952 19808
rect 2004 19796 2010 19848
rect 2222 19836 2228 19848
rect 2183 19808 2228 19836
rect 2222 19796 2228 19808
rect 2280 19796 2286 19848
rect 2866 19836 2872 19848
rect 2827 19808 2872 19836
rect 2866 19796 2872 19808
rect 2924 19796 2930 19848
rect 12802 19796 12808 19848
rect 12860 19836 12866 19848
rect 13265 19839 13323 19845
rect 13265 19836 13277 19839
rect 12860 19808 13277 19836
rect 12860 19796 12866 19808
rect 13265 19805 13277 19808
rect 13311 19805 13323 19839
rect 13265 19799 13323 19805
rect 2590 19728 2596 19780
rect 2648 19768 2654 19780
rect 15764 19768 15792 19876
rect 22922 19836 22928 19848
rect 2648 19740 15792 19768
rect 15948 19808 22928 19836
rect 2648 19728 2654 19740
rect 1670 19660 1676 19712
rect 1728 19700 1734 19712
rect 2685 19703 2743 19709
rect 2685 19700 2697 19703
rect 1728 19672 2697 19700
rect 1728 19660 1734 19672
rect 2685 19669 2697 19672
rect 2731 19669 2743 19703
rect 2685 19663 2743 19669
rect 12710 19660 12716 19712
rect 12768 19700 12774 19712
rect 12805 19703 12863 19709
rect 12805 19700 12817 19703
rect 12768 19672 12817 19700
rect 12768 19660 12774 19672
rect 12805 19669 12817 19672
rect 12851 19669 12863 19703
rect 13170 19700 13176 19712
rect 13083 19672 13176 19700
rect 12805 19663 12863 19669
rect 13170 19660 13176 19672
rect 13228 19700 13234 19712
rect 15948 19700 15976 19808
rect 22922 19796 22928 19808
rect 22980 19796 22986 19848
rect 31726 19768 31754 19876
rect 33134 19864 33140 19916
rect 33192 19904 33198 19916
rect 33229 19907 33287 19913
rect 33229 19904 33241 19907
rect 33192 19876 33241 19904
rect 33192 19864 33198 19876
rect 33229 19873 33241 19876
rect 33275 19904 33287 19907
rect 33410 19904 33416 19916
rect 33275 19876 33416 19904
rect 33275 19873 33287 19876
rect 33229 19867 33287 19873
rect 33410 19864 33416 19876
rect 33468 19864 33474 19916
rect 33321 19839 33379 19845
rect 33321 19805 33333 19839
rect 33367 19836 33379 19839
rect 35434 19836 35440 19848
rect 33367 19808 35440 19836
rect 33367 19805 33379 19808
rect 33321 19799 33379 19805
rect 35434 19796 35440 19808
rect 35492 19796 35498 19848
rect 37292 19836 37320 19935
rect 37829 19839 37887 19845
rect 37829 19836 37841 19839
rect 37292 19808 37841 19836
rect 37829 19805 37841 19808
rect 37875 19805 37887 19839
rect 37829 19799 37887 19805
rect 32493 19771 32551 19777
rect 32493 19768 32505 19771
rect 31726 19740 32505 19768
rect 32493 19737 32505 19740
rect 32539 19768 32551 19771
rect 33413 19771 33471 19777
rect 33413 19768 33425 19771
rect 32539 19740 33425 19768
rect 32539 19737 32551 19740
rect 32493 19731 32551 19737
rect 33413 19737 33425 19740
rect 33459 19737 33471 19771
rect 33413 19731 33471 19737
rect 13228 19672 15976 19700
rect 33781 19703 33839 19709
rect 13228 19660 13234 19672
rect 33781 19669 33793 19703
rect 33827 19700 33839 19703
rect 34238 19700 34244 19712
rect 33827 19672 34244 19700
rect 33827 19669 33839 19672
rect 33781 19663 33839 19669
rect 34238 19660 34244 19672
rect 34296 19660 34302 19712
rect 38010 19700 38016 19712
rect 37971 19672 38016 19700
rect 38010 19660 38016 19672
rect 38068 19660 38074 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 3326 19496 3332 19508
rect 3287 19468 3332 19496
rect 3326 19456 3332 19468
rect 3384 19456 3390 19508
rect 33778 19496 33784 19508
rect 33739 19468 33784 19496
rect 33778 19456 33784 19468
rect 33836 19456 33842 19508
rect 23109 19431 23167 19437
rect 23109 19428 23121 19431
rect 22296 19400 23121 19428
rect 22296 19372 22324 19400
rect 23109 19397 23121 19400
rect 23155 19397 23167 19431
rect 23109 19391 23167 19397
rect 1670 19360 1676 19372
rect 1631 19332 1676 19360
rect 1670 19320 1676 19332
rect 1728 19320 1734 19372
rect 3510 19360 3516 19372
rect 3471 19332 3516 19360
rect 3510 19320 3516 19332
rect 3568 19320 3574 19372
rect 12710 19360 12716 19372
rect 12671 19332 12716 19360
rect 12710 19320 12716 19332
rect 12768 19320 12774 19372
rect 22278 19360 22284 19372
rect 22239 19332 22284 19360
rect 22278 19320 22284 19332
rect 22336 19320 22342 19372
rect 22373 19363 22431 19369
rect 22373 19329 22385 19363
rect 22419 19360 22431 19363
rect 23750 19360 23756 19372
rect 22419 19332 23756 19360
rect 22419 19329 22431 19332
rect 22373 19323 22431 19329
rect 23750 19320 23756 19332
rect 23808 19320 23814 19372
rect 33413 19363 33471 19369
rect 33413 19329 33425 19363
rect 33459 19329 33471 19363
rect 34238 19360 34244 19372
rect 34199 19332 34244 19360
rect 33413 19323 33471 19329
rect 21910 19252 21916 19304
rect 21968 19292 21974 19304
rect 22465 19295 22523 19301
rect 22465 19292 22477 19295
rect 21968 19264 22477 19292
rect 21968 19252 21974 19264
rect 22465 19261 22477 19264
rect 22511 19261 22523 19295
rect 33134 19292 33140 19304
rect 33095 19264 33140 19292
rect 22465 19255 22523 19261
rect 33134 19252 33140 19264
rect 33192 19252 33198 19304
rect 33318 19292 33324 19304
rect 33279 19264 33324 19292
rect 33318 19252 33324 19264
rect 33376 19252 33382 19304
rect 32493 19227 32551 19233
rect 32493 19224 32505 19227
rect 6886 19196 32505 19224
rect 1486 19156 1492 19168
rect 1447 19128 1492 19156
rect 1486 19116 1492 19128
rect 1544 19116 1550 19168
rect 1946 19116 1952 19168
rect 2004 19156 2010 19168
rect 6886 19156 6914 19196
rect 32493 19193 32505 19196
rect 32539 19224 32551 19227
rect 33428 19224 33456 19323
rect 34238 19320 34244 19332
rect 34296 19320 34302 19372
rect 32539 19196 33456 19224
rect 32539 19193 32551 19196
rect 32493 19187 32551 19193
rect 12526 19156 12532 19168
rect 2004 19128 6914 19156
rect 12487 19128 12532 19156
rect 2004 19116 2010 19128
rect 12526 19116 12532 19128
rect 12584 19116 12590 19168
rect 21910 19156 21916 19168
rect 21871 19128 21916 19156
rect 21910 19116 21916 19128
rect 21968 19116 21974 19168
rect 23750 19156 23756 19168
rect 23711 19128 23756 19156
rect 23750 19116 23756 19128
rect 23808 19116 23814 19168
rect 34425 19159 34483 19165
rect 34425 19125 34437 19159
rect 34471 19156 34483 19159
rect 35342 19156 35348 19168
rect 34471 19128 35348 19156
rect 34471 19125 34483 19128
rect 34425 19119 34483 19125
rect 35342 19116 35348 19128
rect 35400 19116 35406 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 32953 18955 33011 18961
rect 32953 18921 32965 18955
rect 32999 18952 33011 18955
rect 33134 18952 33140 18964
rect 32999 18924 33140 18952
rect 32999 18921 33011 18924
rect 32953 18915 33011 18921
rect 33134 18912 33140 18924
rect 33192 18912 33198 18964
rect 10410 18776 10416 18828
rect 10468 18816 10474 18828
rect 21361 18819 21419 18825
rect 10468 18788 17080 18816
rect 10468 18776 10474 18788
rect 1673 18751 1731 18757
rect 1673 18717 1685 18751
rect 1719 18748 1731 18751
rect 12526 18748 12532 18760
rect 1719 18720 12532 18748
rect 1719 18717 1731 18720
rect 1673 18711 1731 18717
rect 12526 18708 12532 18720
rect 12584 18708 12590 18760
rect 17052 18748 17080 18788
rect 21361 18785 21373 18819
rect 21407 18816 21419 18819
rect 21910 18816 21916 18828
rect 21407 18788 21916 18816
rect 21407 18785 21419 18788
rect 21361 18779 21419 18785
rect 21910 18776 21916 18788
rect 21968 18776 21974 18828
rect 21637 18751 21695 18757
rect 21637 18748 21649 18751
rect 17052 18720 21649 18748
rect 21637 18717 21649 18720
rect 21683 18717 21695 18751
rect 21637 18711 21695 18717
rect 35342 18708 35348 18760
rect 35400 18748 35406 18760
rect 37829 18751 37887 18757
rect 37829 18748 37841 18751
rect 35400 18720 37841 18748
rect 35400 18708 35406 18720
rect 37829 18717 37841 18720
rect 37875 18717 37887 18751
rect 37829 18711 37887 18717
rect 1486 18612 1492 18624
rect 1447 18584 1492 18612
rect 1486 18572 1492 18584
rect 1544 18572 1550 18624
rect 9122 18572 9128 18624
rect 9180 18612 9186 18624
rect 26050 18612 26056 18624
rect 9180 18584 26056 18612
rect 9180 18572 9186 18584
rect 26050 18572 26056 18584
rect 26108 18572 26114 18624
rect 33318 18572 33324 18624
rect 33376 18612 33382 18624
rect 33873 18615 33931 18621
rect 33873 18612 33885 18615
rect 33376 18584 33885 18612
rect 33376 18572 33382 18584
rect 33873 18581 33885 18584
rect 33919 18581 33931 18615
rect 38010 18612 38016 18624
rect 37971 18584 38016 18612
rect 33873 18575 33931 18581
rect 38010 18572 38016 18584
rect 38068 18572 38074 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 14274 18408 14280 18420
rect 14235 18380 14280 18408
rect 14274 18368 14280 18380
rect 14332 18368 14338 18420
rect 22462 18368 22468 18420
rect 22520 18408 22526 18420
rect 25133 18411 25191 18417
rect 25133 18408 25145 18411
rect 22520 18380 25145 18408
rect 22520 18368 22526 18380
rect 25133 18377 25145 18380
rect 25179 18377 25191 18411
rect 25133 18371 25191 18377
rect 2225 18343 2283 18349
rect 2225 18340 2237 18343
rect 1688 18312 2237 18340
rect 1688 18281 1716 18312
rect 2225 18309 2237 18312
rect 2271 18340 2283 18343
rect 22646 18340 22652 18352
rect 2271 18312 22652 18340
rect 2271 18309 2283 18312
rect 2225 18303 2283 18309
rect 22646 18300 22652 18312
rect 22704 18300 22710 18352
rect 1673 18275 1731 18281
rect 1673 18241 1685 18275
rect 1719 18241 1731 18275
rect 12986 18272 12992 18284
rect 12947 18244 12992 18272
rect 1673 18235 1731 18241
rect 12986 18232 12992 18244
rect 13044 18232 13050 18284
rect 25148 18204 25176 18371
rect 26053 18275 26111 18281
rect 26053 18272 26065 18275
rect 25884 18244 26065 18272
rect 25777 18207 25835 18213
rect 25777 18204 25789 18207
rect 25148 18176 25789 18204
rect 25777 18173 25789 18176
rect 25823 18173 25835 18207
rect 25777 18167 25835 18173
rect 24578 18096 24584 18148
rect 24636 18136 24642 18148
rect 25884 18136 25912 18244
rect 26053 18241 26065 18244
rect 26099 18272 26111 18275
rect 26973 18275 27031 18281
rect 26973 18272 26985 18275
rect 26099 18244 26985 18272
rect 26099 18241 26111 18244
rect 26053 18235 26111 18241
rect 26973 18241 26985 18244
rect 27019 18241 27031 18275
rect 26973 18235 27031 18241
rect 37461 18275 37519 18281
rect 37461 18241 37473 18275
rect 37507 18272 37519 18275
rect 38102 18272 38108 18284
rect 37507 18244 38108 18272
rect 37507 18241 37519 18244
rect 37461 18235 37519 18241
rect 38102 18232 38108 18244
rect 38160 18232 38166 18284
rect 25961 18207 26019 18213
rect 25961 18173 25973 18207
rect 26007 18204 26019 18207
rect 26007 18176 35894 18204
rect 26007 18173 26019 18176
rect 25961 18167 26019 18173
rect 33778 18136 33784 18148
rect 24636 18108 33784 18136
rect 24636 18096 24642 18108
rect 33778 18096 33784 18108
rect 33836 18096 33842 18148
rect 35866 18136 35894 18176
rect 37921 18139 37979 18145
rect 37921 18136 37933 18139
rect 35866 18108 37933 18136
rect 37921 18105 37933 18108
rect 37967 18105 37979 18139
rect 37921 18099 37979 18105
rect 1486 18068 1492 18080
rect 1447 18040 1492 18068
rect 1486 18028 1492 18040
rect 1544 18028 1550 18080
rect 26421 18071 26479 18077
rect 26421 18037 26433 18071
rect 26467 18068 26479 18071
rect 26510 18068 26516 18080
rect 26467 18040 26516 18068
rect 26467 18037 26479 18040
rect 26421 18031 26479 18037
rect 26510 18028 26516 18040
rect 26568 18028 26574 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 3510 17824 3516 17876
rect 3568 17864 3574 17876
rect 3789 17867 3847 17873
rect 3789 17864 3801 17867
rect 3568 17836 3801 17864
rect 3568 17824 3574 17836
rect 3789 17833 3801 17836
rect 3835 17833 3847 17867
rect 3789 17827 3847 17833
rect 12986 17756 12992 17808
rect 13044 17796 13050 17808
rect 16025 17799 16083 17805
rect 16025 17796 16037 17799
rect 13044 17768 16037 17796
rect 13044 17756 13050 17768
rect 16025 17765 16037 17768
rect 16071 17765 16083 17799
rect 16025 17759 16083 17765
rect 4433 17731 4491 17737
rect 4433 17697 4445 17731
rect 4479 17728 4491 17731
rect 4614 17728 4620 17740
rect 4479 17700 4620 17728
rect 4479 17697 4491 17700
rect 4433 17691 4491 17697
rect 4614 17688 4620 17700
rect 4672 17688 4678 17740
rect 8018 17620 8024 17672
rect 8076 17660 8082 17672
rect 21818 17660 21824 17672
rect 8076 17632 21824 17660
rect 8076 17620 8082 17632
rect 21818 17620 21824 17632
rect 21876 17620 21882 17672
rect 26510 17660 26516 17672
rect 26471 17632 26516 17660
rect 26510 17620 26516 17632
rect 26568 17620 26574 17672
rect 36725 17663 36783 17669
rect 36725 17629 36737 17663
rect 36771 17660 36783 17663
rect 38102 17660 38108 17672
rect 36771 17632 38108 17660
rect 36771 17629 36783 17632
rect 36725 17623 36783 17629
rect 38102 17620 38108 17632
rect 38160 17620 38166 17672
rect 14737 17595 14795 17601
rect 14737 17561 14749 17595
rect 14783 17561 14795 17595
rect 14737 17555 14795 17561
rect 1578 17484 1584 17536
rect 1636 17524 1642 17536
rect 4157 17527 4215 17533
rect 4157 17524 4169 17527
rect 1636 17496 4169 17524
rect 1636 17484 1642 17496
rect 4157 17493 4169 17496
rect 4203 17493 4215 17527
rect 4157 17487 4215 17493
rect 4249 17527 4307 17533
rect 4249 17493 4261 17527
rect 4295 17524 4307 17527
rect 4890 17524 4896 17536
rect 4295 17496 4896 17524
rect 4295 17493 4307 17496
rect 4249 17487 4307 17493
rect 4890 17484 4896 17496
rect 4948 17524 4954 17536
rect 4985 17527 5043 17533
rect 4985 17524 4997 17527
rect 4948 17496 4997 17524
rect 4948 17484 4954 17496
rect 4985 17493 4997 17496
rect 5031 17493 5043 17527
rect 4985 17487 5043 17493
rect 10318 17484 10324 17536
rect 10376 17524 10382 17536
rect 14185 17527 14243 17533
rect 14185 17524 14197 17527
rect 10376 17496 14197 17524
rect 10376 17484 10382 17496
rect 14185 17493 14197 17496
rect 14231 17524 14243 17527
rect 14752 17524 14780 17555
rect 14231 17496 14780 17524
rect 26697 17527 26755 17533
rect 14231 17493 14243 17496
rect 14185 17487 14243 17493
rect 26697 17493 26709 17527
rect 26743 17524 26755 17527
rect 33870 17524 33876 17536
rect 26743 17496 33876 17524
rect 26743 17493 26755 17496
rect 26697 17487 26755 17493
rect 33870 17484 33876 17496
rect 33928 17484 33934 17536
rect 37274 17524 37280 17536
rect 37235 17496 37280 17524
rect 37274 17484 37280 17496
rect 37332 17484 37338 17536
rect 37642 17484 37648 17536
rect 37700 17524 37706 17536
rect 37921 17527 37979 17533
rect 37921 17524 37933 17527
rect 37700 17496 37933 17524
rect 37700 17484 37706 17496
rect 37921 17493 37933 17496
rect 37967 17493 37979 17527
rect 37921 17487 37979 17493
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 1578 17320 1584 17332
rect 1539 17292 1584 17320
rect 1578 17280 1584 17292
rect 1636 17280 1642 17332
rect 4614 17320 4620 17332
rect 4575 17292 4620 17320
rect 4614 17280 4620 17292
rect 4672 17280 4678 17332
rect 21174 17280 21180 17332
rect 21232 17320 21238 17332
rect 35802 17320 35808 17332
rect 21232 17292 35808 17320
rect 21232 17280 21238 17292
rect 35802 17280 35808 17292
rect 35860 17280 35866 17332
rect 37642 17320 37648 17332
rect 37603 17292 37648 17320
rect 37642 17280 37648 17292
rect 37700 17280 37706 17332
rect 37734 17280 37740 17332
rect 37792 17320 37798 17332
rect 37792 17292 37837 17320
rect 37792 17280 37798 17292
rect 21266 17212 21272 17264
rect 21324 17252 21330 17264
rect 36725 17255 36783 17261
rect 21324 17224 22094 17252
rect 21324 17212 21330 17224
rect 1394 17184 1400 17196
rect 1355 17156 1400 17184
rect 1394 17144 1400 17156
rect 1452 17184 1458 17196
rect 2041 17187 2099 17193
rect 2041 17184 2053 17187
rect 1452 17156 2053 17184
rect 1452 17144 1458 17156
rect 2041 17153 2053 17156
rect 2087 17153 2099 17187
rect 22066 17184 22094 17224
rect 36725 17221 36737 17255
rect 36771 17252 36783 17255
rect 37752 17252 37780 17280
rect 36771 17224 37780 17252
rect 36771 17221 36783 17224
rect 36725 17215 36783 17221
rect 37642 17184 37648 17196
rect 22066 17156 37648 17184
rect 2041 17147 2099 17153
rect 37642 17144 37648 17156
rect 37700 17144 37706 17196
rect 26970 17076 26976 17128
rect 27028 17116 27034 17128
rect 37274 17116 37280 17128
rect 27028 17088 37280 17116
rect 27028 17076 27034 17088
rect 37274 17076 37280 17088
rect 37332 17116 37338 17128
rect 37461 17119 37519 17125
rect 37461 17116 37473 17119
rect 37332 17088 37473 17116
rect 37332 17076 37338 17088
rect 37461 17085 37473 17088
rect 37507 17085 37519 17119
rect 37461 17079 37519 17085
rect 1946 16940 1952 16992
rect 2004 16980 2010 16992
rect 8202 16980 8208 16992
rect 2004 16952 8208 16980
rect 2004 16940 2010 16952
rect 8202 16940 8208 16952
rect 8260 16940 8266 16992
rect 38010 16940 38016 16992
rect 38068 16980 38074 16992
rect 38105 16983 38163 16989
rect 38105 16980 38117 16983
rect 38068 16952 38117 16980
rect 38068 16940 38074 16952
rect 38105 16949 38117 16952
rect 38151 16949 38163 16983
rect 38105 16943 38163 16949
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 18046 16708 18052 16720
rect 1964 16680 18052 16708
rect 1964 16649 1992 16680
rect 18046 16668 18052 16680
rect 18104 16668 18110 16720
rect 25148 16680 26004 16708
rect 1949 16643 2007 16649
rect 1949 16609 1961 16643
rect 1995 16609 2007 16643
rect 1949 16603 2007 16609
rect 4062 16600 4068 16652
rect 4120 16640 4126 16652
rect 25148 16649 25176 16680
rect 25976 16649 26004 16680
rect 25133 16643 25191 16649
rect 25133 16640 25145 16643
rect 4120 16612 25145 16640
rect 4120 16600 4126 16612
rect 25133 16609 25145 16612
rect 25179 16609 25191 16643
rect 25133 16603 25191 16609
rect 25869 16643 25927 16649
rect 25869 16609 25881 16643
rect 25915 16609 25927 16643
rect 25869 16603 25927 16609
rect 25961 16643 26019 16649
rect 25961 16609 25973 16643
rect 26007 16609 26019 16643
rect 25961 16603 26019 16609
rect 36725 16643 36783 16649
rect 36725 16609 36737 16643
rect 36771 16609 36783 16643
rect 36725 16603 36783 16609
rect 2038 16532 2044 16584
rect 2096 16572 2102 16584
rect 2225 16575 2283 16581
rect 2225 16572 2237 16575
rect 2096 16544 2237 16572
rect 2096 16532 2102 16544
rect 2225 16541 2237 16544
rect 2271 16541 2283 16575
rect 25884 16572 25912 16603
rect 26142 16572 26148 16584
rect 25884 16544 26148 16572
rect 2225 16535 2283 16541
rect 26142 16532 26148 16544
rect 26200 16532 26206 16584
rect 26881 16575 26939 16581
rect 26881 16572 26893 16575
rect 26436 16544 26893 16572
rect 26053 16439 26111 16445
rect 26053 16405 26065 16439
rect 26099 16436 26111 16439
rect 26326 16436 26332 16448
rect 26099 16408 26332 16436
rect 26099 16405 26111 16408
rect 26053 16399 26111 16405
rect 26326 16396 26332 16408
rect 26384 16396 26390 16448
rect 26436 16445 26464 16544
rect 26881 16541 26893 16544
rect 26927 16541 26939 16575
rect 36740 16572 36768 16603
rect 37182 16572 37188 16584
rect 36740 16544 37188 16572
rect 26881 16535 26939 16541
rect 37182 16532 37188 16544
rect 37240 16572 37246 16584
rect 37369 16575 37427 16581
rect 37369 16572 37381 16575
rect 37240 16544 37381 16572
rect 37240 16532 37246 16544
rect 37369 16541 37381 16544
rect 37415 16541 37427 16575
rect 38010 16572 38016 16584
rect 37971 16544 38016 16572
rect 37369 16535 37427 16541
rect 38010 16532 38016 16544
rect 38068 16532 38074 16584
rect 26421 16439 26479 16445
rect 26421 16405 26433 16439
rect 26467 16405 26479 16439
rect 27062 16436 27068 16448
rect 27023 16408 27068 16436
rect 26421 16399 26479 16405
rect 27062 16396 27068 16408
rect 27120 16396 27126 16448
rect 35434 16396 35440 16448
rect 35492 16436 35498 16448
rect 37185 16439 37243 16445
rect 37185 16436 37197 16439
rect 35492 16408 37197 16436
rect 35492 16396 35498 16408
rect 37185 16405 37197 16408
rect 37231 16405 37243 16439
rect 37185 16399 37243 16405
rect 37734 16396 37740 16448
rect 37792 16436 37798 16448
rect 37829 16439 37887 16445
rect 37829 16436 37841 16439
rect 37792 16408 37841 16436
rect 37792 16396 37798 16408
rect 37829 16405 37841 16408
rect 37875 16405 37887 16439
rect 37829 16399 37887 16405
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 2038 16232 2044 16244
rect 1999 16204 2044 16232
rect 2038 16192 2044 16204
rect 2096 16192 2102 16244
rect 13814 16192 13820 16244
rect 13872 16232 13878 16244
rect 21634 16232 21640 16244
rect 13872 16204 21640 16232
rect 13872 16192 13878 16204
rect 21634 16192 21640 16204
rect 21692 16192 21698 16244
rect 26142 16192 26148 16244
rect 26200 16232 26206 16244
rect 26973 16235 27031 16241
rect 26973 16232 26985 16235
rect 26200 16204 26985 16232
rect 26200 16192 26206 16204
rect 26973 16201 26985 16204
rect 27019 16201 27031 16235
rect 37366 16232 37372 16244
rect 37327 16204 37372 16232
rect 26973 16195 27031 16201
rect 37366 16192 37372 16204
rect 37424 16192 37430 16244
rect 15028 16136 16068 16164
rect 1394 16096 1400 16108
rect 1355 16068 1400 16096
rect 1394 16056 1400 16068
rect 1452 16056 1458 16108
rect 15028 16096 15056 16136
rect 14936 16068 15056 16096
rect 15105 16099 15163 16105
rect 14936 16037 14964 16068
rect 15105 16065 15117 16099
rect 15151 16065 15163 16099
rect 15105 16059 15163 16065
rect 14921 16031 14979 16037
rect 14921 15997 14933 16031
rect 14967 15997 14979 16031
rect 14921 15991 14979 15997
rect 15013 16031 15071 16037
rect 15013 15997 15025 16031
rect 15059 15997 15071 16031
rect 15013 15991 15071 15997
rect 1581 15963 1639 15969
rect 1581 15929 1593 15963
rect 1627 15960 1639 15963
rect 15028 15960 15056 15991
rect 1627 15932 15056 15960
rect 1627 15929 1639 15932
rect 1581 15923 1639 15929
rect 1762 15852 1768 15904
rect 1820 15892 1826 15904
rect 14185 15895 14243 15901
rect 14185 15892 14197 15895
rect 1820 15864 14197 15892
rect 1820 15852 1826 15864
rect 14185 15861 14197 15864
rect 14231 15892 14243 15895
rect 15120 15892 15148 16059
rect 15470 15892 15476 15904
rect 14231 15864 15148 15892
rect 15431 15864 15476 15892
rect 14231 15861 14243 15864
rect 14185 15855 14243 15861
rect 15470 15852 15476 15864
rect 15528 15852 15534 15904
rect 16040 15901 16068 16136
rect 37384 16096 37412 16192
rect 37829 16099 37887 16105
rect 37829 16096 37841 16099
rect 37384 16068 37841 16096
rect 37829 16065 37841 16068
rect 37875 16065 37887 16099
rect 37829 16059 37887 16065
rect 27062 15988 27068 16040
rect 27120 16028 27126 16040
rect 38470 16028 38476 16040
rect 27120 16000 38476 16028
rect 27120 15988 27126 16000
rect 38470 15988 38476 16000
rect 38528 15988 38534 16040
rect 16025 15895 16083 15901
rect 16025 15861 16037 15895
rect 16071 15892 16083 15895
rect 21726 15892 21732 15904
rect 16071 15864 21732 15892
rect 16071 15861 16083 15864
rect 16025 15855 16083 15861
rect 21726 15852 21732 15864
rect 21784 15852 21790 15904
rect 38010 15892 38016 15904
rect 37971 15864 38016 15892
rect 38010 15852 38016 15864
rect 38068 15852 38074 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 1394 15688 1400 15700
rect 1355 15660 1400 15688
rect 1394 15648 1400 15660
rect 1452 15648 1458 15700
rect 15470 15552 15476 15564
rect 15431 15524 15476 15552
rect 15470 15512 15476 15524
rect 15528 15512 15534 15564
rect 15749 15487 15807 15493
rect 15749 15453 15761 15487
rect 15795 15484 15807 15487
rect 16298 15484 16304 15496
rect 15795 15456 16304 15484
rect 15795 15453 15807 15456
rect 15749 15447 15807 15453
rect 16298 15444 16304 15456
rect 16356 15444 16362 15496
rect 37461 15487 37519 15493
rect 37461 15453 37473 15487
rect 37507 15484 37519 15487
rect 38102 15484 38108 15496
rect 37507 15456 38108 15484
rect 37507 15453 37519 15456
rect 37461 15447 37519 15453
rect 38102 15444 38108 15456
rect 38160 15444 38166 15496
rect 26326 15308 26332 15360
rect 26384 15348 26390 15360
rect 26970 15348 26976 15360
rect 26384 15320 26976 15348
rect 26384 15308 26390 15320
rect 26970 15308 26976 15320
rect 27028 15308 27034 15360
rect 37918 15348 37924 15360
rect 37879 15320 37924 15348
rect 37918 15308 37924 15320
rect 37976 15308 37982 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 1762 15104 1768 15156
rect 1820 15144 1826 15156
rect 4798 15144 4804 15156
rect 1820 15116 4804 15144
rect 1820 15104 1826 15116
rect 4798 15104 4804 15116
rect 4856 15104 4862 15156
rect 27062 15104 27068 15156
rect 27120 15144 27126 15156
rect 27341 15147 27399 15153
rect 27341 15144 27353 15147
rect 27120 15116 27353 15144
rect 27120 15104 27126 15116
rect 27341 15113 27353 15116
rect 27387 15113 27399 15147
rect 27341 15107 27399 15113
rect 34793 15147 34851 15153
rect 34793 15113 34805 15147
rect 34839 15144 34851 15147
rect 38010 15144 38016 15156
rect 34839 15116 38016 15144
rect 34839 15113 34851 15116
rect 34793 15107 34851 15113
rect 4798 15008 4804 15020
rect 4759 14980 4804 15008
rect 4798 14968 4804 14980
rect 4856 14968 4862 15020
rect 27356 15008 27384 15107
rect 38010 15104 38016 15116
rect 38068 15104 38074 15156
rect 28261 15079 28319 15085
rect 28261 15045 28273 15079
rect 28307 15076 28319 15079
rect 37918 15076 37924 15088
rect 28307 15048 37924 15076
rect 28307 15045 28319 15048
rect 28261 15039 28319 15045
rect 37918 15036 37924 15048
rect 37976 15036 37982 15088
rect 34606 15008 34612 15020
rect 27356 14980 28488 15008
rect 34567 14980 34612 15008
rect 28350 14940 28356 14952
rect 28311 14912 28356 14940
rect 28350 14900 28356 14912
rect 28408 14900 28414 14952
rect 28460 14949 28488 14980
rect 34606 14968 34612 14980
rect 34664 14968 34670 15020
rect 28445 14943 28503 14949
rect 28445 14909 28457 14943
rect 28491 14909 28503 14943
rect 28445 14903 28503 14909
rect 4985 14875 5043 14881
rect 4985 14841 4997 14875
rect 5031 14872 5043 14875
rect 38562 14872 38568 14884
rect 5031 14844 38568 14872
rect 5031 14841 5043 14844
rect 4985 14835 5043 14841
rect 38562 14832 38568 14844
rect 38620 14832 38626 14884
rect 27890 14804 27896 14816
rect 27851 14776 27896 14804
rect 27890 14764 27896 14776
rect 27948 14764 27954 14816
rect 38102 14804 38108 14816
rect 38063 14776 38108 14804
rect 38102 14764 38108 14776
rect 38160 14764 38166 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 26694 14560 26700 14612
rect 26752 14600 26758 14612
rect 26789 14603 26847 14609
rect 26789 14600 26801 14603
rect 26752 14572 26801 14600
rect 26752 14560 26758 14572
rect 26789 14569 26801 14572
rect 26835 14569 26847 14603
rect 26789 14563 26847 14569
rect 27341 14467 27399 14473
rect 27341 14433 27353 14467
rect 27387 14464 27399 14467
rect 27890 14464 27896 14476
rect 27387 14436 27896 14464
rect 27387 14433 27399 14436
rect 27341 14427 27399 14433
rect 27890 14424 27896 14436
rect 27948 14424 27954 14476
rect 37826 14464 37832 14476
rect 37787 14436 37832 14464
rect 37826 14424 37832 14436
rect 37884 14424 37890 14476
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14396 1731 14399
rect 2225 14399 2283 14405
rect 2225 14396 2237 14399
rect 1719 14368 2237 14396
rect 1719 14365 1731 14368
rect 1673 14359 1731 14365
rect 2225 14365 2237 14368
rect 2271 14396 2283 14399
rect 18966 14396 18972 14408
rect 2271 14368 18972 14396
rect 2271 14365 2283 14368
rect 2225 14359 2283 14365
rect 18966 14356 18972 14368
rect 19024 14356 19030 14408
rect 27614 14396 27620 14408
rect 27575 14368 27620 14396
rect 27614 14356 27620 14368
rect 27672 14356 27678 14408
rect 38102 14396 38108 14408
rect 38063 14368 38108 14396
rect 38102 14356 38108 14368
rect 38160 14356 38166 14408
rect 1486 14260 1492 14272
rect 1447 14232 1492 14260
rect 1486 14220 1492 14232
rect 1544 14220 1550 14272
rect 24118 14220 24124 14272
rect 24176 14260 24182 14272
rect 26418 14260 26424 14272
rect 24176 14232 26424 14260
rect 24176 14220 24182 14232
rect 26418 14220 26424 14232
rect 26476 14220 26482 14272
rect 33689 14263 33747 14269
rect 33689 14229 33701 14263
rect 33735 14260 33747 14263
rect 34422 14260 34428 14272
rect 33735 14232 34428 14260
rect 33735 14229 33747 14232
rect 33689 14223 33747 14229
rect 34422 14220 34428 14232
rect 34480 14220 34486 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 4801 14059 4859 14065
rect 4801 14025 4813 14059
rect 4847 14056 4859 14059
rect 24118 14056 24124 14068
rect 4847 14028 24124 14056
rect 4847 14025 4859 14028
rect 4801 14019 4859 14025
rect 24118 14016 24124 14028
rect 24176 14016 24182 14068
rect 33229 14059 33287 14065
rect 33229 14056 33241 14059
rect 26252 14028 33241 14056
rect 9214 13948 9220 14000
rect 9272 13988 9278 14000
rect 14458 13988 14464 14000
rect 9272 13960 14464 13988
rect 9272 13948 9278 13960
rect 14458 13948 14464 13960
rect 14516 13948 14522 14000
rect 14568 13960 19334 13988
rect 1949 13923 2007 13929
rect 1949 13889 1961 13923
rect 1995 13920 2007 13923
rect 4614 13920 4620 13932
rect 1995 13892 4476 13920
rect 4575 13892 4620 13920
rect 1995 13889 2007 13892
rect 1949 13883 2007 13889
rect 2038 13812 2044 13864
rect 2096 13852 2102 13864
rect 2225 13855 2283 13861
rect 2225 13852 2237 13855
rect 2096 13824 2237 13852
rect 2096 13812 2102 13824
rect 2225 13821 2237 13824
rect 2271 13821 2283 13855
rect 4448 13852 4476 13892
rect 4614 13880 4620 13892
rect 4672 13880 4678 13932
rect 14568 13920 14596 13960
rect 6886 13892 14596 13920
rect 19306 13920 19334 13960
rect 26252 13920 26280 14028
rect 33229 14025 33241 14028
rect 33275 14056 33287 14059
rect 34149 14059 34207 14065
rect 34149 14056 34161 14059
rect 33275 14028 34161 14056
rect 33275 14025 33287 14028
rect 33229 14019 33287 14025
rect 34149 14025 34161 14028
rect 34195 14025 34207 14059
rect 34149 14019 34207 14025
rect 34241 14059 34299 14065
rect 34241 14025 34253 14059
rect 34287 14056 34299 14059
rect 34514 14056 34520 14068
rect 34287 14028 34520 14056
rect 34287 14025 34299 14028
rect 34241 14019 34299 14025
rect 34514 14016 34520 14028
rect 34572 14056 34578 14068
rect 34977 14059 35035 14065
rect 34977 14056 34989 14059
rect 34572 14028 34989 14056
rect 34572 14016 34578 14028
rect 34977 14025 34989 14028
rect 35023 14025 35035 14059
rect 34977 14019 35035 14025
rect 26418 13948 26424 14000
rect 26476 13988 26482 14000
rect 38286 13988 38292 14000
rect 26476 13960 38292 13988
rect 26476 13948 26482 13960
rect 38286 13948 38292 13960
rect 38344 13948 38350 14000
rect 27341 13923 27399 13929
rect 27341 13920 27353 13923
rect 19306 13892 26280 13920
rect 26436 13892 27353 13920
rect 6886 13852 6914 13892
rect 4448 13824 6914 13852
rect 2225 13815 2283 13821
rect 14458 13812 14464 13864
rect 14516 13852 14522 13864
rect 26329 13855 26387 13861
rect 26329 13852 26341 13855
rect 14516 13824 26341 13852
rect 14516 13812 14522 13824
rect 26329 13821 26341 13824
rect 26375 13852 26387 13855
rect 26436 13852 26464 13892
rect 27341 13889 27353 13892
rect 27387 13889 27399 13923
rect 27341 13883 27399 13889
rect 36814 13880 36820 13932
rect 36872 13920 36878 13932
rect 37829 13923 37887 13929
rect 37829 13920 37841 13923
rect 36872 13892 37841 13920
rect 36872 13880 36878 13892
rect 37829 13889 37841 13892
rect 37875 13889 37887 13923
rect 37829 13883 37887 13889
rect 27430 13852 27436 13864
rect 26375 13824 26464 13852
rect 27391 13824 27436 13852
rect 26375 13821 26387 13824
rect 26329 13815 26387 13821
rect 27430 13812 27436 13824
rect 27488 13812 27494 13864
rect 27525 13855 27583 13861
rect 27525 13821 27537 13855
rect 27571 13821 27583 13855
rect 34422 13852 34428 13864
rect 34383 13824 34428 13852
rect 27525 13815 27583 13821
rect 26234 13744 26240 13796
rect 26292 13784 26298 13796
rect 26694 13784 26700 13796
rect 26292 13756 26700 13784
rect 26292 13744 26298 13756
rect 26694 13744 26700 13756
rect 26752 13784 26758 13796
rect 27540 13784 27568 13815
rect 34422 13812 34428 13824
rect 34480 13812 34486 13864
rect 26752 13756 27568 13784
rect 26752 13744 26758 13756
rect 26878 13676 26884 13728
rect 26936 13716 26942 13728
rect 26973 13719 27031 13725
rect 26973 13716 26985 13719
rect 26936 13688 26985 13716
rect 26936 13676 26942 13688
rect 26973 13685 26985 13688
rect 27019 13685 27031 13719
rect 26973 13679 27031 13685
rect 33781 13719 33839 13725
rect 33781 13685 33793 13719
rect 33827 13716 33839 13719
rect 33962 13716 33968 13728
rect 33827 13688 33968 13716
rect 33827 13685 33839 13688
rect 33781 13679 33839 13685
rect 33962 13676 33968 13688
rect 34020 13676 34026 13728
rect 38010 13716 38016 13728
rect 37971 13688 38016 13716
rect 38010 13676 38016 13688
rect 38068 13676 38074 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 2038 13512 2044 13524
rect 1999 13484 2044 13512
rect 2038 13472 2044 13484
rect 2096 13472 2102 13524
rect 4525 13515 4583 13521
rect 4525 13481 4537 13515
rect 4571 13512 4583 13515
rect 4614 13512 4620 13524
rect 4571 13484 4620 13512
rect 4571 13481 4583 13484
rect 4525 13475 4583 13481
rect 4614 13472 4620 13484
rect 4672 13472 4678 13524
rect 34606 13472 34612 13524
rect 34664 13512 34670 13524
rect 34701 13515 34759 13521
rect 34701 13512 34713 13515
rect 34664 13484 34713 13512
rect 34664 13472 34670 13484
rect 34701 13481 34713 13484
rect 34747 13481 34759 13515
rect 34701 13475 34759 13481
rect 37277 13447 37335 13453
rect 37277 13444 37289 13447
rect 22066 13416 37289 13444
rect 3973 13379 4031 13385
rect 3973 13345 3985 13379
rect 4019 13376 4031 13379
rect 4706 13376 4712 13388
rect 4019 13348 4712 13376
rect 4019 13345 4031 13348
rect 3973 13339 4031 13345
rect 4706 13336 4712 13348
rect 4764 13336 4770 13388
rect 7466 13336 7472 13388
rect 7524 13376 7530 13388
rect 22066 13376 22094 13416
rect 37277 13413 37289 13416
rect 37323 13413 37335 13447
rect 37277 13407 37335 13413
rect 7524 13348 22094 13376
rect 7524 13336 7530 13348
rect 34422 13336 34428 13388
rect 34480 13376 34486 13388
rect 35253 13379 35311 13385
rect 35253 13376 35265 13379
rect 34480 13348 35265 13376
rect 34480 13336 34486 13348
rect 35253 13345 35265 13348
rect 35299 13345 35311 13379
rect 35253 13339 35311 13345
rect 1394 13308 1400 13320
rect 1355 13280 1400 13308
rect 1394 13268 1400 13280
rect 1452 13308 1458 13320
rect 2593 13311 2651 13317
rect 2593 13308 2605 13311
rect 1452 13280 2605 13308
rect 1452 13268 1458 13280
rect 2593 13277 2605 13280
rect 2639 13277 2651 13311
rect 2593 13271 2651 13277
rect 4157 13311 4215 13317
rect 4157 13277 4169 13311
rect 4203 13308 4215 13311
rect 5074 13308 5080 13320
rect 4203 13280 5080 13308
rect 4203 13277 4215 13280
rect 4157 13271 4215 13277
rect 5074 13268 5080 13280
rect 5132 13268 5138 13320
rect 26878 13308 26884 13320
rect 26839 13280 26884 13308
rect 26878 13268 26884 13280
rect 26936 13268 26942 13320
rect 33962 13308 33968 13320
rect 33923 13280 33968 13308
rect 33962 13268 33968 13280
rect 34020 13268 34026 13320
rect 35066 13308 35072 13320
rect 34072 13280 35072 13308
rect 4065 13243 4123 13249
rect 4065 13240 4077 13243
rect 1596 13212 4077 13240
rect 1596 13181 1624 13212
rect 4065 13209 4077 13212
rect 4111 13209 4123 13243
rect 4065 13203 4123 13209
rect 1581 13175 1639 13181
rect 1581 13141 1593 13175
rect 1627 13141 1639 13175
rect 1581 13135 1639 13141
rect 4706 13132 4712 13184
rect 4764 13172 4770 13184
rect 4985 13175 5043 13181
rect 4985 13172 4997 13175
rect 4764 13144 4997 13172
rect 4764 13132 4770 13144
rect 4985 13141 4997 13144
rect 5031 13141 5043 13175
rect 4985 13135 5043 13141
rect 27065 13175 27123 13181
rect 27065 13141 27077 13175
rect 27111 13172 27123 13175
rect 34072 13172 34100 13280
rect 35066 13268 35072 13280
rect 35124 13268 35130 13320
rect 35161 13311 35219 13317
rect 35161 13277 35173 13311
rect 35207 13277 35219 13311
rect 35161 13271 35219 13277
rect 34974 13240 34980 13252
rect 34164 13212 34980 13240
rect 34164 13181 34192 13212
rect 34974 13200 34980 13212
rect 35032 13200 35038 13252
rect 35176 13240 35204 13271
rect 35342 13268 35348 13320
rect 35400 13308 35406 13320
rect 36814 13308 36820 13320
rect 35400 13280 36820 13308
rect 35400 13268 35406 13280
rect 36814 13268 36820 13280
rect 36872 13268 36878 13320
rect 37292 13308 37320 13407
rect 37829 13311 37887 13317
rect 37829 13308 37841 13311
rect 37292 13280 37841 13308
rect 37829 13277 37841 13280
rect 37875 13277 37887 13311
rect 37829 13271 37887 13277
rect 37918 13240 37924 13252
rect 35176 13212 37924 13240
rect 37918 13200 37924 13212
rect 37976 13200 37982 13252
rect 27111 13144 34100 13172
rect 34149 13175 34207 13181
rect 27111 13141 27123 13144
rect 27065 13135 27123 13141
rect 34149 13141 34161 13175
rect 34195 13141 34207 13175
rect 34149 13135 34207 13141
rect 34606 13132 34612 13184
rect 34664 13172 34670 13184
rect 35069 13175 35127 13181
rect 35069 13172 35081 13175
rect 34664 13144 35081 13172
rect 34664 13132 34670 13144
rect 35069 13141 35081 13144
rect 35115 13141 35127 13175
rect 35069 13135 35127 13141
rect 35342 13132 35348 13184
rect 35400 13172 35406 13184
rect 37826 13172 37832 13184
rect 35400 13144 37832 13172
rect 35400 13132 35406 13144
rect 37826 13132 37832 13144
rect 37884 13132 37890 13184
rect 38010 13172 38016 13184
rect 37971 13144 38016 13172
rect 38010 13132 38016 13144
rect 38068 13132 38074 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 12986 12900 12992 12912
rect 12947 12872 12992 12900
rect 12986 12860 12992 12872
rect 13044 12860 13050 12912
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12832 1731 12835
rect 10594 12832 10600 12844
rect 1719 12804 10600 12832
rect 1719 12801 1731 12804
rect 1673 12795 1731 12801
rect 10594 12792 10600 12804
rect 10652 12792 10658 12844
rect 37642 12792 37648 12844
rect 37700 12832 37706 12844
rect 37829 12835 37887 12841
rect 37829 12832 37841 12835
rect 37700 12804 37841 12832
rect 37700 12792 37706 12804
rect 37829 12801 37841 12804
rect 37875 12801 37887 12835
rect 37829 12795 37887 12801
rect 38102 12764 38108 12776
rect 38063 12736 38108 12764
rect 38102 12724 38108 12736
rect 38160 12724 38166 12776
rect 1486 12628 1492 12640
rect 1447 12600 1492 12628
rect 1486 12588 1492 12600
rect 1544 12588 1550 12640
rect 13906 12588 13912 12640
rect 13964 12628 13970 12640
rect 14277 12631 14335 12637
rect 14277 12628 14289 12631
rect 13964 12600 14289 12628
rect 13964 12588 13970 12600
rect 14277 12597 14289 12600
rect 14323 12597 14335 12631
rect 14277 12591 14335 12597
rect 34422 12588 34428 12640
rect 34480 12628 34486 12640
rect 34517 12631 34575 12637
rect 34517 12628 34529 12631
rect 34480 12600 34529 12628
rect 34480 12588 34486 12600
rect 34517 12597 34529 12600
rect 34563 12597 34575 12631
rect 34517 12591 34575 12597
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 10594 12424 10600 12436
rect 10555 12396 10600 12424
rect 10594 12384 10600 12396
rect 10652 12384 10658 12436
rect 14642 12384 14648 12436
rect 14700 12424 14706 12436
rect 20162 12424 20168 12436
rect 14700 12396 20168 12424
rect 14700 12384 14706 12396
rect 20162 12384 20168 12396
rect 20220 12424 20226 12436
rect 34422 12424 34428 12436
rect 20220 12396 34428 12424
rect 20220 12384 20226 12396
rect 34422 12384 34428 12396
rect 34480 12384 34486 12436
rect 38102 12356 38108 12368
rect 38063 12328 38108 12356
rect 38102 12316 38108 12328
rect 38160 12316 38166 12368
rect 11790 12288 11796 12300
rect 11751 12260 11796 12288
rect 11790 12248 11796 12260
rect 11848 12248 11854 12300
rect 10781 12223 10839 12229
rect 10781 12189 10793 12223
rect 10827 12220 10839 12223
rect 10827 12192 11284 12220
rect 10827 12189 10839 12192
rect 10781 12183 10839 12189
rect 1486 12084 1492 12096
rect 1447 12056 1492 12084
rect 1486 12044 1492 12056
rect 1544 12044 1550 12096
rect 11256 12093 11284 12192
rect 11241 12087 11299 12093
rect 11241 12053 11253 12087
rect 11287 12053 11299 12087
rect 11606 12084 11612 12096
rect 11567 12056 11612 12084
rect 11241 12047 11299 12053
rect 11606 12044 11612 12056
rect 11664 12044 11670 12096
rect 11701 12087 11759 12093
rect 11701 12053 11713 12087
rect 11747 12084 11759 12087
rect 17770 12084 17776 12096
rect 11747 12056 17776 12084
rect 11747 12053 11759 12056
rect 11701 12047 11759 12053
rect 17770 12044 17776 12056
rect 17828 12044 17834 12096
rect 37274 12044 37280 12096
rect 37332 12084 37338 12096
rect 37461 12087 37519 12093
rect 37461 12084 37473 12087
rect 37332 12056 37473 12084
rect 37332 12044 37338 12056
rect 37461 12053 37473 12056
rect 37507 12053 37519 12087
rect 37461 12047 37519 12053
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 3970 11840 3976 11892
rect 4028 11880 4034 11892
rect 4065 11883 4123 11889
rect 4065 11880 4077 11883
rect 4028 11852 4077 11880
rect 4028 11840 4034 11852
rect 4065 11849 4077 11852
rect 4111 11849 4123 11883
rect 4065 11843 4123 11849
rect 4525 11883 4583 11889
rect 4525 11849 4537 11883
rect 4571 11880 4583 11883
rect 4798 11880 4804 11892
rect 4571 11852 4804 11880
rect 4571 11849 4583 11852
rect 4525 11843 4583 11849
rect 4798 11840 4804 11852
rect 4856 11840 4862 11892
rect 22094 11840 22100 11892
rect 22152 11880 22158 11892
rect 29730 11880 29736 11892
rect 22152 11852 29736 11880
rect 22152 11840 22158 11852
rect 29730 11840 29736 11852
rect 29788 11840 29794 11892
rect 2041 11815 2099 11821
rect 2041 11781 2053 11815
rect 2087 11812 2099 11815
rect 8294 11812 8300 11824
rect 2087 11784 8300 11812
rect 2087 11781 2099 11784
rect 2041 11775 2099 11781
rect 8294 11772 8300 11784
rect 8352 11812 8358 11824
rect 11517 11815 11575 11821
rect 11517 11812 11529 11815
rect 8352 11784 11529 11812
rect 8352 11772 8358 11784
rect 11517 11781 11529 11784
rect 11563 11812 11575 11815
rect 11790 11812 11796 11824
rect 11563 11784 11796 11812
rect 11563 11781 11575 11784
rect 11517 11775 11575 11781
rect 11790 11772 11796 11784
rect 11848 11812 11854 11824
rect 14642 11812 14648 11824
rect 11848 11784 14648 11812
rect 11848 11772 11854 11784
rect 14642 11772 14648 11784
rect 14700 11772 14706 11824
rect 26786 11772 26792 11824
rect 26844 11812 26850 11824
rect 37090 11812 37096 11824
rect 26844 11784 37096 11812
rect 26844 11772 26850 11784
rect 37090 11772 37096 11784
rect 37148 11772 37154 11824
rect 1486 11744 1492 11756
rect 1447 11716 1492 11744
rect 1486 11704 1492 11716
rect 1544 11704 1550 11756
rect 1854 11704 1860 11756
rect 1912 11744 1918 11756
rect 4157 11747 4215 11753
rect 1912 11716 4108 11744
rect 1912 11704 1918 11716
rect 3881 11679 3939 11685
rect 3881 11645 3893 11679
rect 3927 11645 3939 11679
rect 4080 11676 4108 11716
rect 4157 11713 4169 11747
rect 4203 11744 4215 11747
rect 4614 11744 4620 11756
rect 4203 11716 4620 11744
rect 4203 11713 4215 11716
rect 4157 11707 4215 11713
rect 4614 11704 4620 11716
rect 4672 11704 4678 11756
rect 14826 11744 14832 11756
rect 14787 11716 14832 11744
rect 14826 11704 14832 11716
rect 14884 11704 14890 11756
rect 23474 11704 23480 11756
rect 23532 11744 23538 11756
rect 37642 11744 37648 11756
rect 23532 11716 37648 11744
rect 23532 11704 23538 11716
rect 37642 11704 37648 11716
rect 37700 11704 37706 11756
rect 10873 11679 10931 11685
rect 10873 11676 10885 11679
rect 4080 11648 10885 11676
rect 3881 11639 3939 11645
rect 10873 11645 10885 11648
rect 10919 11676 10931 11679
rect 11606 11676 11612 11688
rect 10919 11648 11612 11676
rect 10919 11645 10931 11648
rect 10873 11639 10931 11645
rect 3896 11608 3924 11639
rect 11606 11636 11612 11648
rect 11664 11636 11670 11688
rect 14553 11679 14611 11685
rect 14553 11645 14565 11679
rect 14599 11676 14611 11679
rect 15010 11676 15016 11688
rect 14599 11648 15016 11676
rect 14599 11645 14611 11648
rect 14553 11639 14611 11645
rect 15010 11636 15016 11648
rect 15068 11636 15074 11688
rect 37274 11676 37280 11688
rect 37235 11648 37280 11676
rect 37274 11636 37280 11648
rect 37332 11636 37338 11688
rect 37553 11679 37611 11685
rect 37553 11645 37565 11679
rect 37599 11645 37611 11679
rect 37553 11639 37611 11645
rect 3896 11580 4752 11608
rect 4724 11552 4752 11580
rect 9766 11568 9772 11620
rect 9824 11608 9830 11620
rect 20990 11608 20996 11620
rect 9824 11580 20996 11608
rect 9824 11568 9830 11580
rect 20990 11568 20996 11580
rect 21048 11568 21054 11620
rect 29822 11568 29828 11620
rect 29880 11608 29886 11620
rect 37568 11608 37596 11639
rect 29880 11580 37596 11608
rect 29880 11568 29886 11580
rect 4706 11500 4712 11552
rect 4764 11540 4770 11552
rect 4985 11543 5043 11549
rect 4985 11540 4997 11543
rect 4764 11512 4997 11540
rect 4764 11500 4770 11512
rect 4985 11509 4997 11512
rect 5031 11509 5043 11543
rect 4985 11503 5043 11509
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 1581 11339 1639 11345
rect 1581 11305 1593 11339
rect 1627 11336 1639 11339
rect 1670 11336 1676 11348
rect 1627 11308 1676 11336
rect 1627 11305 1639 11308
rect 1581 11299 1639 11305
rect 1670 11296 1676 11308
rect 1728 11296 1734 11348
rect 37918 11336 37924 11348
rect 37879 11308 37924 11336
rect 37918 11296 37924 11308
rect 37976 11296 37982 11348
rect 1394 11132 1400 11144
rect 1355 11104 1400 11132
rect 1394 11092 1400 11104
rect 1452 11132 1458 11144
rect 2041 11135 2099 11141
rect 2041 11132 2053 11135
rect 1452 11104 2053 11132
rect 1452 11092 1458 11104
rect 2041 11101 2053 11104
rect 2087 11101 2099 11135
rect 2041 11095 2099 11101
rect 37461 11135 37519 11141
rect 37461 11101 37473 11135
rect 37507 11132 37519 11135
rect 38102 11132 38108 11144
rect 37507 11104 38108 11132
rect 37507 11101 37519 11104
rect 37461 11095 37519 11101
rect 38102 11092 38108 11104
rect 38160 11092 38166 11144
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 2406 10752 2412 10804
rect 2464 10792 2470 10804
rect 8294 10792 8300 10804
rect 2464 10764 6914 10792
rect 8255 10764 8300 10792
rect 2464 10752 2470 10764
rect 6886 10724 6914 10764
rect 8294 10752 8300 10764
rect 8352 10752 8358 10804
rect 7745 10727 7803 10733
rect 7745 10724 7757 10727
rect 6886 10696 7757 10724
rect 7745 10693 7757 10696
rect 7791 10724 7803 10727
rect 9033 10727 9091 10733
rect 9033 10724 9045 10727
rect 7791 10696 9045 10724
rect 7791 10693 7803 10696
rect 7745 10687 7803 10693
rect 9033 10693 9045 10696
rect 9079 10693 9091 10727
rect 15565 10727 15623 10733
rect 15565 10724 15577 10727
rect 9033 10687 9091 10693
rect 14568 10696 15577 10724
rect 1394 10656 1400 10668
rect 1355 10628 1400 10656
rect 1394 10616 1400 10628
rect 1452 10656 1458 10668
rect 2041 10659 2099 10665
rect 2041 10656 2053 10659
rect 1452 10628 2053 10656
rect 1452 10616 1458 10628
rect 2041 10625 2053 10628
rect 2087 10625 2099 10659
rect 2041 10619 2099 10625
rect 6178 10616 6184 10668
rect 6236 10656 6242 10668
rect 9125 10659 9183 10665
rect 9125 10656 9137 10659
rect 6236 10628 9137 10656
rect 6236 10616 6242 10628
rect 9125 10625 9137 10628
rect 9171 10625 9183 10659
rect 9125 10619 9183 10625
rect 14568 10600 14596 10696
rect 15565 10693 15577 10696
rect 15611 10693 15623 10727
rect 15565 10687 15623 10693
rect 14734 10656 14740 10668
rect 14695 10628 14740 10656
rect 14734 10616 14740 10628
rect 14792 10616 14798 10668
rect 37461 10659 37519 10665
rect 37461 10625 37473 10659
rect 37507 10656 37519 10659
rect 38102 10656 38108 10668
rect 37507 10628 38108 10656
rect 37507 10625 37519 10628
rect 37461 10619 37519 10625
rect 38102 10616 38108 10628
rect 38160 10616 38166 10668
rect 8294 10548 8300 10600
rect 8352 10588 8358 10600
rect 8849 10591 8907 10597
rect 8849 10588 8861 10591
rect 8352 10560 8861 10588
rect 8352 10548 8358 10560
rect 8849 10557 8861 10560
rect 8895 10557 8907 10591
rect 14550 10588 14556 10600
rect 14511 10560 14556 10588
rect 8849 10551 8907 10557
rect 14550 10548 14556 10560
rect 14608 10548 14614 10600
rect 14645 10591 14703 10597
rect 14645 10557 14657 10591
rect 14691 10557 14703 10591
rect 37274 10588 37280 10600
rect 14645 10551 14703 10557
rect 26206 10560 37280 10588
rect 2498 10480 2504 10532
rect 2556 10520 2562 10532
rect 13817 10523 13875 10529
rect 13817 10520 13829 10523
rect 2556 10492 13829 10520
rect 2556 10480 2562 10492
rect 13817 10489 13829 10492
rect 13863 10520 13875 10523
rect 14660 10520 14688 10551
rect 13863 10492 14688 10520
rect 13863 10489 13875 10492
rect 13817 10483 13875 10489
rect 23382 10480 23388 10532
rect 23440 10520 23446 10532
rect 26206 10520 26234 10560
rect 37274 10548 37280 10560
rect 37332 10548 37338 10600
rect 37921 10523 37979 10529
rect 37921 10520 37933 10523
rect 23440 10492 26234 10520
rect 35866 10492 37933 10520
rect 23440 10480 23446 10492
rect 1578 10452 1584 10464
rect 1539 10424 1584 10452
rect 1578 10412 1584 10424
rect 1636 10412 1642 10464
rect 9493 10455 9551 10461
rect 9493 10421 9505 10455
rect 9539 10452 9551 10455
rect 12158 10452 12164 10464
rect 9539 10424 12164 10452
rect 9539 10421 9551 10424
rect 9493 10415 9551 10421
rect 12158 10412 12164 10424
rect 12216 10412 12222 10464
rect 15102 10452 15108 10464
rect 15063 10424 15108 10452
rect 15102 10412 15108 10424
rect 15160 10412 15166 10464
rect 23750 10412 23756 10464
rect 23808 10452 23814 10464
rect 35866 10452 35894 10492
rect 37921 10489 37933 10492
rect 37967 10489 37979 10523
rect 37921 10483 37979 10489
rect 23808 10424 35894 10452
rect 23808 10412 23814 10424
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 1578 10208 1584 10260
rect 1636 10248 1642 10260
rect 14734 10248 14740 10260
rect 1636 10220 14740 10248
rect 1636 10208 1642 10220
rect 14734 10208 14740 10220
rect 14792 10208 14798 10260
rect 37550 10208 37556 10260
rect 37608 10248 37614 10260
rect 37921 10251 37979 10257
rect 37921 10248 37933 10251
rect 37608 10220 37933 10248
rect 37608 10208 37614 10220
rect 37921 10217 37933 10220
rect 37967 10217 37979 10251
rect 37921 10211 37979 10217
rect 12345 10183 12403 10189
rect 12345 10149 12357 10183
rect 12391 10180 12403 10183
rect 17218 10180 17224 10192
rect 12391 10152 17224 10180
rect 12391 10149 12403 10152
rect 12345 10143 12403 10149
rect 17218 10140 17224 10152
rect 17276 10140 17282 10192
rect 1394 10044 1400 10056
rect 1355 10016 1400 10044
rect 1394 10004 1400 10016
rect 1452 10044 1458 10056
rect 2041 10047 2099 10053
rect 2041 10044 2053 10047
rect 1452 10016 2053 10044
rect 1452 10004 1458 10016
rect 2041 10013 2053 10016
rect 2087 10013 2099 10047
rect 12158 10044 12164 10056
rect 12119 10016 12164 10044
rect 2041 10007 2099 10013
rect 12158 10004 12164 10016
rect 12216 10004 12222 10056
rect 15102 10004 15108 10056
rect 15160 10044 15166 10056
rect 15841 10047 15899 10053
rect 15841 10044 15853 10047
rect 15160 10016 15853 10044
rect 15160 10004 15166 10016
rect 15841 10013 15853 10016
rect 15887 10013 15899 10047
rect 15841 10007 15899 10013
rect 37369 10047 37427 10053
rect 37369 10013 37381 10047
rect 37415 10044 37427 10047
rect 38102 10044 38108 10056
rect 37415 10016 38108 10044
rect 37415 10013 37427 10016
rect 37369 10007 37427 10013
rect 38102 10004 38108 10016
rect 38160 10004 38166 10056
rect 14918 9976 14924 9988
rect 1596 9948 14924 9976
rect 1596 9917 1624 9948
rect 14918 9936 14924 9948
rect 14976 9936 14982 9988
rect 1581 9911 1639 9917
rect 1581 9877 1593 9911
rect 1627 9877 1639 9911
rect 1581 9871 1639 9877
rect 16025 9911 16083 9917
rect 16025 9877 16037 9911
rect 16071 9908 16083 9911
rect 18138 9908 18144 9920
rect 16071 9880 18144 9908
rect 16071 9877 16083 9880
rect 16025 9871 16083 9877
rect 18138 9868 18144 9880
rect 18196 9868 18202 9920
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 14642 9596 14648 9648
rect 14700 9636 14706 9648
rect 14700 9608 15608 9636
rect 14700 9596 14706 9608
rect 15470 9568 15476 9580
rect 15431 9540 15476 9568
rect 15470 9528 15476 9540
rect 15528 9528 15534 9580
rect 15580 9568 15608 9608
rect 15580 9540 15700 9568
rect 14642 9500 14648 9512
rect 14603 9472 14648 9500
rect 14642 9460 14648 9472
rect 14700 9460 14706 9512
rect 15672 9509 15700 9540
rect 15565 9503 15623 9509
rect 15565 9469 15577 9503
rect 15611 9469 15623 9503
rect 15565 9463 15623 9469
rect 15657 9503 15715 9509
rect 15657 9469 15669 9503
rect 15703 9469 15715 9503
rect 15657 9463 15715 9469
rect 15010 9392 15016 9444
rect 15068 9432 15074 9444
rect 15105 9435 15163 9441
rect 15105 9432 15117 9435
rect 15068 9404 15117 9432
rect 15068 9392 15074 9404
rect 15105 9401 15117 9404
rect 15151 9401 15163 9435
rect 15105 9395 15163 9401
rect 15580 9364 15608 9463
rect 16761 9367 16819 9373
rect 16761 9364 16773 9367
rect 15580 9336 16773 9364
rect 16761 9333 16773 9336
rect 16807 9364 16819 9367
rect 30926 9364 30932 9376
rect 16807 9336 30932 9364
rect 16807 9333 16819 9336
rect 16761 9327 16819 9333
rect 30926 9324 30932 9336
rect 30984 9324 30990 9376
rect 38102 9364 38108 9376
rect 38063 9336 38108 9364
rect 38102 9324 38108 9336
rect 38160 9324 38166 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 33778 8984 33784 9036
rect 33836 9024 33842 9036
rect 37829 9027 37887 9033
rect 37829 9024 37841 9027
rect 33836 8996 37841 9024
rect 33836 8984 33842 8996
rect 37829 8993 37841 8996
rect 37875 8993 37887 9027
rect 37829 8987 37887 8993
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8925 1731 8959
rect 38102 8956 38108 8968
rect 38063 8928 38108 8956
rect 1673 8919 1731 8925
rect 1688 8888 1716 8919
rect 38102 8916 38108 8928
rect 38160 8916 38166 8968
rect 2225 8891 2283 8897
rect 2225 8888 2237 8891
rect 1688 8860 2237 8888
rect 2225 8857 2237 8860
rect 2271 8888 2283 8891
rect 19334 8888 19340 8900
rect 2271 8860 19340 8888
rect 2271 8857 2283 8860
rect 2225 8851 2283 8857
rect 19334 8848 19340 8860
rect 19392 8848 19398 8900
rect 1486 8820 1492 8832
rect 1447 8792 1492 8820
rect 1486 8780 1492 8792
rect 1544 8780 1550 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 14918 8576 14924 8628
rect 14976 8616 14982 8628
rect 15657 8619 15715 8625
rect 15657 8616 15669 8619
rect 14976 8588 15669 8616
rect 14976 8576 14982 8588
rect 15657 8585 15669 8588
rect 15703 8585 15715 8619
rect 15657 8579 15715 8585
rect 1949 8483 2007 8489
rect 1949 8449 1961 8483
rect 1995 8480 2007 8483
rect 3694 8480 3700 8492
rect 1995 8452 3700 8480
rect 1995 8449 2007 8452
rect 1949 8443 2007 8449
rect 3694 8440 3700 8452
rect 3752 8440 3758 8492
rect 15749 8483 15807 8489
rect 15749 8449 15761 8483
rect 15795 8480 15807 8483
rect 15930 8480 15936 8492
rect 15795 8452 15936 8480
rect 15795 8449 15807 8452
rect 15749 8443 15807 8449
rect 15930 8440 15936 8452
rect 15988 8440 15994 8492
rect 16298 8440 16304 8492
rect 16356 8480 16362 8492
rect 37277 8483 37335 8489
rect 37277 8480 37289 8483
rect 16356 8452 37289 8480
rect 16356 8440 16362 8452
rect 37277 8449 37289 8452
rect 37323 8480 37335 8483
rect 37829 8483 37887 8489
rect 37829 8480 37841 8483
rect 37323 8452 37841 8480
rect 37323 8449 37335 8452
rect 37277 8443 37335 8449
rect 37829 8449 37841 8452
rect 37875 8449 37887 8483
rect 37829 8443 37887 8449
rect 2222 8412 2228 8424
rect 2183 8384 2228 8412
rect 2222 8372 2228 8384
rect 2280 8412 2286 8424
rect 2685 8415 2743 8421
rect 2685 8412 2697 8415
rect 2280 8384 2697 8412
rect 2280 8372 2286 8384
rect 2685 8381 2697 8384
rect 2731 8381 2743 8415
rect 2685 8375 2743 8381
rect 15565 8415 15623 8421
rect 15565 8381 15577 8415
rect 15611 8381 15623 8415
rect 15565 8375 15623 8381
rect 15580 8344 15608 8375
rect 16761 8347 16819 8353
rect 16761 8344 16773 8347
rect 15580 8316 16773 8344
rect 16761 8313 16773 8316
rect 16807 8344 16819 8347
rect 17954 8344 17960 8356
rect 16807 8316 17960 8344
rect 16807 8313 16819 8316
rect 16761 8307 16819 8313
rect 17954 8304 17960 8316
rect 18012 8304 18018 8356
rect 38010 8344 38016 8356
rect 37971 8316 38016 8344
rect 38010 8304 38016 8316
rect 38068 8304 38074 8356
rect 16114 8276 16120 8288
rect 16075 8248 16120 8276
rect 16114 8236 16120 8248
rect 16172 8236 16178 8288
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 1949 7939 2007 7945
rect 1949 7905 1961 7939
rect 1995 7936 2007 7939
rect 13814 7936 13820 7948
rect 1995 7908 13820 7936
rect 1995 7905 2007 7908
rect 1949 7899 2007 7905
rect 13814 7896 13820 7908
rect 13872 7896 13878 7948
rect 16114 7896 16120 7948
rect 16172 7936 16178 7948
rect 16301 7939 16359 7945
rect 16301 7936 16313 7939
rect 16172 7908 16313 7936
rect 16172 7896 16178 7908
rect 16301 7905 16313 7908
rect 16347 7905 16359 7939
rect 16301 7899 16359 7905
rect 2038 7828 2044 7880
rect 2096 7868 2102 7880
rect 2225 7871 2283 7877
rect 2225 7868 2237 7871
rect 2096 7840 2237 7868
rect 2096 7828 2102 7840
rect 2225 7837 2237 7840
rect 2271 7837 2283 7871
rect 2225 7831 2283 7837
rect 16577 7871 16635 7877
rect 16577 7837 16589 7871
rect 16623 7868 16635 7871
rect 16623 7840 26234 7868
rect 16623 7837 16635 7840
rect 16577 7831 16635 7837
rect 26206 7800 26234 7840
rect 31018 7828 31024 7880
rect 31076 7868 31082 7880
rect 37829 7871 37887 7877
rect 37829 7868 37841 7871
rect 31076 7840 37841 7868
rect 31076 7828 31082 7840
rect 37829 7837 37841 7840
rect 37875 7837 37887 7871
rect 37829 7831 37887 7837
rect 36170 7800 36176 7812
rect 26206 7772 36176 7800
rect 36170 7760 36176 7772
rect 36228 7760 36234 7812
rect 38010 7732 38016 7744
rect 37971 7704 38016 7732
rect 38010 7692 38016 7704
rect 38068 7692 38074 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 2038 7528 2044 7540
rect 1999 7500 2044 7528
rect 2038 7488 2044 7500
rect 2096 7488 2102 7540
rect 1394 7392 1400 7404
rect 1355 7364 1400 7392
rect 1394 7352 1400 7364
rect 1452 7352 1458 7404
rect 22554 7392 22560 7404
rect 22515 7364 22560 7392
rect 22554 7352 22560 7364
rect 22612 7352 22618 7404
rect 37369 7395 37427 7401
rect 37369 7361 37381 7395
rect 37415 7392 37427 7395
rect 38010 7392 38016 7404
rect 37415 7364 38016 7392
rect 37415 7361 37427 7364
rect 37369 7355 37427 7361
rect 38010 7352 38016 7364
rect 38068 7352 38074 7404
rect 4890 7284 4896 7336
rect 4948 7324 4954 7336
rect 37829 7327 37887 7333
rect 37829 7324 37841 7327
rect 4948 7296 37841 7324
rect 4948 7284 4954 7296
rect 37829 7293 37841 7296
rect 37875 7293 37887 7327
rect 37829 7287 37887 7293
rect 1581 7259 1639 7265
rect 1581 7225 1593 7259
rect 1627 7256 1639 7259
rect 4614 7256 4620 7268
rect 1627 7228 4620 7256
rect 1627 7225 1639 7228
rect 1581 7219 1639 7225
rect 4614 7216 4620 7228
rect 4672 7216 4678 7268
rect 22741 7259 22799 7265
rect 22741 7225 22753 7259
rect 22787 7256 22799 7259
rect 31018 7256 31024 7268
rect 22787 7228 31024 7256
rect 22787 7225 22799 7228
rect 22741 7219 22799 7225
rect 31018 7216 31024 7228
rect 31076 7216 31082 7268
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1394 6916 1400 6928
rect 1355 6888 1400 6916
rect 1394 6876 1400 6888
rect 1452 6876 1458 6928
rect 10597 6851 10655 6857
rect 10597 6817 10609 6851
rect 10643 6848 10655 6851
rect 10686 6848 10692 6860
rect 10643 6820 10692 6848
rect 10643 6817 10655 6820
rect 10597 6811 10655 6817
rect 10686 6808 10692 6820
rect 10744 6808 10750 6860
rect 12158 6808 12164 6860
rect 12216 6848 12222 6860
rect 12437 6851 12495 6857
rect 12437 6848 12449 6851
rect 12216 6820 12449 6848
rect 12216 6808 12222 6820
rect 12437 6817 12449 6820
rect 12483 6848 12495 6851
rect 17954 6848 17960 6860
rect 12483 6820 17960 6848
rect 12483 6817 12495 6820
rect 12437 6811 12495 6817
rect 17954 6808 17960 6820
rect 18012 6808 18018 6860
rect 21913 6851 21971 6857
rect 21913 6817 21925 6851
rect 21959 6848 21971 6851
rect 22554 6848 22560 6860
rect 21959 6820 22560 6848
rect 21959 6817 21971 6820
rect 21913 6811 21971 6817
rect 22554 6808 22560 6820
rect 22612 6808 22618 6860
rect 21726 6780 21732 6792
rect 21687 6752 21732 6780
rect 21726 6740 21732 6752
rect 21784 6780 21790 6792
rect 21784 6752 22094 6780
rect 21784 6740 21790 6752
rect 10781 6715 10839 6721
rect 10781 6681 10793 6715
rect 10827 6712 10839 6715
rect 11514 6712 11520 6724
rect 10827 6684 11520 6712
rect 10827 6681 10839 6684
rect 10781 6675 10839 6681
rect 11514 6672 11520 6684
rect 11572 6672 11578 6724
rect 21542 6712 21548 6724
rect 21503 6684 21548 6712
rect 21542 6672 21548 6684
rect 21600 6672 21606 6724
rect 22066 6644 22094 6752
rect 22465 6647 22523 6653
rect 22465 6644 22477 6647
rect 22066 6616 22477 6644
rect 22465 6613 22477 6616
rect 22511 6644 22523 6647
rect 30466 6644 30472 6656
rect 22511 6616 30472 6644
rect 22511 6613 22523 6616
rect 22465 6607 22523 6613
rect 30466 6604 30472 6616
rect 30524 6604 30530 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 11514 6440 11520 6452
rect 11475 6412 11520 6440
rect 11514 6400 11520 6412
rect 11572 6400 11578 6452
rect 17954 6400 17960 6452
rect 18012 6440 18018 6452
rect 24213 6443 24271 6449
rect 24213 6440 24225 6443
rect 18012 6412 24225 6440
rect 18012 6400 18018 6412
rect 24213 6409 24225 6412
rect 24259 6440 24271 6443
rect 24946 6440 24952 6452
rect 24259 6412 24952 6440
rect 24259 6409 24271 6412
rect 24213 6403 24271 6409
rect 24946 6400 24952 6412
rect 25004 6400 25010 6452
rect 37274 6440 37280 6452
rect 37235 6412 37280 6440
rect 37274 6400 37280 6412
rect 37332 6400 37338 6452
rect 2314 6332 2320 6384
rect 2372 6372 2378 6384
rect 20714 6372 20720 6384
rect 2372 6344 20720 6372
rect 2372 6332 2378 6344
rect 20714 6332 20720 6344
rect 20772 6332 20778 6384
rect 1673 6307 1731 6313
rect 1673 6273 1685 6307
rect 1719 6304 1731 6307
rect 1762 6304 1768 6316
rect 1719 6276 1768 6304
rect 1719 6273 1731 6276
rect 1673 6267 1731 6273
rect 1762 6264 1768 6276
rect 1820 6304 1826 6316
rect 2133 6307 2191 6313
rect 2133 6304 2145 6307
rect 1820 6276 2145 6304
rect 1820 6264 1826 6276
rect 2133 6273 2145 6276
rect 2179 6273 2191 6307
rect 2133 6267 2191 6273
rect 11885 6307 11943 6313
rect 11885 6273 11897 6307
rect 11931 6273 11943 6307
rect 11885 6267 11943 6273
rect 13817 6307 13875 6313
rect 13817 6273 13829 6307
rect 13863 6304 13875 6307
rect 14737 6307 14795 6313
rect 14737 6304 14749 6307
rect 13863 6276 14749 6304
rect 13863 6273 13875 6276
rect 13817 6267 13875 6273
rect 14737 6273 14749 6276
rect 14783 6304 14795 6307
rect 37292 6304 37320 6400
rect 37829 6307 37887 6313
rect 37829 6304 37841 6307
rect 14783 6276 26234 6304
rect 37292 6276 37841 6304
rect 14783 6273 14795 6276
rect 14737 6267 14795 6273
rect 1486 6168 1492 6180
rect 1447 6140 1492 6168
rect 1486 6128 1492 6140
rect 1544 6128 1550 6180
rect 11900 6100 11928 6267
rect 11974 6196 11980 6248
rect 12032 6236 12038 6248
rect 12158 6236 12164 6248
rect 12032 6208 12077 6236
rect 12119 6208 12164 6236
rect 12032 6196 12038 6208
rect 12158 6196 12164 6208
rect 12216 6196 12222 6248
rect 12250 6196 12256 6248
rect 12308 6236 12314 6248
rect 13909 6239 13967 6245
rect 13909 6236 13921 6239
rect 12308 6208 13921 6236
rect 12308 6196 12314 6208
rect 13909 6205 13921 6208
rect 13955 6205 13967 6239
rect 13909 6199 13967 6205
rect 14093 6239 14151 6245
rect 14093 6205 14105 6239
rect 14139 6236 14151 6239
rect 14550 6236 14556 6248
rect 14139 6208 14556 6236
rect 14139 6205 14151 6208
rect 14093 6199 14151 6205
rect 14550 6196 14556 6208
rect 14608 6196 14614 6248
rect 26206 6236 26234 6276
rect 37829 6273 37841 6276
rect 37875 6273 37887 6307
rect 37829 6267 37887 6273
rect 38378 6236 38384 6248
rect 26206 6208 38384 6236
rect 38378 6196 38384 6208
rect 38436 6196 38442 6248
rect 38010 6168 38016 6180
rect 37971 6140 38016 6168
rect 38010 6128 38016 6140
rect 38068 6128 38074 6180
rect 12802 6100 12808 6112
rect 11900 6072 12808 6100
rect 12802 6060 12808 6072
rect 12860 6060 12866 6112
rect 12986 6060 12992 6112
rect 13044 6100 13050 6112
rect 13449 6103 13507 6109
rect 13449 6100 13461 6103
rect 13044 6072 13461 6100
rect 13044 6060 13050 6072
rect 13449 6069 13461 6072
rect 13495 6069 13507 6103
rect 13449 6063 13507 6069
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 14369 5899 14427 5905
rect 14369 5865 14381 5899
rect 14415 5896 14427 5899
rect 14550 5896 14556 5908
rect 14415 5868 14556 5896
rect 14415 5865 14427 5868
rect 14369 5859 14427 5865
rect 14550 5856 14556 5868
rect 14608 5896 14614 5908
rect 17310 5896 17316 5908
rect 14608 5868 17316 5896
rect 14608 5856 14614 5868
rect 17310 5856 17316 5868
rect 17368 5856 17374 5908
rect 25406 5856 25412 5908
rect 25464 5896 25470 5908
rect 25593 5899 25651 5905
rect 25593 5896 25605 5899
rect 25464 5868 25605 5896
rect 25464 5856 25470 5868
rect 25593 5865 25605 5868
rect 25639 5865 25651 5899
rect 25593 5859 25651 5865
rect 4614 5788 4620 5840
rect 4672 5828 4678 5840
rect 7193 5831 7251 5837
rect 7193 5828 7205 5831
rect 4672 5800 7205 5828
rect 4672 5788 4678 5800
rect 6564 5769 6592 5800
rect 7193 5797 7205 5800
rect 7239 5797 7251 5831
rect 27614 5828 27620 5840
rect 7193 5791 7251 5797
rect 12406 5800 27620 5828
rect 2225 5763 2283 5769
rect 2225 5729 2237 5763
rect 2271 5760 2283 5763
rect 6549 5763 6607 5769
rect 2271 5732 6500 5760
rect 2271 5729 2283 5732
rect 2225 5723 2283 5729
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5692 1731 5695
rect 2240 5692 2268 5723
rect 1719 5664 2268 5692
rect 5537 5695 5595 5701
rect 1719 5661 1731 5664
rect 1673 5655 1731 5661
rect 5537 5661 5549 5695
rect 5583 5692 5595 5695
rect 6362 5692 6368 5704
rect 5583 5664 6368 5692
rect 5583 5661 5595 5664
rect 5537 5655 5595 5661
rect 6362 5652 6368 5664
rect 6420 5652 6426 5704
rect 6472 5692 6500 5732
rect 6549 5729 6561 5763
rect 6595 5760 6607 5763
rect 6595 5732 6629 5760
rect 6595 5729 6607 5732
rect 6549 5723 6607 5729
rect 6472 5664 11744 5692
rect 6457 5627 6515 5633
rect 6457 5593 6469 5627
rect 6503 5624 6515 5627
rect 8478 5624 8484 5636
rect 6503 5596 8484 5624
rect 6503 5593 6515 5596
rect 6457 5587 6515 5593
rect 8478 5584 8484 5596
rect 8536 5584 8542 5636
rect 11716 5624 11744 5664
rect 12406 5624 12434 5800
rect 27614 5788 27620 5800
rect 27672 5788 27678 5840
rect 12802 5720 12808 5772
rect 12860 5760 12866 5772
rect 24946 5760 24952 5772
rect 12860 5732 22094 5760
rect 24907 5732 24952 5760
rect 12860 5720 12866 5732
rect 12986 5692 12992 5704
rect 12947 5664 12992 5692
rect 12986 5652 12992 5664
rect 13044 5652 13050 5704
rect 22066 5692 22094 5732
rect 24946 5720 24952 5732
rect 25004 5760 25010 5772
rect 26326 5760 26332 5772
rect 25004 5732 26332 5760
rect 25004 5720 25010 5732
rect 26326 5720 26332 5732
rect 26384 5760 26390 5772
rect 26605 5763 26663 5769
rect 26605 5760 26617 5763
rect 26384 5732 26617 5760
rect 26384 5720 26390 5732
rect 26605 5729 26617 5732
rect 26651 5729 26663 5763
rect 26605 5723 26663 5729
rect 26694 5692 26700 5704
rect 22066 5664 26700 5692
rect 26694 5652 26700 5664
rect 26752 5652 26758 5704
rect 26881 5695 26939 5701
rect 26881 5661 26893 5695
rect 26927 5692 26939 5695
rect 27614 5692 27620 5704
rect 26927 5664 27620 5692
rect 26927 5661 26939 5664
rect 26881 5655 26939 5661
rect 27614 5652 27620 5664
rect 27672 5652 27678 5704
rect 37826 5692 37832 5704
rect 37787 5664 37832 5692
rect 37826 5652 37832 5664
rect 37884 5652 37890 5704
rect 24765 5627 24823 5633
rect 11716 5596 12434 5624
rect 23768 5596 24532 5624
rect 23768 5568 23796 5596
rect 1486 5556 1492 5568
rect 1447 5528 1492 5556
rect 1486 5516 1492 5528
rect 1544 5516 1550 5568
rect 2777 5559 2835 5565
rect 2777 5525 2789 5559
rect 2823 5556 2835 5559
rect 2958 5556 2964 5568
rect 2823 5528 2964 5556
rect 2823 5525 2835 5528
rect 2777 5519 2835 5525
rect 2958 5516 2964 5528
rect 3016 5516 3022 5568
rect 5810 5516 5816 5568
rect 5868 5556 5874 5568
rect 5997 5559 6055 5565
rect 5997 5556 6009 5559
rect 5868 5528 6009 5556
rect 5868 5516 5874 5528
rect 5997 5525 6009 5528
rect 6043 5525 6055 5559
rect 5997 5519 6055 5525
rect 9582 5516 9588 5568
rect 9640 5556 9646 5568
rect 12805 5559 12863 5565
rect 12805 5556 12817 5559
rect 9640 5528 12817 5556
rect 9640 5516 9646 5528
rect 12805 5525 12817 5528
rect 12851 5525 12863 5559
rect 23750 5556 23756 5568
rect 23711 5528 23756 5556
rect 12805 5519 12863 5525
rect 23750 5516 23756 5528
rect 23808 5516 23814 5568
rect 24394 5556 24400 5568
rect 24355 5528 24400 5556
rect 24394 5516 24400 5528
rect 24452 5516 24458 5568
rect 24504 5556 24532 5596
rect 24765 5593 24777 5627
rect 24811 5624 24823 5627
rect 25406 5624 25412 5636
rect 24811 5596 25412 5624
rect 24811 5593 24823 5596
rect 24765 5587 24823 5593
rect 25406 5584 25412 5596
rect 25464 5584 25470 5636
rect 26789 5627 26847 5633
rect 26789 5593 26801 5627
rect 26835 5624 26847 5627
rect 27801 5627 27859 5633
rect 27801 5624 27813 5627
rect 26835 5596 27813 5624
rect 26835 5593 26847 5596
rect 26789 5587 26847 5593
rect 27801 5593 27813 5596
rect 27847 5624 27859 5627
rect 38194 5624 38200 5636
rect 27847 5596 38200 5624
rect 27847 5593 27859 5596
rect 27801 5587 27859 5593
rect 38194 5584 38200 5596
rect 38252 5584 38258 5636
rect 24857 5559 24915 5565
rect 24857 5556 24869 5559
rect 24504 5528 24869 5556
rect 24857 5525 24869 5528
rect 24903 5525 24915 5559
rect 24857 5519 24915 5525
rect 27062 5516 27068 5568
rect 27120 5556 27126 5568
rect 27249 5559 27307 5565
rect 27249 5556 27261 5559
rect 27120 5528 27261 5556
rect 27120 5516 27126 5528
rect 27249 5525 27261 5528
rect 27295 5525 27307 5559
rect 37366 5556 37372 5568
rect 37327 5528 37372 5556
rect 27249 5519 27307 5525
rect 37366 5516 37372 5528
rect 37424 5516 37430 5568
rect 38010 5556 38016 5568
rect 37971 5528 38016 5556
rect 38010 5516 38016 5528
rect 38068 5516 38074 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5352 1639 5355
rect 6178 5352 6184 5364
rect 1627 5324 6184 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 6178 5312 6184 5324
rect 6236 5312 6242 5364
rect 26326 5352 26332 5364
rect 26287 5324 26332 5352
rect 26326 5312 26332 5324
rect 26384 5312 26390 5364
rect 37369 5355 37427 5361
rect 37369 5321 37381 5355
rect 37415 5352 37427 5355
rect 37826 5352 37832 5364
rect 37415 5324 37832 5352
rect 37415 5321 37427 5324
rect 37369 5315 37427 5321
rect 37826 5312 37832 5324
rect 37884 5352 37890 5364
rect 38470 5352 38476 5364
rect 37884 5324 38476 5352
rect 37884 5312 37890 5324
rect 38470 5312 38476 5324
rect 38528 5312 38534 5364
rect 1394 5216 1400 5228
rect 1355 5188 1400 5216
rect 1394 5176 1400 5188
rect 1452 5216 1458 5228
rect 2041 5219 2099 5225
rect 2041 5216 2053 5219
rect 1452 5188 2053 5216
rect 1452 5176 1458 5188
rect 2041 5185 2053 5188
rect 2087 5185 2099 5219
rect 5810 5216 5816 5228
rect 5771 5188 5816 5216
rect 2041 5179 2099 5185
rect 5810 5176 5816 5188
rect 5868 5176 5874 5228
rect 23661 5219 23719 5225
rect 23661 5185 23673 5219
rect 23707 5216 23719 5219
rect 24394 5216 24400 5228
rect 23707 5188 24400 5216
rect 23707 5185 23719 5188
rect 23661 5179 23719 5185
rect 24394 5176 24400 5188
rect 24452 5176 24458 5228
rect 27062 5216 27068 5228
rect 27023 5188 27068 5216
rect 27062 5176 27068 5188
rect 27120 5176 27126 5228
rect 37734 5176 37740 5228
rect 37792 5216 37798 5228
rect 37829 5219 37887 5225
rect 37829 5216 37841 5219
rect 37792 5188 37841 5216
rect 37792 5176 37798 5188
rect 37829 5185 37841 5188
rect 37875 5185 37887 5219
rect 37829 5179 37887 5185
rect 1670 4972 1676 5024
rect 1728 5012 1734 5024
rect 2593 5015 2651 5021
rect 2593 5012 2605 5015
rect 1728 4984 2605 5012
rect 1728 4972 1734 4984
rect 2593 4981 2605 4984
rect 2639 4981 2651 5015
rect 2593 4975 2651 4981
rect 2866 4972 2872 5024
rect 2924 5012 2930 5024
rect 3145 5015 3203 5021
rect 3145 5012 3157 5015
rect 2924 4984 3157 5012
rect 2924 4972 2930 4984
rect 3145 4981 3157 4984
rect 3191 4981 3203 5015
rect 3145 4975 3203 4981
rect 4798 4972 4804 5024
rect 4856 5012 4862 5024
rect 5629 5015 5687 5021
rect 5629 5012 5641 5015
rect 4856 4984 5641 5012
rect 4856 4972 4862 4984
rect 5629 4981 5641 4984
rect 5675 4981 5687 5015
rect 5629 4975 5687 4981
rect 23845 5015 23903 5021
rect 23845 4981 23857 5015
rect 23891 5012 23903 5015
rect 25590 5012 25596 5024
rect 23891 4984 25596 5012
rect 23891 4981 23903 4984
rect 23845 4975 23903 4981
rect 25590 4972 25596 4984
rect 25648 4972 25654 5024
rect 27249 5015 27307 5021
rect 27249 4981 27261 5015
rect 27295 5012 27307 5015
rect 28902 5012 28908 5024
rect 27295 4984 28908 5012
rect 27295 4981 27307 4984
rect 27249 4975 27307 4981
rect 28902 4972 28908 4984
rect 28960 4972 28966 5024
rect 36630 5012 36636 5024
rect 36591 4984 36636 5012
rect 36630 4972 36636 4984
rect 36688 4972 36694 5024
rect 38010 5012 38016 5024
rect 37971 4984 38016 5012
rect 38010 4972 38016 4984
rect 38068 4972 38074 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 2130 4808 2136 4820
rect 2091 4780 2136 4808
rect 2130 4768 2136 4780
rect 2188 4768 2194 4820
rect 36170 4808 36176 4820
rect 36131 4780 36176 4808
rect 36170 4768 36176 4780
rect 36228 4768 36234 4820
rect 37642 4700 37648 4752
rect 37700 4740 37706 4752
rect 37829 4743 37887 4749
rect 37829 4740 37841 4743
rect 37700 4712 37841 4740
rect 37700 4700 37706 4712
rect 37829 4709 37841 4712
rect 37875 4709 37887 4743
rect 37829 4703 37887 4709
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4604 1731 4607
rect 2130 4604 2136 4616
rect 1719 4576 2136 4604
rect 1719 4573 1731 4576
rect 1673 4567 1731 4573
rect 2130 4564 2136 4576
rect 2188 4564 2194 4616
rect 17589 4607 17647 4613
rect 17589 4573 17601 4607
rect 17635 4604 17647 4607
rect 17954 4604 17960 4616
rect 17635 4576 17960 4604
rect 17635 4573 17647 4576
rect 17589 4567 17647 4573
rect 17954 4564 17960 4576
rect 18012 4564 18018 4616
rect 37369 4539 37427 4545
rect 37369 4505 37381 4539
rect 37415 4536 37427 4539
rect 38010 4536 38016 4548
rect 37415 4508 38016 4536
rect 37415 4505 37427 4508
rect 37369 4499 37427 4505
rect 38010 4496 38016 4508
rect 38068 4496 38074 4548
rect 1486 4468 1492 4480
rect 1447 4440 1492 4468
rect 1486 4428 1492 4440
rect 1544 4428 1550 4480
rect 2774 4468 2780 4480
rect 2735 4440 2780 4468
rect 2774 4428 2780 4440
rect 2832 4428 2838 4480
rect 3878 4468 3884 4480
rect 3839 4440 3884 4468
rect 3878 4428 3884 4440
rect 3936 4428 3942 4480
rect 15562 4468 15568 4480
rect 15523 4440 15568 4468
rect 15562 4428 15568 4440
rect 15620 4428 15626 4480
rect 17773 4471 17831 4477
rect 17773 4437 17785 4471
rect 17819 4468 17831 4471
rect 34790 4468 34796 4480
rect 17819 4440 34796 4468
rect 17819 4437 17831 4440
rect 17773 4431 17831 4437
rect 34790 4428 34796 4440
rect 34848 4428 34854 4480
rect 35710 4468 35716 4480
rect 35671 4440 35716 4468
rect 35710 4428 35716 4440
rect 35768 4428 35774 4480
rect 36722 4468 36728 4480
rect 36683 4440 36728 4468
rect 36722 4428 36728 4440
rect 36780 4428 36786 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 37366 4156 37372 4208
rect 37424 4196 37430 4208
rect 38013 4199 38071 4205
rect 38013 4196 38025 4199
rect 37424 4168 38025 4196
rect 37424 4156 37430 4168
rect 38013 4165 38025 4168
rect 38059 4196 38071 4199
rect 39298 4196 39304 4208
rect 38059 4168 39304 4196
rect 38059 4165 38071 4168
rect 38013 4159 38071 4165
rect 39298 4156 39304 4168
rect 39356 4156 39362 4208
rect 658 4088 664 4140
rect 716 4128 722 4140
rect 1397 4131 1455 4137
rect 1397 4128 1409 4131
rect 716 4100 1409 4128
rect 716 4088 722 4100
rect 1397 4097 1409 4100
rect 1443 4128 1455 4131
rect 1670 4128 1676 4140
rect 1443 4100 1676 4128
rect 1443 4097 1455 4100
rect 1397 4091 1455 4097
rect 1670 4088 1676 4100
rect 1728 4088 1734 4140
rect 2041 4131 2099 4137
rect 2041 4097 2053 4131
rect 2087 4128 2099 4131
rect 2774 4128 2780 4140
rect 2087 4100 2780 4128
rect 2087 4097 2099 4100
rect 2041 4091 2099 4097
rect 2774 4088 2780 4100
rect 2832 4088 2838 4140
rect 3326 4088 3332 4140
rect 3384 4128 3390 4140
rect 10318 4128 10324 4140
rect 3384 4100 10324 4128
rect 3384 4088 3390 4100
rect 10318 4088 10324 4100
rect 10376 4088 10382 4140
rect 13446 4088 13452 4140
rect 13504 4128 13510 4140
rect 18046 4128 18052 4140
rect 13504 4100 18052 4128
rect 13504 4088 13510 4100
rect 18046 4088 18052 4100
rect 18104 4088 18110 4140
rect 24489 4131 24547 4137
rect 24489 4097 24501 4131
rect 24535 4128 24547 4131
rect 24670 4128 24676 4140
rect 24535 4100 24676 4128
rect 24535 4097 24547 4100
rect 24489 4091 24547 4097
rect 24670 4088 24676 4100
rect 24728 4128 24734 4140
rect 26234 4128 26240 4140
rect 24728 4100 26240 4128
rect 24728 4088 24734 4100
rect 26234 4088 26240 4100
rect 26292 4088 26298 4140
rect 30834 4128 30840 4140
rect 30795 4100 30840 4128
rect 30834 4088 30840 4100
rect 30892 4088 30898 4140
rect 37090 4088 37096 4140
rect 37148 4128 37154 4140
rect 37277 4131 37335 4137
rect 37277 4128 37289 4131
rect 37148 4100 37289 4128
rect 37148 4088 37154 4100
rect 37277 4097 37289 4100
rect 37323 4097 37335 4131
rect 37277 4091 37335 4097
rect 1596 4032 9812 4060
rect 1596 4001 1624 4032
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3961 1639 3995
rect 1581 3955 1639 3961
rect 2225 3995 2283 4001
rect 2225 3961 2237 3995
rect 2271 3992 2283 3995
rect 9674 3992 9680 4004
rect 2271 3964 9680 3992
rect 2271 3961 2283 3964
rect 2225 3955 2283 3961
rect 9674 3952 9680 3964
rect 9732 3952 9738 4004
rect 9784 3992 9812 4032
rect 15286 4020 15292 4072
rect 15344 4060 15350 4072
rect 15473 4063 15531 4069
rect 15473 4060 15485 4063
rect 15344 4032 15485 4060
rect 15344 4020 15350 4032
rect 15473 4029 15485 4032
rect 15519 4029 15531 4063
rect 15473 4023 15531 4029
rect 17494 3992 17500 4004
rect 9784 3964 17500 3992
rect 17494 3952 17500 3964
rect 17552 3952 17558 4004
rect 25222 3952 25228 4004
rect 25280 3992 25286 4004
rect 37829 3995 37887 4001
rect 37829 3992 37841 3995
rect 25280 3964 37841 3992
rect 25280 3952 25286 3964
rect 37829 3961 37841 3964
rect 37875 3961 37887 3995
rect 37829 3955 37887 3961
rect 2682 3924 2688 3936
rect 2643 3896 2688 3924
rect 2682 3884 2688 3896
rect 2740 3884 2746 3936
rect 3694 3924 3700 3936
rect 3655 3896 3700 3924
rect 3694 3884 3700 3896
rect 3752 3884 3758 3936
rect 4062 3884 4068 3936
rect 4120 3924 4126 3936
rect 4157 3927 4215 3933
rect 4157 3924 4169 3927
rect 4120 3896 4169 3924
rect 4120 3884 4126 3896
rect 4157 3893 4169 3896
rect 4203 3893 4215 3927
rect 4706 3924 4712 3936
rect 4667 3896 4712 3924
rect 4157 3887 4215 3893
rect 4706 3884 4712 3896
rect 4764 3884 4770 3936
rect 16114 3924 16120 3936
rect 16075 3896 16120 3924
rect 16114 3884 16120 3896
rect 16172 3884 16178 3936
rect 35434 3924 35440 3936
rect 35395 3896 35440 3924
rect 35434 3884 35440 3896
rect 35492 3884 35498 3936
rect 36078 3924 36084 3936
rect 36039 3896 36084 3924
rect 36078 3884 36084 3896
rect 36136 3884 36142 3936
rect 36446 3884 36452 3936
rect 36504 3924 36510 3936
rect 36541 3927 36599 3933
rect 36541 3924 36553 3927
rect 36504 3896 36553 3924
rect 36504 3884 36510 3896
rect 36541 3893 36553 3896
rect 36587 3893 36599 3927
rect 36541 3887 36599 3893
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 3970 3720 3976 3732
rect 3931 3692 3976 3720
rect 3970 3680 3976 3692
rect 4028 3680 4034 3732
rect 5626 3720 5632 3732
rect 5587 3692 5632 3720
rect 5626 3680 5632 3692
rect 5684 3680 5690 3732
rect 13446 3720 13452 3732
rect 13407 3692 13452 3720
rect 13446 3680 13452 3692
rect 13504 3680 13510 3732
rect 14369 3723 14427 3729
rect 14369 3689 14381 3723
rect 14415 3720 14427 3723
rect 14458 3720 14464 3732
rect 14415 3692 14464 3720
rect 14415 3689 14427 3692
rect 14369 3683 14427 3689
rect 14458 3680 14464 3692
rect 14516 3720 14522 3732
rect 17954 3720 17960 3732
rect 14516 3692 16344 3720
rect 17915 3692 17960 3720
rect 14516 3680 14522 3692
rect 2869 3655 2927 3661
rect 2869 3621 2881 3655
rect 2915 3652 2927 3655
rect 4614 3652 4620 3664
rect 2915 3624 4620 3652
rect 2915 3621 2927 3624
rect 2869 3615 2927 3621
rect 4614 3612 4620 3624
rect 4672 3612 4678 3664
rect 16316 3652 16344 3692
rect 17954 3680 17960 3692
rect 18012 3680 18018 3732
rect 18046 3680 18052 3732
rect 18104 3720 18110 3732
rect 26602 3720 26608 3732
rect 18104 3692 26608 3720
rect 18104 3680 18110 3692
rect 26602 3680 26608 3692
rect 26660 3680 26666 3732
rect 30466 3720 30472 3732
rect 30427 3692 30472 3720
rect 30466 3680 30472 3692
rect 30524 3680 30530 3732
rect 31018 3720 31024 3732
rect 30979 3692 31024 3720
rect 31018 3680 31024 3692
rect 31076 3680 31082 3732
rect 33870 3720 33876 3732
rect 33831 3692 33876 3720
rect 33870 3680 33876 3692
rect 33928 3680 33934 3732
rect 16316 3624 18000 3652
rect 1946 3584 1952 3596
rect 1907 3556 1952 3584
rect 1946 3544 1952 3556
rect 2004 3544 2010 3596
rect 2222 3584 2228 3596
rect 2135 3556 2228 3584
rect 2222 3544 2228 3556
rect 2280 3584 2286 3596
rect 4706 3584 4712 3596
rect 2280 3556 4712 3584
rect 2280 3544 2286 3556
rect 4706 3544 4712 3556
rect 4764 3544 4770 3596
rect 13906 3544 13912 3596
rect 13964 3584 13970 3596
rect 15381 3587 15439 3593
rect 15381 3584 15393 3587
rect 13964 3556 15393 3584
rect 13964 3544 13970 3556
rect 15381 3553 15393 3556
rect 15427 3553 15439 3587
rect 17310 3584 17316 3596
rect 17271 3556 17316 3584
rect 15381 3547 15439 3553
rect 17310 3544 17316 3556
rect 17368 3544 17374 3596
rect 17494 3584 17500 3596
rect 17455 3556 17500 3584
rect 17494 3544 17500 3556
rect 17552 3544 17558 3596
rect 17972 3584 18000 3624
rect 18414 3612 18420 3664
rect 18472 3652 18478 3664
rect 24670 3652 24676 3664
rect 18472 3624 24676 3652
rect 18472 3612 18478 3624
rect 24670 3612 24676 3624
rect 24728 3612 24734 3664
rect 33318 3612 33324 3664
rect 33376 3652 33382 3664
rect 35713 3655 35771 3661
rect 35713 3652 35725 3655
rect 33376 3624 35725 3652
rect 33376 3612 33382 3624
rect 35713 3621 35725 3624
rect 35759 3621 35771 3655
rect 35713 3615 35771 3621
rect 37277 3655 37335 3661
rect 37277 3621 37289 3655
rect 37323 3652 37335 3655
rect 38654 3652 38660 3664
rect 37323 3624 38660 3652
rect 37323 3621 37335 3624
rect 37277 3615 37335 3621
rect 38654 3612 38660 3624
rect 38712 3612 38718 3664
rect 22738 3584 22744 3596
rect 17972 3556 22744 3584
rect 22738 3544 22744 3556
rect 22796 3544 22802 3596
rect 24762 3544 24768 3596
rect 24820 3584 24826 3596
rect 36538 3584 36544 3596
rect 24820 3556 36544 3584
rect 24820 3544 24826 3556
rect 36538 3544 36544 3556
rect 36596 3544 36602 3596
rect 2682 3516 2688 3528
rect 1964 3488 2688 3516
rect 1964 3460 1992 3488
rect 2682 3476 2688 3488
rect 2740 3476 2746 3528
rect 3694 3476 3700 3528
rect 3752 3516 3758 3528
rect 3789 3519 3847 3525
rect 3789 3516 3801 3519
rect 3752 3488 3801 3516
rect 3752 3476 3758 3488
rect 3789 3485 3801 3488
rect 3835 3485 3847 3519
rect 3789 3479 3847 3485
rect 1946 3408 1952 3460
rect 2004 3408 2010 3460
rect 2590 3408 2596 3460
rect 2648 3448 2654 3460
rect 3804 3448 3832 3479
rect 9490 3476 9496 3528
rect 9548 3516 9554 3528
rect 14366 3516 14372 3528
rect 9548 3488 14372 3516
rect 9548 3476 9554 3488
rect 14366 3476 14372 3488
rect 14424 3476 14430 3528
rect 15648 3519 15706 3525
rect 15648 3485 15660 3519
rect 15694 3516 15706 3519
rect 16114 3516 16120 3528
rect 15694 3488 16120 3516
rect 15694 3485 15706 3488
rect 15648 3479 15706 3485
rect 16114 3476 16120 3488
rect 16172 3476 16178 3528
rect 24581 3519 24639 3525
rect 24581 3516 24593 3519
rect 17420 3488 24593 3516
rect 2648 3420 3832 3448
rect 2648 3408 2654 3420
rect 4614 3340 4620 3392
rect 4672 3380 4678 3392
rect 4893 3383 4951 3389
rect 4893 3380 4905 3383
rect 4672 3352 4905 3380
rect 4672 3340 4678 3352
rect 4893 3349 4905 3352
rect 4939 3349 4951 3383
rect 6178 3380 6184 3392
rect 6139 3352 6184 3380
rect 4893 3343 4951 3349
rect 6178 3340 6184 3352
rect 6236 3340 6242 3392
rect 11606 3380 11612 3392
rect 11567 3352 11612 3380
rect 11606 3340 11612 3352
rect 11664 3340 11670 3392
rect 14918 3380 14924 3392
rect 14879 3352 14924 3380
rect 14918 3340 14924 3352
rect 14976 3340 14982 3392
rect 16761 3383 16819 3389
rect 16761 3349 16773 3383
rect 16807 3380 16819 3383
rect 17420 3380 17448 3488
rect 24581 3485 24593 3488
rect 24627 3485 24639 3519
rect 24581 3479 24639 3485
rect 27706 3476 27712 3528
rect 27764 3516 27770 3528
rect 28445 3519 28503 3525
rect 28445 3516 28457 3519
rect 27764 3488 28457 3516
rect 27764 3476 27770 3488
rect 28445 3485 28457 3488
rect 28491 3485 28503 3519
rect 28445 3479 28503 3485
rect 30926 3476 30932 3528
rect 30984 3516 30990 3528
rect 31205 3519 31263 3525
rect 31205 3516 31217 3519
rect 30984 3488 31217 3516
rect 30984 3476 30990 3488
rect 31205 3485 31217 3488
rect 31251 3516 31263 3519
rect 31665 3519 31723 3525
rect 31665 3516 31677 3519
rect 31251 3488 31677 3516
rect 31251 3485 31263 3488
rect 31205 3479 31263 3485
rect 31665 3485 31677 3488
rect 31711 3485 31723 3519
rect 31665 3479 31723 3485
rect 35897 3519 35955 3525
rect 35897 3485 35909 3519
rect 35943 3516 35955 3519
rect 36078 3516 36084 3528
rect 35943 3488 36084 3516
rect 35943 3485 35955 3488
rect 35897 3479 35955 3485
rect 36078 3476 36084 3488
rect 36136 3476 36142 3528
rect 36357 3519 36415 3525
rect 36357 3485 36369 3519
rect 36403 3485 36415 3519
rect 37090 3516 37096 3528
rect 37051 3488 37096 3516
rect 36357 3479 36415 3485
rect 17494 3408 17500 3460
rect 17552 3448 17558 3460
rect 18414 3448 18420 3460
rect 17552 3420 18420 3448
rect 17552 3408 17558 3420
rect 18414 3408 18420 3420
rect 18472 3408 18478 3460
rect 25958 3408 25964 3460
rect 26016 3448 26022 3460
rect 36372 3448 36400 3479
rect 37090 3476 37096 3488
rect 37148 3476 37154 3528
rect 37826 3516 37832 3528
rect 37787 3488 37832 3516
rect 37826 3476 37832 3488
rect 37884 3476 37890 3528
rect 26016 3420 36400 3448
rect 26016 3408 26022 3420
rect 16807 3352 17448 3380
rect 16807 3349 16819 3352
rect 16761 3343 16819 3349
rect 17586 3340 17592 3392
rect 17644 3380 17650 3392
rect 17644 3352 17689 3380
rect 17644 3340 17650 3352
rect 21082 3340 21088 3392
rect 21140 3380 21146 3392
rect 21361 3383 21419 3389
rect 21361 3380 21373 3383
rect 21140 3352 21373 3380
rect 21140 3340 21146 3352
rect 21361 3349 21373 3352
rect 21407 3349 21419 3383
rect 23198 3380 23204 3392
rect 23159 3352 23204 3380
rect 21361 3343 21419 3349
rect 23198 3340 23204 3352
rect 23256 3340 23262 3392
rect 23658 3380 23664 3392
rect 23619 3352 23664 3380
rect 23658 3340 23664 3352
rect 23716 3340 23722 3392
rect 24486 3340 24492 3392
rect 24544 3380 24550 3392
rect 24765 3383 24823 3389
rect 24765 3380 24777 3383
rect 24544 3352 24777 3380
rect 24544 3340 24550 3352
rect 24765 3349 24777 3352
rect 24811 3349 24823 3383
rect 24765 3343 24823 3349
rect 26418 3340 26424 3392
rect 26476 3380 26482 3392
rect 26789 3383 26847 3389
rect 26789 3380 26801 3383
rect 26476 3352 26801 3380
rect 26476 3340 26482 3352
rect 26789 3349 26801 3352
rect 26835 3349 26847 3383
rect 26789 3343 26847 3349
rect 27154 3340 27160 3392
rect 27212 3380 27218 3392
rect 27341 3383 27399 3389
rect 27341 3380 27353 3383
rect 27212 3352 27353 3380
rect 27212 3340 27218 3352
rect 27341 3349 27353 3352
rect 27387 3349 27399 3383
rect 27341 3343 27399 3349
rect 27522 3340 27528 3392
rect 27580 3380 27586 3392
rect 27893 3383 27951 3389
rect 27893 3380 27905 3383
rect 27580 3352 27905 3380
rect 27580 3340 27586 3352
rect 27893 3349 27905 3352
rect 27939 3349 27951 3383
rect 27893 3343 27951 3349
rect 28902 3340 28908 3392
rect 28960 3380 28966 3392
rect 32030 3380 32036 3392
rect 28960 3352 32036 3380
rect 28960 3340 28966 3352
rect 32030 3340 32036 3352
rect 32088 3340 32094 3392
rect 32214 3380 32220 3392
rect 32175 3352 32220 3380
rect 32214 3340 32220 3352
rect 32272 3340 32278 3392
rect 32766 3380 32772 3392
rect 32727 3352 32772 3380
rect 32766 3340 32772 3352
rect 32824 3340 32830 3392
rect 32858 3340 32864 3392
rect 32916 3380 32922 3392
rect 33321 3383 33379 3389
rect 33321 3380 33333 3383
rect 32916 3352 33333 3380
rect 32916 3340 32922 3352
rect 33321 3349 33333 3352
rect 33367 3349 33379 3383
rect 33321 3343 33379 3349
rect 34146 3340 34152 3392
rect 34204 3380 34210 3392
rect 34701 3383 34759 3389
rect 34701 3380 34713 3383
rect 34204 3352 34713 3380
rect 34204 3340 34210 3352
rect 34701 3349 34713 3352
rect 34747 3349 34759 3383
rect 34701 3343 34759 3349
rect 36541 3383 36599 3389
rect 36541 3349 36553 3383
rect 36587 3380 36599 3383
rect 36814 3380 36820 3392
rect 36587 3352 36820 3380
rect 36587 3349 36599 3352
rect 36541 3343 36599 3349
rect 36814 3340 36820 3352
rect 36872 3340 36878 3392
rect 38010 3380 38016 3392
rect 37971 3352 38016 3380
rect 38010 3340 38016 3352
rect 38068 3340 38074 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 2314 3176 2320 3188
rect 2275 3148 2320 3176
rect 2314 3136 2320 3148
rect 2372 3136 2378 3188
rect 8478 3176 8484 3188
rect 8439 3148 8484 3176
rect 8478 3136 8484 3148
rect 8536 3136 8542 3188
rect 9766 3176 9772 3188
rect 9727 3148 9772 3176
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 10410 3176 10416 3188
rect 10371 3148 10416 3176
rect 10410 3136 10416 3148
rect 10468 3136 10474 3188
rect 11701 3179 11759 3185
rect 11701 3145 11713 3179
rect 11747 3176 11759 3179
rect 12710 3176 12716 3188
rect 11747 3148 12716 3176
rect 11747 3145 11759 3148
rect 11701 3139 11759 3145
rect 12710 3136 12716 3148
rect 12768 3136 12774 3188
rect 13173 3179 13231 3185
rect 13173 3145 13185 3179
rect 13219 3176 13231 3179
rect 15286 3176 15292 3188
rect 13219 3148 15148 3176
rect 15247 3148 15292 3176
rect 13219 3145 13231 3148
rect 13173 3139 13231 3145
rect 14 3068 20 3120
rect 72 3108 78 3120
rect 3145 3111 3203 3117
rect 72 3080 3096 3108
rect 72 3068 78 3080
rect 2225 3043 2283 3049
rect 2225 3009 2237 3043
rect 2271 3040 2283 3043
rect 2866 3040 2872 3052
rect 2271 3012 2872 3040
rect 2271 3009 2283 3012
rect 2225 3003 2283 3009
rect 2866 3000 2872 3012
rect 2924 3000 2930 3052
rect 2961 3043 3019 3049
rect 2961 3009 2973 3043
rect 3007 3009 3019 3043
rect 3068 3040 3096 3080
rect 3145 3077 3157 3111
rect 3191 3108 3203 3111
rect 3234 3108 3240 3120
rect 3191 3080 3240 3108
rect 3191 3077 3203 3080
rect 3145 3071 3203 3077
rect 3234 3068 3240 3080
rect 3292 3068 3298 3120
rect 4801 3111 4859 3117
rect 4801 3077 4813 3111
rect 4847 3108 4859 3111
rect 9490 3108 9496 3120
rect 4847 3080 9496 3108
rect 4847 3077 4859 3080
rect 4801 3071 4859 3077
rect 9490 3068 9496 3080
rect 9548 3068 9554 3120
rect 9674 3068 9680 3120
rect 9732 3108 9738 3120
rect 14154 3111 14212 3117
rect 14154 3108 14166 3111
rect 9732 3080 14166 3108
rect 9732 3068 9738 3080
rect 14154 3077 14166 3080
rect 14200 3077 14212 3111
rect 15120 3108 15148 3148
rect 15286 3136 15292 3148
rect 15344 3136 15350 3188
rect 17497 3179 17555 3185
rect 17497 3145 17509 3179
rect 17543 3176 17555 3179
rect 17586 3176 17592 3188
rect 17543 3148 17592 3176
rect 17543 3145 17555 3148
rect 17497 3139 17555 3145
rect 17586 3136 17592 3148
rect 17644 3136 17650 3188
rect 17770 3136 17776 3188
rect 17828 3176 17834 3188
rect 18785 3179 18843 3185
rect 18785 3176 18797 3179
rect 17828 3148 18797 3176
rect 17828 3136 17834 3148
rect 18785 3145 18797 3148
rect 18831 3145 18843 3179
rect 20530 3176 20536 3188
rect 20491 3148 20536 3176
rect 18785 3139 18843 3145
rect 20530 3136 20536 3148
rect 20588 3136 20594 3188
rect 21269 3179 21327 3185
rect 21269 3145 21281 3179
rect 21315 3176 21327 3179
rect 24949 3179 25007 3185
rect 24949 3176 24961 3179
rect 21315 3148 24961 3176
rect 21315 3145 21327 3148
rect 21269 3139 21327 3145
rect 24949 3145 24961 3148
rect 24995 3145 25007 3179
rect 25958 3176 25964 3188
rect 25919 3148 25964 3176
rect 24949 3139 25007 3145
rect 25958 3136 25964 3148
rect 26016 3136 26022 3188
rect 26970 3176 26976 3188
rect 26931 3148 26976 3176
rect 26970 3136 26976 3148
rect 27028 3136 27034 3188
rect 27430 3136 27436 3188
rect 27488 3176 27494 3188
rect 27617 3179 27675 3185
rect 27617 3176 27629 3179
rect 27488 3148 27629 3176
rect 27488 3136 27494 3148
rect 27617 3145 27629 3148
rect 27663 3145 27675 3179
rect 27617 3139 27675 3145
rect 28350 3136 28356 3188
rect 28408 3176 28414 3188
rect 28445 3179 28503 3185
rect 28445 3176 28457 3179
rect 28408 3148 28457 3176
rect 28408 3136 28414 3148
rect 28445 3145 28457 3148
rect 28491 3145 28503 3179
rect 28445 3139 28503 3145
rect 31573 3179 31631 3185
rect 31573 3145 31585 3179
rect 31619 3145 31631 3179
rect 31573 3139 31631 3145
rect 30377 3111 30435 3117
rect 30377 3108 30389 3111
rect 15120 3080 30389 3108
rect 14154 3071 14212 3077
rect 30377 3077 30389 3080
rect 30423 3108 30435 3111
rect 31205 3111 31263 3117
rect 31205 3108 31217 3111
rect 30423 3080 31217 3108
rect 30423 3077 30435 3080
rect 30377 3071 30435 3077
rect 31205 3077 31217 3080
rect 31251 3077 31263 3111
rect 31205 3071 31263 3077
rect 3605 3043 3663 3049
rect 3605 3040 3617 3043
rect 3068 3012 3617 3040
rect 2961 3003 3019 3009
rect 3605 3009 3617 3012
rect 3651 3040 3663 3043
rect 4062 3040 4068 3052
rect 3651 3012 4068 3040
rect 3651 3009 3663 3012
rect 3605 3003 3663 3009
rect 2976 2972 3004 3003
rect 4062 3000 4068 3012
rect 4120 3000 4126 3052
rect 4614 3040 4620 3052
rect 4575 3012 4620 3040
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 5537 3043 5595 3049
rect 5537 3009 5549 3043
rect 5583 3040 5595 3043
rect 5626 3040 5632 3052
rect 5583 3012 5632 3040
rect 5583 3009 5595 3012
rect 5537 3003 5595 3009
rect 5626 3000 5632 3012
rect 5684 3000 5690 3052
rect 6733 3043 6791 3049
rect 6733 3009 6745 3043
rect 6779 3040 6791 3043
rect 7098 3040 7104 3052
rect 6779 3012 7104 3040
rect 6779 3009 6791 3012
rect 6733 3003 6791 3009
rect 7098 3000 7104 3012
rect 7156 3040 7162 3052
rect 7193 3043 7251 3049
rect 7193 3040 7205 3043
rect 7156 3012 7205 3040
rect 7156 3000 7162 3012
rect 7193 3009 7205 3012
rect 7239 3009 7251 3043
rect 7193 3003 7251 3009
rect 8386 3000 8392 3052
rect 8444 3040 8450 3052
rect 8665 3043 8723 3049
rect 8665 3040 8677 3043
rect 8444 3012 8677 3040
rect 8444 3000 8450 3012
rect 8665 3009 8677 3012
rect 8711 3009 8723 3043
rect 8665 3003 8723 3009
rect 10962 3000 10968 3052
rect 11020 3040 11026 3052
rect 11517 3043 11575 3049
rect 11517 3040 11529 3043
rect 11020 3012 11529 3040
rect 11020 3000 11026 3012
rect 11517 3009 11529 3012
rect 11563 3009 11575 3043
rect 11517 3003 11575 3009
rect 12529 3043 12587 3049
rect 12529 3009 12541 3043
rect 12575 3040 12587 3043
rect 12894 3040 12900 3052
rect 12575 3012 12900 3040
rect 12575 3009 12587 3012
rect 12529 3003 12587 3009
rect 12894 3000 12900 3012
rect 12952 3040 12958 3052
rect 12989 3043 13047 3049
rect 12989 3040 13001 3043
rect 12952 3012 13001 3040
rect 12952 3000 12958 3012
rect 12989 3009 13001 3012
rect 13035 3009 13047 3043
rect 13906 3040 13912 3052
rect 13867 3012 13912 3040
rect 12989 3003 13047 3009
rect 13906 3000 13912 3012
rect 13964 3000 13970 3052
rect 14918 3000 14924 3052
rect 14976 3040 14982 3052
rect 15749 3043 15807 3049
rect 15749 3040 15761 3043
rect 14976 3012 15761 3040
rect 14976 3000 14982 3012
rect 15749 3009 15761 3012
rect 15795 3009 15807 3043
rect 15749 3003 15807 3009
rect 17402 3000 17408 3052
rect 17460 3040 17466 3052
rect 17681 3043 17739 3049
rect 17681 3040 17693 3043
rect 17460 3012 17693 3040
rect 17460 3000 17466 3012
rect 17681 3009 17693 3012
rect 17727 3040 17739 3043
rect 18141 3043 18199 3049
rect 18141 3040 18153 3043
rect 17727 3012 18153 3040
rect 17727 3009 17739 3012
rect 17681 3003 17739 3009
rect 18141 3009 18153 3012
rect 18187 3009 18199 3043
rect 18141 3003 18199 3009
rect 18690 3000 18696 3052
rect 18748 3040 18754 3052
rect 18969 3043 19027 3049
rect 18969 3040 18981 3043
rect 18748 3012 18981 3040
rect 18748 3000 18754 3012
rect 18969 3009 18981 3012
rect 19015 3040 19027 3043
rect 19429 3043 19487 3049
rect 19429 3040 19441 3043
rect 19015 3012 19441 3040
rect 19015 3009 19027 3012
rect 18969 3003 19027 3009
rect 19429 3009 19441 3012
rect 19475 3009 19487 3043
rect 21082 3040 21088 3052
rect 21043 3012 21088 3040
rect 19429 3003 19487 3009
rect 21082 3000 21088 3012
rect 21140 3000 21146 3052
rect 22097 3043 22155 3049
rect 22097 3009 22109 3043
rect 22143 3040 22155 3043
rect 24394 3040 24400 3052
rect 22143 3012 24400 3040
rect 22143 3009 22155 3012
rect 22097 3003 22155 3009
rect 24394 3000 24400 3012
rect 24452 3000 24458 3052
rect 25777 3043 25835 3049
rect 25777 3040 25789 3043
rect 25332 3012 25789 3040
rect 12250 2972 12256 2984
rect 1596 2944 3004 2972
rect 6886 2944 12256 2972
rect 1302 2796 1308 2848
rect 1360 2836 1366 2848
rect 1596 2845 1624 2944
rect 3789 2907 3847 2913
rect 3789 2873 3801 2907
rect 3835 2904 3847 2907
rect 6886 2904 6914 2944
rect 12250 2932 12256 2944
rect 12308 2932 12314 2984
rect 21450 2932 21456 2984
rect 21508 2972 21514 2984
rect 21508 2944 22094 2972
rect 21508 2932 21514 2944
rect 3835 2876 6914 2904
rect 7377 2907 7435 2913
rect 3835 2873 3847 2876
rect 3789 2867 3847 2873
rect 7377 2873 7389 2907
rect 7423 2904 7435 2907
rect 11974 2904 11980 2916
rect 7423 2876 11980 2904
rect 7423 2873 7435 2876
rect 7377 2867 7435 2873
rect 11974 2864 11980 2876
rect 12032 2864 12038 2916
rect 15933 2907 15991 2913
rect 15933 2873 15945 2907
rect 15979 2904 15991 2907
rect 21542 2904 21548 2916
rect 15979 2876 21548 2904
rect 15979 2873 15991 2876
rect 15933 2867 15991 2873
rect 21542 2864 21548 2876
rect 21600 2864 21606 2916
rect 22066 2904 22094 2944
rect 23198 2932 23204 2984
rect 23256 2972 23262 2984
rect 23293 2975 23351 2981
rect 23293 2972 23305 2975
rect 23256 2944 23305 2972
rect 23256 2932 23262 2944
rect 23293 2941 23305 2944
rect 23339 2941 23351 2975
rect 23293 2935 23351 2941
rect 23569 2975 23627 2981
rect 23569 2941 23581 2975
rect 23615 2941 23627 2975
rect 24670 2972 24676 2984
rect 24631 2944 24676 2972
rect 23569 2935 23627 2941
rect 23584 2904 23612 2935
rect 24670 2932 24676 2944
rect 24728 2932 24734 2984
rect 24857 2975 24915 2981
rect 24857 2941 24869 2975
rect 24903 2941 24915 2975
rect 24857 2935 24915 2941
rect 22066 2876 23612 2904
rect 1581 2839 1639 2845
rect 1581 2836 1593 2839
rect 1360 2808 1593 2836
rect 1360 2796 1366 2808
rect 1581 2805 1593 2808
rect 1627 2805 1639 2839
rect 1581 2799 1639 2805
rect 5166 2796 5172 2848
rect 5224 2836 5230 2848
rect 5353 2839 5411 2845
rect 5353 2836 5365 2839
rect 5224 2808 5365 2836
rect 5224 2796 5230 2808
rect 5353 2805 5365 2808
rect 5399 2805 5411 2839
rect 5353 2799 5411 2805
rect 8021 2839 8079 2845
rect 8021 2805 8033 2839
rect 8067 2836 8079 2839
rect 8386 2836 8392 2848
rect 8067 2808 8392 2836
rect 8067 2805 8079 2808
rect 8021 2799 8079 2805
rect 8386 2796 8392 2808
rect 8444 2796 8450 2848
rect 9030 2796 9036 2848
rect 9088 2836 9094 2848
rect 9217 2839 9275 2845
rect 9217 2836 9229 2839
rect 9088 2808 9229 2836
rect 9088 2796 9094 2808
rect 9217 2805 9229 2808
rect 9263 2805 9275 2839
rect 10962 2836 10968 2848
rect 10923 2808 10968 2836
rect 9217 2799 9275 2805
rect 10962 2796 10968 2808
rect 11020 2796 11026 2848
rect 16114 2796 16120 2848
rect 16172 2836 16178 2848
rect 16669 2839 16727 2845
rect 16669 2836 16681 2839
rect 16172 2808 16681 2836
rect 16172 2796 16178 2808
rect 16669 2805 16681 2808
rect 16715 2805 16727 2839
rect 21910 2836 21916 2848
rect 21871 2808 21916 2836
rect 16669 2799 16727 2805
rect 21910 2796 21916 2808
rect 21968 2796 21974 2848
rect 22002 2796 22008 2848
rect 22060 2836 22066 2848
rect 22557 2839 22615 2845
rect 22557 2836 22569 2839
rect 22060 2808 22569 2836
rect 22060 2796 22066 2808
rect 22557 2805 22569 2808
rect 22603 2805 22615 2839
rect 24872 2836 24900 2935
rect 25332 2913 25360 3012
rect 25777 3009 25789 3012
rect 25823 3009 25835 3043
rect 25777 3003 25835 3009
rect 26418 3000 26424 3052
rect 26476 3040 26482 3052
rect 27157 3043 27215 3049
rect 27157 3040 27169 3043
rect 26476 3012 27169 3040
rect 26476 3000 26482 3012
rect 27157 3009 27169 3012
rect 27203 3009 27215 3043
rect 27157 3003 27215 3009
rect 27801 3043 27859 3049
rect 27801 3009 27813 3043
rect 27847 3009 27859 3043
rect 27801 3003 27859 3009
rect 27062 2932 27068 2984
rect 27120 2972 27126 2984
rect 27522 2972 27528 2984
rect 27120 2944 27528 2972
rect 27120 2932 27126 2944
rect 27522 2932 27528 2944
rect 27580 2972 27586 2984
rect 27816 2972 27844 3003
rect 28534 3000 28540 3052
rect 28592 3040 28598 3052
rect 28629 3043 28687 3049
rect 28629 3040 28641 3043
rect 28592 3012 28641 3040
rect 28592 3000 28598 3012
rect 28629 3009 28641 3012
rect 28675 3040 28687 3043
rect 29089 3043 29147 3049
rect 29089 3040 29101 3043
rect 28675 3012 29101 3040
rect 28675 3009 28687 3012
rect 28629 3003 28687 3009
rect 29089 3009 29101 3012
rect 29135 3009 29147 3043
rect 31588 3040 31616 3139
rect 31662 3136 31668 3188
rect 31720 3176 31726 3188
rect 33413 3179 33471 3185
rect 33413 3176 33425 3179
rect 31720 3148 33425 3176
rect 31720 3136 31726 3148
rect 33413 3145 33425 3148
rect 33459 3145 33471 3179
rect 33413 3139 33471 3145
rect 34425 3179 34483 3185
rect 34425 3145 34437 3179
rect 34471 3176 34483 3179
rect 34606 3176 34612 3188
rect 34471 3148 34612 3176
rect 34471 3145 34483 3148
rect 34425 3139 34483 3145
rect 34606 3136 34612 3148
rect 34664 3136 34670 3188
rect 36538 3176 36544 3188
rect 36499 3148 36544 3176
rect 36538 3136 36544 3148
rect 36596 3136 36602 3188
rect 32030 3068 32036 3120
rect 32088 3108 32094 3120
rect 32088 3080 35756 3108
rect 32088 3068 32094 3080
rect 32125 3043 32183 3049
rect 32125 3040 32137 3043
rect 31588 3012 32137 3040
rect 29089 3003 29147 3009
rect 32125 3009 32137 3012
rect 32171 3009 32183 3043
rect 32125 3003 32183 3009
rect 32306 3000 32312 3052
rect 32364 3040 32370 3052
rect 32766 3040 32772 3052
rect 32364 3012 32772 3040
rect 32364 3000 32370 3012
rect 32766 3000 32772 3012
rect 32824 3040 32830 3052
rect 32953 3043 33011 3049
rect 32953 3040 32965 3043
rect 32824 3012 32965 3040
rect 32824 3000 32830 3012
rect 32953 3009 32965 3012
rect 32999 3009 33011 3043
rect 32953 3003 33011 3009
rect 33597 3043 33655 3049
rect 33597 3009 33609 3043
rect 33643 3009 33655 3043
rect 33597 3003 33655 3009
rect 27580 2944 27844 2972
rect 27580 2932 27586 2944
rect 30466 2932 30472 2984
rect 30524 2972 30530 2984
rect 30929 2975 30987 2981
rect 30929 2972 30941 2975
rect 30524 2944 30941 2972
rect 30524 2932 30530 2944
rect 30929 2941 30941 2944
rect 30975 2941 30987 2975
rect 30929 2935 30987 2941
rect 31113 2975 31171 2981
rect 31113 2941 31125 2975
rect 31159 2941 31171 2975
rect 31113 2935 31171 2941
rect 25317 2907 25375 2913
rect 25317 2873 25329 2907
rect 25363 2873 25375 2907
rect 25317 2867 25375 2873
rect 27798 2836 27804 2848
rect 24872 2808 27804 2836
rect 22557 2799 22615 2805
rect 27798 2796 27804 2808
rect 27856 2796 27862 2848
rect 29638 2836 29644 2848
rect 29599 2808 29644 2836
rect 29638 2796 29644 2808
rect 29696 2796 29702 2848
rect 31128 2836 31156 2935
rect 32858 2932 32864 2984
rect 32916 2972 32922 2984
rect 33612 2972 33640 3003
rect 34146 3000 34152 3052
rect 34204 3040 34210 3052
rect 34241 3043 34299 3049
rect 34241 3040 34253 3043
rect 34204 3012 34253 3040
rect 34204 3000 34210 3012
rect 34241 3009 34253 3012
rect 34287 3009 34299 3043
rect 34241 3003 34299 3009
rect 35253 3043 35311 3049
rect 35253 3009 35265 3043
rect 35299 3040 35311 3043
rect 35434 3040 35440 3052
rect 35299 3012 35440 3040
rect 35299 3009 35311 3012
rect 35253 3003 35311 3009
rect 35434 3000 35440 3012
rect 35492 3000 35498 3052
rect 35728 3049 35756 3080
rect 36170 3068 36176 3120
rect 36228 3108 36234 3120
rect 36228 3080 37504 3108
rect 36228 3068 36234 3080
rect 37476 3049 37504 3080
rect 35713 3043 35771 3049
rect 35713 3009 35725 3043
rect 35759 3009 35771 3043
rect 35713 3003 35771 3009
rect 36633 3043 36691 3049
rect 36633 3009 36645 3043
rect 36679 3009 36691 3043
rect 36633 3003 36691 3009
rect 37461 3043 37519 3049
rect 37461 3009 37473 3043
rect 37507 3009 37519 3043
rect 37461 3003 37519 3009
rect 36648 2972 36676 3003
rect 36722 2972 36728 2984
rect 32916 2944 33640 2972
rect 36635 2944 36728 2972
rect 32916 2932 32922 2944
rect 36722 2932 36728 2944
rect 36780 2972 36786 2984
rect 37918 2972 37924 2984
rect 36780 2944 37924 2972
rect 36780 2932 36786 2944
rect 37918 2932 37924 2944
rect 37976 2932 37982 2984
rect 32769 2907 32827 2913
rect 32769 2904 32781 2907
rect 31680 2876 32781 2904
rect 31680 2836 31708 2876
rect 32769 2873 32781 2876
rect 32815 2873 32827 2907
rect 34790 2904 34796 2916
rect 32769 2867 32827 2873
rect 33336 2876 34796 2904
rect 31128 2808 31708 2836
rect 32309 2839 32367 2845
rect 32309 2805 32321 2839
rect 32355 2836 32367 2839
rect 33336 2836 33364 2876
rect 34790 2864 34796 2876
rect 34848 2864 34854 2916
rect 32355 2808 33364 2836
rect 32355 2805 32367 2808
rect 32309 2799 32367 2805
rect 34514 2796 34520 2848
rect 34572 2836 34578 2848
rect 35069 2839 35127 2845
rect 35069 2836 35081 2839
rect 34572 2808 35081 2836
rect 34572 2796 34578 2808
rect 35069 2805 35081 2808
rect 35115 2805 35127 2839
rect 35069 2799 35127 2805
rect 35894 2796 35900 2848
rect 35952 2836 35958 2848
rect 35952 2808 35997 2836
rect 35952 2796 35958 2808
rect 37366 2796 37372 2848
rect 37424 2836 37430 2848
rect 37645 2839 37703 2845
rect 37645 2836 37657 2839
rect 37424 2808 37657 2836
rect 37424 2796 37430 2808
rect 37645 2805 37657 2808
rect 37691 2805 37703 2839
rect 37645 2799 37703 2805
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 8018 2632 8024 2644
rect 7979 2604 8024 2632
rect 8018 2592 8024 2604
rect 8076 2592 8082 2644
rect 9122 2632 9128 2644
rect 9083 2604 9128 2632
rect 9122 2592 9128 2604
rect 9180 2592 9186 2644
rect 15470 2632 15476 2644
rect 15431 2604 15476 2632
rect 15470 2592 15476 2604
rect 15528 2592 15534 2644
rect 15930 2632 15936 2644
rect 15891 2604 15936 2632
rect 15930 2592 15936 2604
rect 15988 2592 15994 2644
rect 23750 2632 23756 2644
rect 16040 2604 23756 2632
rect 16040 2564 16068 2604
rect 23750 2592 23756 2604
rect 23808 2592 23814 2644
rect 24394 2632 24400 2644
rect 24355 2604 24400 2632
rect 24394 2592 24400 2604
rect 24452 2592 24458 2644
rect 26694 2592 26700 2644
rect 26752 2632 26758 2644
rect 26973 2635 27031 2641
rect 26973 2632 26985 2635
rect 26752 2604 26985 2632
rect 26752 2592 26758 2604
rect 26973 2601 26985 2604
rect 27019 2601 27031 2635
rect 27614 2632 27620 2644
rect 27575 2604 27620 2632
rect 26973 2595 27031 2601
rect 27614 2592 27620 2604
rect 27672 2592 27678 2644
rect 27798 2592 27804 2644
rect 27856 2632 27862 2644
rect 28261 2635 28319 2641
rect 28261 2632 28273 2635
rect 27856 2604 28273 2632
rect 27856 2592 27862 2604
rect 28261 2601 28273 2604
rect 28307 2601 28319 2635
rect 28261 2595 28319 2601
rect 28442 2592 28448 2644
rect 28500 2632 28506 2644
rect 34514 2632 34520 2644
rect 28500 2604 34520 2632
rect 28500 2592 28506 2604
rect 34514 2592 34520 2604
rect 34572 2592 34578 2644
rect 35802 2632 35808 2644
rect 35763 2604 35808 2632
rect 35802 2592 35808 2604
rect 35860 2592 35866 2644
rect 18598 2564 18604 2576
rect 1964 2536 16068 2564
rect 16546 2536 18604 2564
rect 1964 2505 1992 2536
rect 1949 2499 2007 2505
rect 1949 2465 1961 2499
rect 1995 2465 2007 2499
rect 1949 2459 2007 2465
rect 3878 2456 3884 2508
rect 3936 2496 3942 2508
rect 3973 2499 4031 2505
rect 3973 2496 3985 2499
rect 3936 2468 3985 2496
rect 3936 2456 3942 2468
rect 3973 2465 3985 2468
rect 4019 2465 4031 2499
rect 3973 2459 4031 2465
rect 4249 2499 4307 2505
rect 4249 2465 4261 2499
rect 4295 2496 4307 2499
rect 10502 2496 10508 2508
rect 4295 2468 10508 2496
rect 4295 2465 4307 2468
rect 4249 2459 4307 2465
rect 10502 2456 10508 2468
rect 10560 2456 10566 2508
rect 11977 2499 12035 2505
rect 11977 2465 11989 2499
rect 12023 2496 12035 2499
rect 16546 2496 16574 2536
rect 18598 2524 18604 2536
rect 18656 2524 18662 2576
rect 23842 2524 23848 2576
rect 23900 2564 23906 2576
rect 25777 2567 25835 2573
rect 25777 2564 25789 2567
rect 23900 2536 25789 2564
rect 23900 2524 23906 2536
rect 25777 2533 25789 2536
rect 25823 2533 25835 2567
rect 28905 2567 28963 2573
rect 28905 2564 28917 2567
rect 25777 2527 25835 2533
rect 27816 2536 28917 2564
rect 12023 2468 16574 2496
rect 12023 2465 12035 2468
rect 11977 2459 12035 2465
rect 17218 2456 17224 2508
rect 17276 2496 17282 2508
rect 21910 2496 21916 2508
rect 17276 2468 19288 2496
rect 17276 2456 17282 2468
rect 2225 2431 2283 2437
rect 2225 2397 2237 2431
rect 2271 2428 2283 2431
rect 2958 2428 2964 2440
rect 2271 2400 2964 2428
rect 2271 2397 2283 2400
rect 2225 2391 2283 2397
rect 2958 2388 2964 2400
rect 3016 2388 3022 2440
rect 3237 2431 3295 2437
rect 3237 2397 3249 2431
rect 3283 2428 3295 2431
rect 4798 2428 4804 2440
rect 3283 2400 4804 2428
rect 3283 2397 3295 2400
rect 3237 2391 3295 2397
rect 4798 2388 4804 2400
rect 4856 2388 4862 2440
rect 5629 2431 5687 2437
rect 5629 2397 5641 2431
rect 5675 2428 5687 2431
rect 5810 2428 5816 2440
rect 5675 2400 5816 2428
rect 5675 2397 5687 2400
rect 5629 2391 5687 2397
rect 5810 2388 5816 2400
rect 5868 2428 5874 2440
rect 6178 2428 6184 2440
rect 5868 2400 6184 2428
rect 5868 2388 5874 2400
rect 6178 2388 6184 2400
rect 6236 2388 6242 2440
rect 6825 2431 6883 2437
rect 6825 2397 6837 2431
rect 6871 2428 6883 2431
rect 9582 2428 9588 2440
rect 6871 2400 9588 2428
rect 6871 2397 6883 2400
rect 6825 2391 6883 2397
rect 9582 2388 9588 2400
rect 9640 2388 9646 2440
rect 9766 2388 9772 2440
rect 9824 2428 9830 2440
rect 9953 2431 10011 2437
rect 9953 2428 9965 2431
rect 9824 2400 9965 2428
rect 9824 2388 9830 2400
rect 9953 2397 9965 2400
rect 9999 2397 10011 2431
rect 9953 2391 10011 2397
rect 10410 2388 10416 2440
rect 10468 2428 10474 2440
rect 10689 2431 10747 2437
rect 10689 2428 10701 2431
rect 10468 2400 10701 2428
rect 10468 2388 10474 2400
rect 10689 2397 10701 2400
rect 10735 2397 10747 2431
rect 10689 2391 10747 2397
rect 11606 2388 11612 2440
rect 11664 2428 11670 2440
rect 11701 2431 11759 2437
rect 11701 2428 11713 2431
rect 11664 2400 11713 2428
rect 11664 2388 11670 2400
rect 11701 2397 11713 2400
rect 11747 2397 11759 2431
rect 13262 2428 13268 2440
rect 13223 2400 13268 2428
rect 11701 2391 11759 2397
rect 13262 2388 13268 2400
rect 13320 2388 13326 2440
rect 14369 2431 14427 2437
rect 14369 2397 14381 2431
rect 14415 2428 14427 2431
rect 14458 2428 14464 2440
rect 14415 2400 14464 2428
rect 14415 2397 14427 2400
rect 14369 2391 14427 2397
rect 14458 2388 14464 2400
rect 14516 2388 14522 2440
rect 15289 2431 15347 2437
rect 15289 2397 15301 2431
rect 15335 2428 15347 2431
rect 15562 2428 15568 2440
rect 15335 2400 15568 2428
rect 15335 2397 15347 2400
rect 15289 2391 15347 2397
rect 15562 2388 15568 2400
rect 15620 2388 15626 2440
rect 16114 2428 16120 2440
rect 16075 2400 16120 2428
rect 16114 2388 16120 2400
rect 16172 2388 16178 2440
rect 17129 2431 17187 2437
rect 17129 2397 17141 2431
rect 17175 2428 17187 2431
rect 17678 2428 17684 2440
rect 17175 2400 17684 2428
rect 17175 2397 17187 2400
rect 17129 2391 17187 2397
rect 17678 2388 17684 2400
rect 17736 2388 17742 2440
rect 18138 2428 18144 2440
rect 18099 2400 18144 2428
rect 18138 2388 18144 2400
rect 18196 2388 18202 2440
rect 19260 2437 19288 2468
rect 20272 2468 21916 2496
rect 20272 2437 20300 2468
rect 21910 2456 21916 2468
rect 21968 2456 21974 2508
rect 22278 2496 22284 2508
rect 22239 2468 22284 2496
rect 22278 2456 22284 2468
rect 22336 2456 22342 2508
rect 25041 2499 25099 2505
rect 25041 2465 25053 2499
rect 25087 2496 25099 2499
rect 26142 2496 26148 2508
rect 25087 2468 26148 2496
rect 25087 2465 25099 2468
rect 25041 2459 25099 2465
rect 26142 2456 26148 2468
rect 26200 2496 26206 2508
rect 26329 2499 26387 2505
rect 26329 2496 26341 2499
rect 26200 2468 26341 2496
rect 26200 2456 26206 2468
rect 26329 2465 26341 2468
rect 26375 2465 26387 2499
rect 26329 2459 26387 2465
rect 19245 2431 19303 2437
rect 19245 2397 19257 2431
rect 19291 2397 19303 2431
rect 19245 2391 19303 2397
rect 20257 2431 20315 2437
rect 20257 2397 20269 2431
rect 20303 2397 20315 2431
rect 20257 2391 20315 2397
rect 20530 2388 20536 2440
rect 20588 2428 20594 2440
rect 20717 2431 20775 2437
rect 20717 2428 20729 2431
rect 20588 2400 20729 2428
rect 20588 2388 20594 2400
rect 20717 2397 20729 2400
rect 20763 2397 20775 2431
rect 20717 2391 20775 2397
rect 22005 2431 22063 2437
rect 22005 2397 22017 2431
rect 22051 2397 22063 2431
rect 25590 2428 25596 2440
rect 25551 2400 25596 2428
rect 22005 2391 22063 2397
rect 7377 2363 7435 2369
rect 7377 2329 7389 2363
rect 7423 2360 7435 2363
rect 7742 2360 7748 2372
rect 7423 2332 7748 2360
rect 7423 2329 7435 2332
rect 7377 2323 7435 2329
rect 7742 2320 7748 2332
rect 7800 2360 7806 2372
rect 7929 2363 7987 2369
rect 7929 2360 7941 2363
rect 7800 2332 7941 2360
rect 7800 2320 7806 2332
rect 7929 2329 7941 2332
rect 7975 2329 7987 2363
rect 9030 2360 9036 2372
rect 8991 2332 9036 2360
rect 7929 2323 7987 2329
rect 9030 2320 9036 2332
rect 9088 2320 9094 2372
rect 9140 2332 21036 2360
rect 3053 2295 3111 2301
rect 3053 2261 3065 2295
rect 3099 2292 3111 2295
rect 3234 2292 3240 2304
rect 3099 2264 3240 2292
rect 3099 2261 3111 2264
rect 3053 2255 3111 2261
rect 3234 2252 3240 2264
rect 3292 2252 3298 2304
rect 5718 2292 5724 2304
rect 5679 2264 5724 2292
rect 5718 2252 5724 2264
rect 5776 2252 5782 2304
rect 6454 2252 6460 2304
rect 6512 2292 6518 2304
rect 6641 2295 6699 2301
rect 6641 2292 6653 2295
rect 6512 2264 6653 2292
rect 6512 2252 6518 2264
rect 6641 2261 6653 2264
rect 6687 2261 6699 2295
rect 6641 2255 6699 2261
rect 8754 2252 8760 2304
rect 8812 2292 8818 2304
rect 9140 2292 9168 2332
rect 8812 2264 9168 2292
rect 8812 2252 8818 2264
rect 9674 2252 9680 2304
rect 9732 2292 9738 2304
rect 9769 2295 9827 2301
rect 9769 2292 9781 2295
rect 9732 2264 9781 2292
rect 9732 2252 9738 2264
rect 9769 2261 9781 2264
rect 9815 2261 9827 2295
rect 9769 2255 9827 2261
rect 10318 2252 10324 2304
rect 10376 2292 10382 2304
rect 10505 2295 10563 2301
rect 10505 2292 10517 2295
rect 10376 2264 10517 2292
rect 10376 2252 10382 2264
rect 10505 2261 10517 2264
rect 10551 2261 10563 2295
rect 10505 2255 10563 2261
rect 12250 2252 12256 2304
rect 12308 2292 12314 2304
rect 13081 2295 13139 2301
rect 13081 2292 13093 2295
rect 12308 2264 13093 2292
rect 12308 2252 12314 2264
rect 13081 2261 13093 2264
rect 13127 2261 13139 2295
rect 13081 2255 13139 2261
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 14185 2295 14243 2301
rect 14185 2292 14197 2295
rect 13596 2264 14197 2292
rect 13596 2252 13602 2264
rect 14185 2261 14197 2264
rect 14231 2261 14243 2295
rect 14185 2255 14243 2261
rect 16758 2252 16764 2304
rect 16816 2292 16822 2304
rect 16945 2295 17003 2301
rect 16945 2292 16957 2295
rect 16816 2264 16957 2292
rect 16816 2252 16822 2264
rect 16945 2261 16957 2264
rect 16991 2261 17003 2295
rect 16945 2255 17003 2261
rect 18046 2252 18052 2304
rect 18104 2292 18110 2304
rect 18325 2295 18383 2301
rect 18325 2292 18337 2295
rect 18104 2264 18337 2292
rect 18104 2252 18110 2264
rect 18325 2261 18337 2264
rect 18371 2261 18383 2295
rect 18325 2255 18383 2261
rect 19334 2252 19340 2304
rect 19392 2292 19398 2304
rect 19429 2295 19487 2301
rect 19429 2292 19441 2295
rect 19392 2264 19441 2292
rect 19392 2252 19398 2264
rect 19429 2261 19441 2264
rect 19475 2261 19487 2295
rect 19429 2255 19487 2261
rect 19978 2252 19984 2304
rect 20036 2292 20042 2304
rect 20073 2295 20131 2301
rect 20073 2292 20085 2295
rect 20036 2264 20085 2292
rect 20036 2252 20042 2264
rect 20073 2261 20085 2264
rect 20119 2261 20131 2295
rect 20073 2255 20131 2261
rect 20622 2252 20628 2304
rect 20680 2292 20686 2304
rect 20901 2295 20959 2301
rect 20901 2292 20913 2295
rect 20680 2264 20913 2292
rect 20680 2252 20686 2264
rect 20901 2261 20913 2264
rect 20947 2261 20959 2295
rect 21008 2292 21036 2332
rect 21910 2320 21916 2372
rect 21968 2360 21974 2372
rect 22020 2360 22048 2391
rect 25590 2388 25596 2400
rect 25648 2388 25654 2440
rect 27154 2428 27160 2440
rect 27115 2400 27160 2428
rect 27154 2388 27160 2400
rect 27212 2388 27218 2440
rect 27816 2437 27844 2536
rect 28905 2533 28917 2536
rect 28951 2533 28963 2567
rect 28905 2527 28963 2533
rect 29730 2524 29736 2576
rect 29788 2564 29794 2576
rect 36449 2567 36507 2573
rect 36449 2564 36461 2567
rect 29788 2536 36461 2564
rect 29788 2524 29794 2536
rect 36449 2533 36461 2536
rect 36495 2533 36507 2567
rect 36449 2527 36507 2533
rect 27982 2456 27988 2508
rect 28040 2496 28046 2508
rect 32401 2499 32459 2505
rect 32401 2496 32413 2499
rect 28040 2468 32413 2496
rect 28040 2456 28046 2468
rect 32401 2465 32413 2468
rect 32447 2465 32459 2499
rect 32401 2459 32459 2465
rect 35710 2456 35716 2508
rect 35768 2496 35774 2508
rect 37277 2499 37335 2505
rect 37277 2496 37289 2499
rect 35768 2468 37289 2496
rect 35768 2456 35774 2468
rect 37277 2465 37289 2468
rect 37323 2496 37335 2499
rect 37642 2496 37648 2508
rect 37323 2468 37648 2496
rect 37323 2465 37335 2468
rect 37277 2459 37335 2465
rect 37642 2456 37648 2468
rect 37700 2456 37706 2508
rect 27801 2431 27859 2437
rect 27801 2428 27813 2431
rect 27540 2400 27813 2428
rect 21968 2332 22048 2360
rect 23477 2363 23535 2369
rect 21968 2320 21974 2332
rect 23477 2329 23489 2363
rect 23523 2360 23535 2363
rect 23658 2360 23664 2372
rect 23523 2332 23664 2360
rect 23523 2329 23535 2332
rect 23477 2323 23535 2329
rect 23658 2320 23664 2332
rect 23716 2320 23722 2372
rect 24765 2363 24823 2369
rect 24765 2329 24777 2363
rect 24811 2360 24823 2363
rect 24811 2332 25728 2360
rect 24811 2329 24823 2332
rect 24765 2323 24823 2329
rect 23385 2295 23443 2301
rect 23385 2292 23397 2295
rect 21008 2264 23397 2292
rect 20901 2255 20959 2261
rect 23385 2261 23397 2264
rect 23431 2261 23443 2295
rect 24854 2292 24860 2304
rect 24815 2264 24860 2292
rect 23385 2255 23443 2261
rect 24854 2252 24860 2264
rect 24912 2252 24918 2304
rect 25700 2292 25728 2332
rect 25774 2320 25780 2372
rect 25832 2360 25838 2372
rect 27540 2360 27568 2400
rect 27801 2397 27813 2400
rect 27847 2397 27859 2431
rect 27801 2391 27859 2397
rect 28445 2431 28503 2437
rect 28445 2397 28457 2431
rect 28491 2397 28503 2431
rect 28445 2391 28503 2397
rect 25832 2332 27568 2360
rect 25832 2320 25838 2332
rect 27706 2320 27712 2372
rect 27764 2360 27770 2372
rect 28460 2360 28488 2391
rect 29638 2388 29644 2440
rect 29696 2428 29702 2440
rect 29733 2431 29791 2437
rect 29733 2428 29745 2431
rect 29696 2400 29745 2428
rect 29696 2388 29702 2400
rect 29733 2397 29745 2400
rect 29779 2397 29791 2431
rect 30006 2428 30012 2440
rect 29967 2400 30012 2428
rect 29733 2391 29791 2397
rect 30006 2388 30012 2400
rect 30064 2388 30070 2440
rect 30834 2388 30840 2440
rect 30892 2428 30898 2440
rect 31021 2431 31079 2437
rect 31021 2428 31033 2431
rect 30892 2400 31033 2428
rect 30892 2388 30898 2400
rect 31021 2397 31033 2400
rect 31067 2397 31079 2431
rect 31021 2391 31079 2397
rect 31754 2388 31760 2440
rect 31812 2428 31818 2440
rect 32125 2431 32183 2437
rect 32125 2428 32137 2431
rect 31812 2400 32137 2428
rect 31812 2388 31818 2400
rect 32125 2397 32137 2400
rect 32171 2428 32183 2431
rect 32214 2428 32220 2440
rect 32171 2400 32220 2428
rect 32171 2397 32183 2400
rect 32125 2391 32183 2397
rect 32214 2388 32220 2400
rect 32272 2388 32278 2440
rect 33870 2428 33876 2440
rect 33831 2400 33876 2428
rect 33870 2388 33876 2400
rect 33928 2388 33934 2440
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34848 2400 34897 2428
rect 34848 2388 34854 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 36630 2428 36636 2440
rect 36591 2400 36636 2428
rect 34885 2391 34943 2397
rect 36630 2388 36636 2400
rect 36688 2388 36694 2440
rect 37553 2431 37611 2437
rect 37553 2397 37565 2431
rect 37599 2397 37611 2431
rect 37553 2391 37611 2397
rect 27764 2332 28488 2360
rect 35897 2363 35955 2369
rect 27764 2320 27770 2332
rect 35897 2329 35909 2363
rect 35943 2360 35955 2363
rect 36446 2360 36452 2372
rect 35943 2332 36452 2360
rect 35943 2329 35955 2332
rect 35897 2323 35955 2329
rect 36446 2320 36452 2332
rect 36504 2320 36510 2372
rect 28442 2292 28448 2304
rect 25700 2264 28448 2292
rect 28442 2252 28448 2264
rect 28500 2252 28506 2304
rect 30282 2252 30288 2304
rect 30340 2292 30346 2304
rect 31205 2295 31263 2301
rect 31205 2292 31217 2295
rect 30340 2264 31217 2292
rect 30340 2252 30346 2264
rect 31205 2261 31217 2264
rect 31251 2261 31263 2295
rect 31205 2255 31263 2261
rect 33502 2252 33508 2304
rect 33560 2292 33566 2304
rect 33689 2295 33747 2301
rect 33689 2292 33701 2295
rect 33560 2264 33701 2292
rect 33560 2252 33566 2264
rect 33689 2261 33701 2264
rect 33735 2261 33747 2295
rect 33689 2255 33747 2261
rect 34790 2252 34796 2304
rect 34848 2292 34854 2304
rect 35069 2295 35127 2301
rect 35069 2292 35081 2295
rect 34848 2264 35081 2292
rect 34848 2252 34854 2264
rect 35069 2261 35081 2264
rect 35115 2261 35127 2295
rect 35069 2255 35127 2261
rect 35158 2252 35164 2304
rect 35216 2292 35222 2304
rect 37568 2292 37596 2391
rect 35216 2264 37596 2292
rect 35216 2252 35222 2264
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
rect 20070 2048 20076 2100
rect 20128 2088 20134 2100
rect 30006 2088 30012 2100
rect 20128 2060 30012 2088
rect 20128 2048 20134 2060
rect 30006 2048 30012 2060
rect 30064 2048 30070 2100
rect 5718 1980 5724 2032
rect 5776 2020 5782 2032
rect 24302 2020 24308 2032
rect 5776 1992 24308 2020
rect 5776 1980 5782 1992
rect 24302 1980 24308 1992
rect 24360 1980 24366 2032
rect 29914 1980 29920 2032
rect 29972 2020 29978 2032
rect 35158 2020 35164 2032
rect 29972 1992 35164 2020
rect 29972 1980 29978 1992
rect 35158 1980 35164 1992
rect 35216 1980 35222 2032
rect 24854 1912 24860 1964
rect 24912 1952 24918 1964
rect 31478 1952 31484 1964
rect 24912 1924 31484 1952
rect 24912 1912 24918 1924
rect 31478 1912 31484 1924
rect 31536 1912 31542 1964
rect 25130 1844 25136 1896
rect 25188 1884 25194 1896
rect 27154 1884 27160 1896
rect 25188 1856 27160 1884
rect 25188 1844 25194 1856
rect 27154 1844 27160 1856
rect 27212 1844 27218 1896
rect 22554 1708 22560 1760
rect 22612 1748 22618 1760
rect 23658 1748 23664 1760
rect 22612 1720 23664 1748
rect 22612 1708 22618 1720
rect 23658 1708 23664 1720
rect 23716 1708 23722 1760
<< via1 >>
rect 13820 47472 13872 47524
rect 20076 47472 20128 47524
rect 20 47404 72 47456
rect 940 47404 992 47456
rect 10968 47404 11020 47456
rect 24308 47404 24360 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 4620 47243 4672 47252
rect 4620 47209 4629 47243
rect 4629 47209 4663 47243
rect 4663 47209 4672 47243
rect 4620 47200 4672 47209
rect 9864 47243 9916 47252
rect 6460 47132 6512 47184
rect 9864 47209 9873 47243
rect 9873 47209 9907 47243
rect 9907 47209 9916 47243
rect 9864 47200 9916 47209
rect 10968 47243 11020 47252
rect 10968 47209 10977 47243
rect 10977 47209 11011 47243
rect 11011 47209 11020 47243
rect 10968 47200 11020 47209
rect 14464 47200 14516 47252
rect 16764 47200 16816 47252
rect 17960 47200 18012 47252
rect 20076 47243 20128 47252
rect 20076 47209 20085 47243
rect 20085 47209 20119 47243
rect 20119 47209 20128 47243
rect 20076 47200 20128 47209
rect 20720 47200 20772 47252
rect 22468 47243 22520 47252
rect 22468 47209 22477 47243
rect 22477 47209 22511 47243
rect 22511 47209 22520 47243
rect 22468 47200 22520 47209
rect 26424 47200 26476 47252
rect 27344 47200 27396 47252
rect 30380 47200 30432 47252
rect 30932 47200 30984 47252
rect 31760 47200 31812 47252
rect 36636 47243 36688 47252
rect 36636 47209 36645 47243
rect 36645 47209 36679 47243
rect 36679 47209 36688 47243
rect 36636 47200 36688 47209
rect 7196 47107 7248 47116
rect 2044 47039 2096 47048
rect 2044 47005 2053 47039
rect 2053 47005 2087 47039
rect 2087 47005 2096 47039
rect 2044 46996 2096 47005
rect 2596 46996 2648 47048
rect 3240 46996 3292 47048
rect 4804 47039 4856 47048
rect 2688 46860 2740 46912
rect 3792 46860 3844 46912
rect 3976 46928 4028 46980
rect 4804 47005 4813 47039
rect 4813 47005 4847 47039
rect 4847 47005 4856 47039
rect 4804 46996 4856 47005
rect 5356 47039 5408 47048
rect 5356 47005 5365 47039
rect 5365 47005 5399 47039
rect 5399 47005 5408 47039
rect 5356 46996 5408 47005
rect 6552 47039 6604 47048
rect 6552 47005 6561 47039
rect 6561 47005 6595 47039
rect 6595 47005 6604 47039
rect 6552 46996 6604 47005
rect 7196 47073 7205 47107
rect 7205 47073 7239 47107
rect 7239 47073 7248 47107
rect 7196 47064 7248 47073
rect 7472 47039 7524 47048
rect 7472 47005 7481 47039
rect 7481 47005 7515 47039
rect 7515 47005 7524 47039
rect 7472 46996 7524 47005
rect 8392 46996 8444 47048
rect 8944 46996 8996 47048
rect 10048 47039 10100 47048
rect 10048 47005 10057 47039
rect 10057 47005 10091 47039
rect 10091 47005 10100 47039
rect 10048 46996 10100 47005
rect 10784 47039 10836 47048
rect 10784 47005 10793 47039
rect 10793 47005 10827 47039
rect 10827 47005 10836 47039
rect 10784 46996 10836 47005
rect 11980 47039 12032 47048
rect 11980 47005 11989 47039
rect 11989 47005 12023 47039
rect 12023 47005 12032 47039
rect 11980 46996 12032 47005
rect 12440 46996 12492 47048
rect 12624 47039 12676 47048
rect 12624 47005 12633 47039
rect 12633 47005 12667 47039
rect 12667 47005 12676 47039
rect 12624 46996 12676 47005
rect 5540 46971 5592 46980
rect 5540 46937 5549 46971
rect 5549 46937 5583 46971
rect 5583 46937 5592 46971
rect 5540 46928 5592 46937
rect 9220 46928 9272 46980
rect 13268 47039 13320 47048
rect 13268 47005 13277 47039
rect 13277 47005 13311 47039
rect 13311 47005 13320 47039
rect 13268 46996 13320 47005
rect 13912 47064 13964 47116
rect 14280 47107 14332 47116
rect 14280 47073 14289 47107
rect 14289 47073 14323 47107
rect 14323 47073 14332 47107
rect 14280 47064 14332 47073
rect 15384 47064 15436 47116
rect 18052 47132 18104 47184
rect 14648 46996 14700 47048
rect 16672 47039 16724 47048
rect 16672 47005 16681 47039
rect 16681 47005 16715 47039
rect 16715 47005 16724 47039
rect 16672 46996 16724 47005
rect 16948 47039 17000 47048
rect 16948 47005 16957 47039
rect 16957 47005 16991 47039
rect 16991 47005 17000 47039
rect 16948 46996 17000 47005
rect 17408 46928 17460 46980
rect 20444 47064 20496 47116
rect 17960 47039 18012 47048
rect 17960 47005 17969 47039
rect 17969 47005 18003 47039
rect 18003 47005 18012 47039
rect 17960 46996 18012 47005
rect 19340 46996 19392 47048
rect 19616 47039 19668 47048
rect 19616 47005 19625 47039
rect 19625 47005 19659 47039
rect 19659 47005 19668 47039
rect 19616 46996 19668 47005
rect 20260 47039 20312 47048
rect 20260 47005 20269 47039
rect 20269 47005 20303 47039
rect 20303 47005 20312 47039
rect 20260 46996 20312 47005
rect 26148 47132 26200 47184
rect 27712 47132 27764 47184
rect 34796 47132 34848 47184
rect 23020 47107 23072 47116
rect 23020 47073 23029 47107
rect 23029 47073 23063 47107
rect 23063 47073 23072 47107
rect 23020 47064 23072 47073
rect 23848 47064 23900 47116
rect 24400 47107 24452 47116
rect 24400 47073 24409 47107
rect 24409 47073 24443 47107
rect 24443 47073 24452 47107
rect 24400 47064 24452 47073
rect 24860 47064 24912 47116
rect 32956 47107 33008 47116
rect 21088 46996 21140 47048
rect 22836 46996 22888 47048
rect 23296 47039 23348 47048
rect 23296 47005 23305 47039
rect 23305 47005 23339 47039
rect 23339 47005 23348 47039
rect 23296 46996 23348 47005
rect 24676 47039 24728 47048
rect 24676 47005 24685 47039
rect 24685 47005 24719 47039
rect 24719 47005 24728 47039
rect 24676 46996 24728 47005
rect 26056 47039 26108 47048
rect 26056 47005 26065 47039
rect 26065 47005 26099 47039
rect 26099 47005 26108 47039
rect 26056 46996 26108 47005
rect 26976 47039 27028 47048
rect 26976 47005 26985 47039
rect 26985 47005 27019 47039
rect 27019 47005 27028 47039
rect 26976 46996 27028 47005
rect 27344 46996 27396 47048
rect 27896 46996 27948 47048
rect 29000 46996 29052 47048
rect 29644 46996 29696 47048
rect 25412 46928 25464 46980
rect 27436 46928 27488 46980
rect 30932 46996 30984 47048
rect 31484 46996 31536 47048
rect 32956 47073 32965 47107
rect 32965 47073 32999 47107
rect 32999 47073 33008 47107
rect 32956 47064 33008 47073
rect 35624 47064 35676 47116
rect 34520 46996 34572 47048
rect 36084 46996 36136 47048
rect 16120 46860 16172 46912
rect 16672 46860 16724 46912
rect 29552 46903 29604 46912
rect 29552 46869 29561 46903
rect 29561 46869 29595 46903
rect 29595 46869 29604 46903
rect 29552 46860 29604 46869
rect 36360 46860 36412 46912
rect 37280 46860 37332 46912
rect 37648 46860 37700 46912
rect 39304 46860 39356 46912
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 664 46656 716 46708
rect 3884 46656 3936 46708
rect 5356 46656 5408 46708
rect 5816 46699 5868 46708
rect 5816 46665 5825 46699
rect 5825 46665 5859 46699
rect 5859 46665 5868 46699
rect 5816 46656 5868 46665
rect 7196 46656 7248 46708
rect 7932 46699 7984 46708
rect 7932 46665 7941 46699
rect 7941 46665 7975 46699
rect 7975 46665 7984 46699
rect 7932 46656 7984 46665
rect 10784 46656 10836 46708
rect 13820 46699 13872 46708
rect 13820 46665 13829 46699
rect 13829 46665 13863 46699
rect 13863 46665 13872 46699
rect 13820 46656 13872 46665
rect 15476 46656 15528 46708
rect 17408 46699 17460 46708
rect 17408 46665 17417 46699
rect 17417 46665 17451 46699
rect 17451 46665 17460 46699
rect 17408 46656 17460 46665
rect 20260 46656 20312 46708
rect 21272 46699 21324 46708
rect 21272 46665 21281 46699
rect 21281 46665 21315 46699
rect 21315 46665 21324 46699
rect 21272 46656 21324 46665
rect 23020 46656 23072 46708
rect 26056 46656 26108 46708
rect 35440 46656 35492 46708
rect 37372 46656 37424 46708
rect 37464 46656 37516 46708
rect 3056 46588 3108 46640
rect 3148 46520 3200 46572
rect 14372 46588 14424 46640
rect 8300 46520 8352 46572
rect 9128 46563 9180 46572
rect 9128 46529 9137 46563
rect 9137 46529 9171 46563
rect 9171 46529 9180 46563
rect 9128 46520 9180 46529
rect 11704 46563 11756 46572
rect 11704 46529 11713 46563
rect 11713 46529 11747 46563
rect 11747 46529 11756 46563
rect 11704 46520 11756 46529
rect 13728 46563 13780 46572
rect 13728 46529 13737 46563
rect 13737 46529 13771 46563
rect 13771 46529 13780 46563
rect 13728 46520 13780 46529
rect 8392 46452 8444 46504
rect 15292 46452 15344 46504
rect 2504 46384 2556 46436
rect 16212 46520 16264 46572
rect 18788 46563 18840 46572
rect 16488 46452 16540 46504
rect 18788 46529 18797 46563
rect 18797 46529 18831 46563
rect 18831 46529 18840 46563
rect 18788 46520 18840 46529
rect 32220 46588 32272 46640
rect 21916 46520 21968 46572
rect 24768 46563 24820 46572
rect 24768 46529 24777 46563
rect 24777 46529 24811 46563
rect 24811 46529 24820 46563
rect 24768 46520 24820 46529
rect 28632 46563 28684 46572
rect 28632 46529 28641 46563
rect 28641 46529 28675 46563
rect 28675 46529 28684 46563
rect 28632 46520 28684 46529
rect 29920 46563 29972 46572
rect 29920 46529 29929 46563
rect 29929 46529 29963 46563
rect 29963 46529 29972 46563
rect 29920 46520 29972 46529
rect 33784 46563 33836 46572
rect 33784 46529 33793 46563
rect 33793 46529 33827 46563
rect 33827 46529 33836 46563
rect 33784 46520 33836 46529
rect 34428 46563 34480 46572
rect 34428 46529 34437 46563
rect 34437 46529 34471 46563
rect 34471 46529 34480 46563
rect 34428 46520 34480 46529
rect 34796 46520 34848 46572
rect 35900 46563 35952 46572
rect 35900 46529 35909 46563
rect 35909 46529 35943 46563
rect 35943 46529 35952 46563
rect 35900 46520 35952 46529
rect 36268 46520 36320 46572
rect 29552 46452 29604 46504
rect 35532 46452 35584 46504
rect 37464 46452 37516 46504
rect 2320 46316 2372 46368
rect 3056 46359 3108 46368
rect 3056 46325 3065 46359
rect 3065 46325 3099 46359
rect 3099 46325 3108 46359
rect 3056 46316 3108 46325
rect 5356 46316 5408 46368
rect 6552 46359 6604 46368
rect 6552 46325 6561 46359
rect 6561 46325 6595 46359
rect 6595 46325 6604 46359
rect 6552 46316 6604 46325
rect 10048 46316 10100 46368
rect 10692 46316 10744 46368
rect 12716 46316 12768 46368
rect 13452 46316 13504 46368
rect 14280 46316 14332 46368
rect 27160 46384 27212 46436
rect 31576 46384 31628 46436
rect 35440 46384 35492 46436
rect 15200 46316 15252 46368
rect 17776 46316 17828 46368
rect 18972 46359 19024 46368
rect 18972 46325 18981 46359
rect 18981 46325 19015 46359
rect 19015 46325 19024 46359
rect 18972 46316 19024 46325
rect 22100 46316 22152 46368
rect 22192 46316 22244 46368
rect 27896 46359 27948 46368
rect 27896 46325 27905 46359
rect 27905 46325 27939 46359
rect 27939 46325 27948 46359
rect 27896 46316 27948 46325
rect 28448 46359 28500 46368
rect 28448 46325 28457 46359
rect 28457 46325 28491 46359
rect 28491 46325 28500 46359
rect 28448 46316 28500 46325
rect 30932 46359 30984 46368
rect 30932 46325 30941 46359
rect 30941 46325 30975 46359
rect 30975 46325 30984 46359
rect 30932 46316 30984 46325
rect 31484 46359 31536 46368
rect 31484 46325 31493 46359
rect 31493 46325 31527 46359
rect 31527 46325 31536 46359
rect 31484 46316 31536 46325
rect 32588 46359 32640 46368
rect 32588 46325 32597 46359
rect 32597 46325 32631 46359
rect 32631 46325 32640 46359
rect 32588 46316 32640 46325
rect 33600 46359 33652 46368
rect 33600 46325 33609 46359
rect 33609 46325 33643 46359
rect 33643 46325 33652 46359
rect 33600 46316 33652 46325
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 2780 46112 2832 46164
rect 2964 46155 3016 46164
rect 2964 46121 2973 46155
rect 2973 46121 3007 46155
rect 3007 46121 3016 46155
rect 2964 46112 3016 46121
rect 3884 46112 3936 46164
rect 4804 46112 4856 46164
rect 5080 46112 5132 46164
rect 6644 46112 6696 46164
rect 8944 46155 8996 46164
rect 8944 46121 8953 46155
rect 8953 46121 8987 46155
rect 8987 46121 8996 46155
rect 8944 46112 8996 46121
rect 11704 46112 11756 46164
rect 11980 46112 12032 46164
rect 12716 46112 12768 46164
rect 15108 46155 15160 46164
rect 3240 46044 3292 46096
rect 15108 46121 15117 46155
rect 15117 46121 15151 46155
rect 15151 46121 15160 46155
rect 15108 46112 15160 46121
rect 15200 46112 15252 46164
rect 17132 46112 17184 46164
rect 19340 46155 19392 46164
rect 19340 46121 19349 46155
rect 19349 46121 19383 46155
rect 19383 46121 19392 46155
rect 19340 46112 19392 46121
rect 24400 46155 24452 46164
rect 24400 46121 24409 46155
rect 24409 46121 24443 46155
rect 24443 46121 24452 46155
rect 24400 46112 24452 46121
rect 29644 46155 29696 46164
rect 29644 46121 29653 46155
rect 29653 46121 29687 46155
rect 29687 46121 29696 46155
rect 29644 46112 29696 46121
rect 32220 46112 32272 46164
rect 32956 46155 33008 46164
rect 32956 46121 32965 46155
rect 32965 46121 32999 46155
rect 32999 46121 33008 46155
rect 32956 46112 33008 46121
rect 33784 46112 33836 46164
rect 34428 46112 34480 46164
rect 35808 46112 35860 46164
rect 2320 45908 2372 45960
rect 2688 45908 2740 45960
rect 3240 45908 3292 45960
rect 13268 45908 13320 45960
rect 13452 45951 13504 45960
rect 13452 45917 13461 45951
rect 13461 45917 13495 45951
rect 13495 45917 13504 45951
rect 13452 45908 13504 45917
rect 14280 45951 14332 45960
rect 14280 45917 14289 45951
rect 14289 45917 14323 45951
rect 14323 45917 14332 45951
rect 14280 45908 14332 45917
rect 20812 46044 20864 46096
rect 23480 46044 23532 46096
rect 33600 46044 33652 46096
rect 35716 46044 35768 46096
rect 16028 45976 16080 46028
rect 16488 45976 16540 46028
rect 18052 45976 18104 46028
rect 35256 45976 35308 46028
rect 35532 45976 35584 46028
rect 37648 45976 37700 46028
rect 15384 45908 15436 45960
rect 18328 45951 18380 45960
rect 18328 45917 18337 45951
rect 18337 45917 18371 45951
rect 18371 45917 18380 45951
rect 18328 45908 18380 45917
rect 35348 45951 35400 45960
rect 35348 45917 35357 45951
rect 35357 45917 35391 45951
rect 35391 45917 35400 45951
rect 35348 45908 35400 45917
rect 8300 45883 8352 45892
rect 8300 45849 8309 45883
rect 8309 45849 8343 45883
rect 8343 45849 8352 45883
rect 8300 45840 8352 45849
rect 9036 45840 9088 45892
rect 34612 45840 34664 45892
rect 35992 45908 36044 45960
rect 37556 45951 37608 45960
rect 37556 45917 37565 45951
rect 37565 45917 37599 45951
rect 37599 45917 37608 45951
rect 37556 45908 37608 45917
rect 1492 45815 1544 45824
rect 1492 45781 1501 45815
rect 1501 45781 1535 45815
rect 1535 45781 1544 45815
rect 1492 45772 1544 45781
rect 2964 45772 3016 45824
rect 3148 45772 3200 45824
rect 16028 45815 16080 45824
rect 16028 45781 16037 45815
rect 16037 45781 16071 45815
rect 16071 45781 16080 45815
rect 16028 45772 16080 45781
rect 17316 45815 17368 45824
rect 17316 45781 17325 45815
rect 17325 45781 17359 45815
rect 17359 45781 17368 45815
rect 17316 45772 17368 45781
rect 17868 45772 17920 45824
rect 35624 45772 35676 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 18788 45568 18840 45620
rect 35348 45568 35400 45620
rect 20 45500 72 45552
rect 112 45432 164 45484
rect 1308 45432 1360 45484
rect 2964 45500 3016 45552
rect 12624 45500 12676 45552
rect 13912 45543 13964 45552
rect 13912 45509 13921 45543
rect 13921 45509 13955 45543
rect 13955 45509 13964 45543
rect 13912 45500 13964 45509
rect 17316 45500 17368 45552
rect 34704 45500 34756 45552
rect 37372 45543 37424 45552
rect 2596 45432 2648 45484
rect 17776 45475 17828 45484
rect 17776 45441 17785 45475
rect 17785 45441 17819 45475
rect 17819 45441 17828 45475
rect 17776 45432 17828 45441
rect 35256 45432 35308 45484
rect 37372 45509 37381 45543
rect 37381 45509 37415 45543
rect 37415 45509 37424 45543
rect 37372 45500 37424 45509
rect 36820 45432 36872 45484
rect 2412 45296 2464 45348
rect 13728 45296 13780 45348
rect 17592 45296 17644 45348
rect 17960 45339 18012 45348
rect 17960 45305 17969 45339
rect 17969 45305 18003 45339
rect 18003 45305 18012 45339
rect 17960 45296 18012 45305
rect 22008 45296 22060 45348
rect 35992 45339 36044 45348
rect 35992 45305 36001 45339
rect 36001 45305 36035 45339
rect 36035 45305 36044 45339
rect 35992 45296 36044 45305
rect 3240 45271 3292 45280
rect 3240 45237 3249 45271
rect 3249 45237 3283 45271
rect 3283 45237 3292 45271
rect 3240 45228 3292 45237
rect 14372 45271 14424 45280
rect 14372 45237 14381 45271
rect 14381 45237 14415 45271
rect 14415 45237 14424 45271
rect 14372 45228 14424 45237
rect 15200 45228 15252 45280
rect 16028 45271 16080 45280
rect 16028 45237 16037 45271
rect 16037 45237 16071 45271
rect 16071 45237 16080 45271
rect 16028 45228 16080 45237
rect 34796 45271 34848 45280
rect 34796 45237 34805 45271
rect 34805 45237 34839 45271
rect 34839 45237 34848 45271
rect 34796 45228 34848 45237
rect 36544 45271 36596 45280
rect 36544 45237 36553 45271
rect 36553 45237 36587 45271
rect 36587 45237 36596 45271
rect 36544 45228 36596 45237
rect 38016 45271 38068 45280
rect 38016 45237 38025 45271
rect 38025 45237 38059 45271
rect 38059 45237 38068 45271
rect 38016 45228 38068 45237
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 3792 45067 3844 45076
rect 3792 45033 3801 45067
rect 3801 45033 3835 45067
rect 3835 45033 3844 45067
rect 3792 45024 3844 45033
rect 16672 45067 16724 45076
rect 16672 45033 16681 45067
rect 16681 45033 16715 45067
rect 16715 45033 16724 45067
rect 16672 45024 16724 45033
rect 18328 45024 18380 45076
rect 35900 45024 35952 45076
rect 30380 44956 30432 45008
rect 33600 44931 33652 44940
rect 33600 44897 33609 44931
rect 33609 44897 33643 44931
rect 33643 44897 33652 44931
rect 33600 44888 33652 44897
rect 2780 44820 2832 44872
rect 36544 44820 36596 44872
rect 37188 44820 37240 44872
rect 38108 44888 38160 44940
rect 2872 44752 2924 44804
rect 7472 44752 7524 44804
rect 37648 44752 37700 44804
rect 1952 44727 2004 44736
rect 1952 44693 1961 44727
rect 1961 44693 1995 44727
rect 1995 44693 2004 44727
rect 1952 44684 2004 44693
rect 4620 44684 4672 44736
rect 16212 44727 16264 44736
rect 16212 44693 16221 44727
rect 16221 44693 16255 44727
rect 16255 44693 16264 44727
rect 16212 44684 16264 44693
rect 34704 44684 34756 44736
rect 38200 44684 38252 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 2872 44480 2924 44532
rect 1308 44412 1360 44464
rect 1400 44387 1452 44396
rect 1400 44353 1409 44387
rect 1409 44353 1443 44387
rect 1443 44353 1452 44387
rect 1400 44344 1452 44353
rect 1768 44140 1820 44192
rect 22100 44251 22152 44260
rect 22100 44217 22109 44251
rect 22109 44217 22143 44251
rect 22143 44217 22152 44251
rect 22100 44208 22152 44217
rect 38016 44251 38068 44260
rect 38016 44217 38025 44251
rect 38025 44217 38059 44251
rect 38059 44217 38068 44251
rect 38016 44208 38068 44217
rect 22468 44140 22520 44192
rect 33600 44140 33652 44192
rect 35532 44140 35584 44192
rect 36084 44140 36136 44192
rect 36268 44183 36320 44192
rect 36268 44149 36277 44183
rect 36277 44149 36311 44183
rect 36311 44149 36320 44183
rect 36268 44140 36320 44149
rect 37280 44183 37332 44192
rect 37280 44149 37289 44183
rect 37289 44149 37323 44183
rect 37323 44149 37332 44183
rect 37280 44140 37332 44149
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 22468 43979 22520 43988
rect 22468 43945 22477 43979
rect 22477 43945 22511 43979
rect 22511 43945 22520 43979
rect 22468 43936 22520 43945
rect 37372 43936 37424 43988
rect 1400 43775 1452 43784
rect 1400 43741 1409 43775
rect 1409 43741 1443 43775
rect 1443 43741 1452 43775
rect 1400 43732 1452 43741
rect 34704 43775 34756 43784
rect 34704 43741 34713 43775
rect 34713 43741 34747 43775
rect 34747 43741 34756 43775
rect 34704 43732 34756 43741
rect 37280 43775 37332 43784
rect 37280 43741 37289 43775
rect 37289 43741 37323 43775
rect 37323 43741 37332 43775
rect 37280 43732 37332 43741
rect 23756 43664 23808 43716
rect 2596 43596 2648 43648
rect 27988 43596 28040 43648
rect 35348 43596 35400 43648
rect 36728 43639 36780 43648
rect 36728 43605 36737 43639
rect 36737 43605 36771 43639
rect 36771 43605 36780 43639
rect 36728 43596 36780 43605
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 26148 43392 26200 43444
rect 31576 43392 31628 43444
rect 1400 43299 1452 43308
rect 1400 43265 1409 43299
rect 1409 43265 1443 43299
rect 1443 43265 1452 43299
rect 1400 43256 1452 43265
rect 35532 43324 35584 43376
rect 26424 43299 26476 43308
rect 26424 43265 26433 43299
rect 26433 43265 26467 43299
rect 26467 43265 26476 43299
rect 26424 43256 26476 43265
rect 30380 43256 30432 43308
rect 38016 43299 38068 43308
rect 38016 43265 38025 43299
rect 38025 43265 38059 43299
rect 38059 43265 38068 43299
rect 38016 43256 38068 43265
rect 4896 43231 4948 43240
rect 4896 43197 4905 43231
rect 4905 43197 4939 43231
rect 4939 43197 4948 43231
rect 4896 43188 4948 43197
rect 27988 43188 28040 43240
rect 4988 43120 5040 43172
rect 37648 43120 37700 43172
rect 27068 43095 27120 43104
rect 27068 43061 27077 43095
rect 27077 43061 27111 43095
rect 27111 43061 27120 43095
rect 27068 43052 27120 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 4896 42848 4948 42900
rect 4988 42848 5040 42900
rect 20628 42848 20680 42900
rect 26424 42848 26476 42900
rect 1400 42687 1452 42696
rect 1400 42653 1409 42687
rect 1409 42653 1443 42687
rect 1443 42653 1452 42687
rect 1400 42644 1452 42653
rect 4620 42712 4672 42764
rect 12440 42712 12492 42764
rect 18512 42712 18564 42764
rect 27988 42755 28040 42764
rect 27988 42721 27997 42755
rect 27997 42721 28031 42755
rect 28031 42721 28040 42755
rect 27988 42712 28040 42721
rect 4712 42644 4764 42696
rect 27068 42644 27120 42696
rect 37372 42644 37424 42696
rect 38108 42687 38160 42696
rect 38108 42653 38117 42687
rect 38117 42653 38151 42687
rect 38151 42653 38160 42687
rect 38108 42644 38160 42653
rect 3700 42576 3752 42628
rect 9496 42576 9548 42628
rect 35624 42576 35676 42628
rect 4712 42508 4764 42560
rect 26608 42508 26660 42560
rect 37832 42508 37884 42560
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 20628 42304 20680 42356
rect 27344 42347 27396 42356
rect 27344 42313 27353 42347
rect 27353 42313 27387 42347
rect 27387 42313 27396 42347
rect 27344 42304 27396 42313
rect 27160 42211 27212 42220
rect 27160 42177 27169 42211
rect 27169 42177 27203 42211
rect 27203 42177 27212 42211
rect 27160 42168 27212 42177
rect 1860 41964 1912 42016
rect 3700 41964 3752 42016
rect 26148 41964 26200 42016
rect 27988 41964 28040 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 26976 41760 27028 41812
rect 37372 41760 37424 41812
rect 21640 41624 21692 41676
rect 1860 41599 1912 41608
rect 1860 41565 1869 41599
rect 1869 41565 1903 41599
rect 1903 41565 1912 41599
rect 1860 41556 1912 41565
rect 20628 41556 20680 41608
rect 4068 41488 4120 41540
rect 21732 41420 21784 41472
rect 38108 41599 38160 41608
rect 38108 41565 38117 41599
rect 38117 41565 38151 41599
rect 38151 41565 38160 41599
rect 38108 41556 38160 41565
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 27160 41216 27212 41268
rect 27344 41080 27396 41132
rect 35716 41216 35768 41268
rect 2228 41055 2280 41064
rect 2228 41021 2237 41055
rect 2237 41021 2271 41055
rect 2271 41021 2280 41055
rect 2228 41012 2280 41021
rect 21640 41012 21692 41064
rect 19248 40944 19300 40996
rect 38108 41123 38160 41132
rect 38108 41089 38117 41123
rect 38117 41089 38151 41123
rect 38151 41089 38160 41123
rect 38108 41080 38160 41089
rect 20904 40919 20956 40928
rect 20904 40885 20913 40919
rect 20913 40885 20947 40919
rect 20947 40885 20956 40919
rect 20904 40876 20956 40885
rect 21732 40876 21784 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 38108 40511 38160 40520
rect 38108 40477 38117 40511
rect 38117 40477 38151 40511
rect 38151 40477 38160 40511
rect 38108 40468 38160 40477
rect 1860 40443 1912 40452
rect 1860 40409 1869 40443
rect 1869 40409 1903 40443
rect 1903 40409 1912 40443
rect 1860 40400 1912 40409
rect 2044 40443 2096 40452
rect 2044 40409 2053 40443
rect 2053 40409 2087 40443
rect 2087 40409 2096 40443
rect 2044 40400 2096 40409
rect 22744 40400 22796 40452
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 38292 39992 38344 40044
rect 1400 39967 1452 39976
rect 1400 39933 1409 39967
rect 1409 39933 1443 39967
rect 1443 39933 1452 39967
rect 1400 39924 1452 39933
rect 1584 39924 1636 39976
rect 38016 39831 38068 39840
rect 38016 39797 38025 39831
rect 38025 39797 38059 39831
rect 38059 39797 38068 39831
rect 38016 39788 38068 39797
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 21916 39584 21968 39636
rect 24860 39584 24912 39636
rect 1400 39559 1452 39568
rect 1400 39525 1409 39559
rect 1409 39525 1443 39559
rect 1443 39525 1452 39559
rect 1400 39516 1452 39525
rect 20812 39448 20864 39500
rect 21916 39448 21968 39500
rect 2688 39380 2740 39432
rect 10324 39380 10376 39432
rect 19432 39380 19484 39432
rect 20628 39423 20680 39432
rect 20628 39389 20637 39423
rect 20637 39389 20671 39423
rect 20671 39389 20680 39423
rect 20628 39380 20680 39389
rect 22008 39380 22060 39432
rect 1952 39312 2004 39364
rect 12256 39312 12308 39364
rect 20996 39312 21048 39364
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 20628 39040 20680 39092
rect 15476 38904 15528 38956
rect 19432 38904 19484 38956
rect 21272 38904 21324 38956
rect 20812 38836 20864 38888
rect 1492 38811 1544 38820
rect 1492 38777 1501 38811
rect 1501 38777 1535 38811
rect 1535 38777 1544 38811
rect 1492 38768 1544 38777
rect 27620 38700 27672 38752
rect 38016 38811 38068 38820
rect 38016 38777 38025 38811
rect 38025 38777 38059 38811
rect 38059 38777 38068 38811
rect 38016 38768 38068 38777
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 20996 38496 21048 38548
rect 21916 38539 21968 38548
rect 21916 38505 21925 38539
rect 21925 38505 21959 38539
rect 21959 38505 21968 38539
rect 21916 38496 21968 38505
rect 2228 38335 2280 38344
rect 2228 38301 2237 38335
rect 2237 38301 2271 38335
rect 2271 38301 2280 38335
rect 2228 38292 2280 38301
rect 14464 38292 14516 38344
rect 15016 38292 15068 38344
rect 21272 38335 21324 38344
rect 21272 38301 21281 38335
rect 21281 38301 21315 38335
rect 21315 38301 21324 38335
rect 21272 38292 21324 38301
rect 38108 38335 38160 38344
rect 38108 38301 38117 38335
rect 38117 38301 38151 38335
rect 38151 38301 38160 38335
rect 38108 38292 38160 38301
rect 20996 38224 21048 38276
rect 37740 38156 37792 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 8392 37995 8444 38004
rect 8392 37961 8401 37995
rect 8401 37961 8435 37995
rect 8435 37961 8444 37995
rect 8392 37952 8444 37961
rect 15476 37952 15528 38004
rect 22284 37952 22336 38004
rect 4068 37884 4120 37936
rect 24952 37884 25004 37936
rect 8576 37859 8628 37868
rect 8576 37825 8585 37859
rect 8585 37825 8619 37859
rect 8619 37825 8628 37859
rect 8576 37816 8628 37825
rect 35348 37816 35400 37868
rect 2228 37791 2280 37800
rect 2228 37757 2237 37791
rect 2237 37757 2271 37791
rect 2271 37757 2280 37791
rect 2228 37748 2280 37757
rect 22560 37680 22612 37732
rect 38016 37655 38068 37664
rect 38016 37621 38025 37655
rect 38025 37621 38059 37655
rect 38059 37621 38068 37655
rect 38016 37612 38068 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 8576 37408 8628 37460
rect 22744 37451 22796 37460
rect 22744 37417 22753 37451
rect 22753 37417 22787 37451
rect 22787 37417 22796 37451
rect 22744 37408 22796 37417
rect 9956 37272 10008 37324
rect 9496 37247 9548 37256
rect 9496 37213 9505 37247
rect 9505 37213 9539 37247
rect 9539 37213 9548 37247
rect 9496 37204 9548 37213
rect 22100 37204 22152 37256
rect 38108 37247 38160 37256
rect 38108 37213 38117 37247
rect 38117 37213 38151 37247
rect 38151 37213 38160 37247
rect 38108 37204 38160 37213
rect 1492 37111 1544 37120
rect 1492 37077 1501 37111
rect 1501 37077 1535 37111
rect 1535 37077 1544 37111
rect 1492 37068 1544 37077
rect 2136 37111 2188 37120
rect 2136 37077 2145 37111
rect 2145 37077 2179 37111
rect 2179 37077 2188 37111
rect 2136 37068 2188 37077
rect 31484 37068 31536 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 22192 36907 22244 36916
rect 22192 36873 22201 36907
rect 22201 36873 22235 36907
rect 22235 36873 22244 36907
rect 22192 36864 22244 36873
rect 22744 36864 22796 36916
rect 23480 36907 23532 36916
rect 23480 36873 23489 36907
rect 23489 36873 23523 36907
rect 23523 36873 23532 36907
rect 23480 36864 23532 36873
rect 38108 36839 38160 36848
rect 38108 36805 38117 36839
rect 38117 36805 38151 36839
rect 38151 36805 38160 36839
rect 38108 36796 38160 36805
rect 9956 36567 10008 36576
rect 9956 36533 9965 36567
rect 9965 36533 9999 36567
rect 9999 36533 10008 36567
rect 21732 36660 21784 36712
rect 9956 36524 10008 36533
rect 21824 36567 21876 36576
rect 21824 36533 21833 36567
rect 21833 36533 21867 36567
rect 21867 36533 21876 36567
rect 21824 36524 21876 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 22100 36363 22152 36372
rect 22100 36329 22109 36363
rect 22109 36329 22143 36363
rect 22143 36329 22152 36363
rect 23756 36363 23808 36372
rect 22100 36320 22152 36329
rect 23756 36329 23765 36363
rect 23765 36329 23799 36363
rect 23799 36329 23808 36363
rect 23756 36320 23808 36329
rect 24308 36320 24360 36372
rect 22008 36252 22060 36304
rect 1676 36159 1728 36168
rect 1676 36125 1685 36159
rect 1685 36125 1719 36159
rect 1719 36125 1728 36159
rect 1676 36116 1728 36125
rect 22008 36116 22060 36168
rect 1492 36023 1544 36032
rect 1492 35989 1501 36023
rect 1501 35989 1535 36023
rect 1535 35989 1544 36023
rect 1492 35980 1544 35989
rect 17224 35980 17276 36032
rect 35992 36116 36044 36168
rect 23020 35980 23072 36032
rect 38016 36023 38068 36032
rect 38016 35989 38025 36023
rect 38025 35989 38059 36023
rect 38059 35989 38068 36023
rect 38016 35980 38068 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 23480 35776 23532 35828
rect 24308 35776 24360 35828
rect 28448 35776 28500 35828
rect 23756 35708 23808 35760
rect 8760 35640 8812 35692
rect 38108 35683 38160 35692
rect 38108 35649 38117 35683
rect 38117 35649 38151 35683
rect 38151 35649 38160 35683
rect 38108 35640 38160 35649
rect 6552 35572 6604 35624
rect 5448 35504 5500 35556
rect 1492 35479 1544 35488
rect 1492 35445 1501 35479
rect 1501 35445 1535 35479
rect 1535 35445 1544 35479
rect 1492 35436 1544 35445
rect 2228 35479 2280 35488
rect 2228 35445 2237 35479
rect 2237 35445 2271 35479
rect 2271 35445 2280 35479
rect 2228 35436 2280 35445
rect 8760 35479 8812 35488
rect 8760 35445 8769 35479
rect 8769 35445 8803 35479
rect 8803 35445 8812 35479
rect 8760 35436 8812 35445
rect 21640 35572 21692 35624
rect 22008 35572 22060 35624
rect 23112 35572 23164 35624
rect 15200 35436 15252 35488
rect 22376 35436 22428 35488
rect 24860 35479 24912 35488
rect 24860 35445 24869 35479
rect 24869 35445 24903 35479
rect 24903 35445 24912 35479
rect 24860 35436 24912 35445
rect 37924 35479 37976 35488
rect 37924 35445 37933 35479
rect 37933 35445 37967 35479
rect 37967 35445 37976 35479
rect 37924 35436 37976 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 1676 35232 1728 35284
rect 27344 35232 27396 35284
rect 2228 35096 2280 35148
rect 2320 35071 2372 35080
rect 2320 35037 2329 35071
rect 2329 35037 2363 35071
rect 2363 35037 2372 35071
rect 2320 35028 2372 35037
rect 23756 35096 23808 35148
rect 20812 35028 20864 35080
rect 20904 35028 20956 35080
rect 24860 35071 24912 35080
rect 22100 34960 22152 35012
rect 24860 35037 24869 35071
rect 24869 35037 24903 35071
rect 24903 35037 24912 35071
rect 24860 35028 24912 35037
rect 26884 34960 26936 35012
rect 1492 34935 1544 34944
rect 1492 34901 1501 34935
rect 1501 34901 1535 34935
rect 1535 34901 1544 34935
rect 1492 34892 1544 34901
rect 22836 34935 22888 34944
rect 22836 34901 22845 34935
rect 22845 34901 22879 34935
rect 22879 34901 22888 34935
rect 22836 34892 22888 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 22376 34663 22428 34672
rect 22376 34629 22385 34663
rect 22385 34629 22419 34663
rect 22419 34629 22428 34663
rect 22376 34620 22428 34629
rect 23756 34688 23808 34740
rect 27436 34688 27488 34740
rect 36912 34688 36964 34740
rect 23664 34620 23716 34672
rect 2228 34527 2280 34536
rect 2228 34493 2237 34527
rect 2237 34493 2271 34527
rect 2271 34493 2280 34527
rect 2228 34484 2280 34493
rect 4804 34484 4856 34536
rect 27344 34595 27396 34604
rect 27344 34561 27353 34595
rect 27353 34561 27387 34595
rect 27387 34561 27396 34595
rect 27344 34552 27396 34561
rect 38108 34595 38160 34604
rect 38108 34561 38117 34595
rect 38117 34561 38151 34595
rect 38151 34561 38160 34595
rect 38108 34552 38160 34561
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 2320 34187 2372 34196
rect 2320 34153 2329 34187
rect 2329 34153 2363 34187
rect 2363 34153 2372 34187
rect 2320 34144 2372 34153
rect 22652 34144 22704 34196
rect 27344 34187 27396 34196
rect 27344 34153 27353 34187
rect 27353 34153 27387 34187
rect 27387 34153 27396 34187
rect 27344 34144 27396 34153
rect 22744 34076 22796 34128
rect 21824 34051 21876 34060
rect 1768 33940 1820 33992
rect 1676 33804 1728 33856
rect 21824 34017 21833 34051
rect 21833 34017 21867 34051
rect 21867 34017 21876 34051
rect 21824 34008 21876 34017
rect 21548 33983 21600 33992
rect 21548 33949 21557 33983
rect 21557 33949 21591 33983
rect 21591 33949 21600 33983
rect 21548 33940 21600 33949
rect 22284 33940 22336 33992
rect 4620 33804 4672 33856
rect 23756 33804 23808 33856
rect 37832 33940 37884 33992
rect 26148 33847 26200 33856
rect 26148 33813 26157 33847
rect 26157 33813 26191 33847
rect 26191 33813 26200 33847
rect 26148 33804 26200 33813
rect 36912 33872 36964 33924
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 17868 33643 17920 33652
rect 17868 33609 17877 33643
rect 17877 33609 17911 33643
rect 17911 33609 17920 33643
rect 17868 33600 17920 33609
rect 22284 33643 22336 33652
rect 22284 33609 22293 33643
rect 22293 33609 22327 33643
rect 22327 33609 22336 33643
rect 22284 33600 22336 33609
rect 22744 33643 22796 33652
rect 22744 33609 22753 33643
rect 22753 33609 22787 33643
rect 22787 33609 22796 33643
rect 22744 33600 22796 33609
rect 1400 33507 1452 33516
rect 1400 33473 1409 33507
rect 1409 33473 1443 33507
rect 1443 33473 1452 33507
rect 1400 33464 1452 33473
rect 23296 33532 23348 33584
rect 17132 33464 17184 33516
rect 5448 33396 5500 33448
rect 20260 33396 20312 33448
rect 15108 33328 15160 33380
rect 38108 33507 38160 33516
rect 38108 33473 38117 33507
rect 38117 33473 38151 33507
rect 38151 33473 38160 33507
rect 38108 33464 38160 33473
rect 5172 33260 5224 33312
rect 18236 33303 18288 33312
rect 18236 33269 18245 33303
rect 18245 33269 18279 33303
rect 18279 33269 18288 33303
rect 18236 33260 18288 33269
rect 20260 33260 20312 33312
rect 23296 33328 23348 33380
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 5448 33056 5500 33108
rect 17132 33099 17184 33108
rect 17132 33065 17141 33099
rect 17141 33065 17175 33099
rect 17175 33065 17184 33099
rect 17132 33056 17184 33065
rect 27620 33056 27672 33108
rect 35992 33056 36044 33108
rect 23388 32988 23440 33040
rect 22836 32920 22888 32972
rect 1400 32895 1452 32904
rect 1400 32861 1409 32895
rect 1409 32861 1443 32895
rect 1443 32861 1452 32895
rect 1400 32852 1452 32861
rect 22560 32852 22612 32904
rect 29368 32852 29420 32904
rect 38108 32895 38160 32904
rect 38108 32861 38117 32895
rect 38117 32861 38151 32895
rect 38151 32861 38160 32895
rect 38108 32852 38160 32861
rect 15108 32784 15160 32836
rect 21732 32784 21784 32836
rect 23756 32784 23808 32836
rect 20720 32716 20772 32768
rect 22652 32716 22704 32768
rect 36544 32716 36596 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 19248 32512 19300 32564
rect 20996 32512 21048 32564
rect 21916 32512 21968 32564
rect 22560 32555 22612 32564
rect 22560 32521 22569 32555
rect 22569 32521 22603 32555
rect 22603 32521 22612 32555
rect 22560 32512 22612 32521
rect 27068 32512 27120 32564
rect 29368 32555 29420 32564
rect 29368 32521 29377 32555
rect 29377 32521 29411 32555
rect 29411 32521 29420 32555
rect 29368 32512 29420 32521
rect 20720 32444 20772 32496
rect 23572 32487 23624 32496
rect 23572 32453 23581 32487
rect 23581 32453 23615 32487
rect 23615 32453 23624 32487
rect 23572 32444 23624 32453
rect 2688 32376 2740 32428
rect 21364 32376 21416 32428
rect 21732 32308 21784 32360
rect 23756 32351 23808 32360
rect 23756 32317 23765 32351
rect 23765 32317 23799 32351
rect 23799 32317 23808 32351
rect 23756 32308 23808 32317
rect 1492 32215 1544 32224
rect 1492 32181 1501 32215
rect 1501 32181 1535 32215
rect 1535 32181 1544 32215
rect 1492 32172 1544 32181
rect 23204 32215 23256 32224
rect 23204 32181 23213 32215
rect 23213 32181 23247 32215
rect 23247 32181 23256 32215
rect 23204 32172 23256 32181
rect 23848 32240 23900 32292
rect 38108 32419 38160 32428
rect 38108 32385 38117 32419
rect 38117 32385 38151 32419
rect 38151 32385 38160 32419
rect 38108 32376 38160 32385
rect 28724 32351 28776 32360
rect 28724 32317 28733 32351
rect 28733 32317 28767 32351
rect 28767 32317 28776 32351
rect 28724 32308 28776 32317
rect 29828 32351 29880 32360
rect 29828 32317 29837 32351
rect 29837 32317 29871 32351
rect 29871 32317 29880 32351
rect 29828 32308 29880 32317
rect 27896 32172 27948 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 2688 32011 2740 32020
rect 2688 31977 2697 32011
rect 2697 31977 2731 32011
rect 2731 31977 2740 32011
rect 2688 31968 2740 31977
rect 21364 32011 21416 32020
rect 5540 31900 5592 31952
rect 15016 31900 15068 31952
rect 4068 31832 4120 31884
rect 1400 31807 1452 31816
rect 1400 31773 1409 31807
rect 1409 31773 1443 31807
rect 1443 31773 1452 31807
rect 1400 31764 1452 31773
rect 2872 31807 2924 31816
rect 2872 31773 2881 31807
rect 2881 31773 2915 31807
rect 2915 31773 2924 31807
rect 2872 31764 2924 31773
rect 15292 31764 15344 31816
rect 19248 31900 19300 31952
rect 18236 31832 18288 31884
rect 20168 31875 20220 31884
rect 20168 31841 20177 31875
rect 20177 31841 20211 31875
rect 20211 31841 20220 31875
rect 20168 31832 20220 31841
rect 20996 31764 21048 31816
rect 21364 31977 21373 32011
rect 21373 31977 21407 32011
rect 21407 31977 21416 32011
rect 21364 31968 21416 31977
rect 21916 32011 21968 32020
rect 21916 31977 21925 32011
rect 21925 31977 21959 32011
rect 21959 31977 21968 32011
rect 21916 31968 21968 31977
rect 23112 31968 23164 32020
rect 23388 32011 23440 32020
rect 23388 31977 23397 32011
rect 23397 31977 23431 32011
rect 23431 31977 23440 32011
rect 23388 31968 23440 31977
rect 21640 31832 21692 31884
rect 22008 31764 22060 31816
rect 23112 31875 23164 31884
rect 23112 31841 23121 31875
rect 23121 31841 23155 31875
rect 23155 31841 23164 31875
rect 23112 31832 23164 31841
rect 23572 31832 23624 31884
rect 38384 31832 38436 31884
rect 28724 31764 28776 31816
rect 38016 31807 38068 31816
rect 38016 31773 38025 31807
rect 38025 31773 38059 31807
rect 38059 31773 38068 31807
rect 38016 31764 38068 31773
rect 16764 31671 16816 31680
rect 16764 31637 16773 31671
rect 16773 31637 16807 31671
rect 16807 31637 16816 31671
rect 16764 31628 16816 31637
rect 20996 31671 21048 31680
rect 20996 31637 21005 31671
rect 21005 31637 21039 31671
rect 21039 31637 21048 31671
rect 20996 31628 21048 31637
rect 23848 31628 23900 31680
rect 24308 31628 24360 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 2872 31424 2924 31476
rect 3976 31424 4028 31476
rect 20996 31424 21048 31476
rect 21732 31424 21784 31476
rect 23112 31424 23164 31476
rect 23848 31467 23900 31476
rect 23848 31433 23857 31467
rect 23857 31433 23891 31467
rect 23891 31433 23900 31467
rect 23848 31424 23900 31433
rect 2596 31356 2648 31408
rect 5448 31356 5500 31408
rect 15292 31356 15344 31408
rect 23204 31356 23256 31408
rect 5172 31331 5224 31340
rect 5172 31297 5181 31331
rect 5181 31297 5215 31331
rect 5215 31297 5224 31331
rect 5172 31288 5224 31297
rect 14280 31288 14332 31340
rect 20812 31288 20864 31340
rect 22928 31288 22980 31340
rect 1860 31263 1912 31272
rect 1860 31229 1869 31263
rect 1869 31229 1903 31263
rect 1903 31229 1912 31263
rect 1860 31220 1912 31229
rect 14556 31263 14608 31272
rect 14556 31229 14565 31263
rect 14565 31229 14599 31263
rect 14599 31229 14608 31263
rect 14556 31220 14608 31229
rect 18052 31220 18104 31272
rect 20904 31152 20956 31204
rect 37372 31152 37424 31204
rect 1584 31084 1636 31136
rect 1768 31084 1820 31136
rect 4988 31127 5040 31136
rect 4988 31093 4997 31127
rect 4997 31093 5031 31127
rect 5031 31093 5040 31127
rect 4988 31084 5040 31093
rect 15752 31084 15804 31136
rect 18236 31084 18288 31136
rect 21732 31084 21784 31136
rect 24492 31127 24544 31136
rect 24492 31093 24501 31127
rect 24501 31093 24535 31127
rect 24535 31093 24544 31127
rect 24492 31084 24544 31093
rect 37464 31084 37516 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 1400 30923 1452 30932
rect 1400 30889 1409 30923
rect 1409 30889 1443 30923
rect 1443 30889 1452 30923
rect 1400 30880 1452 30889
rect 14556 30923 14608 30932
rect 14556 30889 14565 30923
rect 14565 30889 14599 30923
rect 14599 30889 14608 30923
rect 14556 30880 14608 30889
rect 17224 30812 17276 30864
rect 14280 30744 14332 30796
rect 15752 30787 15804 30796
rect 15752 30753 15761 30787
rect 15761 30753 15795 30787
rect 15795 30753 15804 30787
rect 15752 30744 15804 30753
rect 24492 30812 24544 30864
rect 16764 30608 16816 30660
rect 22468 30583 22520 30592
rect 22468 30549 22477 30583
rect 22477 30549 22511 30583
rect 22511 30549 22520 30583
rect 22468 30540 22520 30549
rect 23020 30583 23072 30592
rect 23020 30549 23029 30583
rect 23029 30549 23063 30583
rect 23063 30549 23072 30583
rect 23020 30540 23072 30549
rect 24308 30540 24360 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 23020 30268 23072 30320
rect 23664 30268 23716 30320
rect 17224 30200 17276 30252
rect 22744 30132 22796 30184
rect 23020 30132 23072 30184
rect 21180 30064 21232 30116
rect 27528 30243 27580 30252
rect 24860 30132 24912 30184
rect 1492 30039 1544 30048
rect 1492 30005 1501 30039
rect 1501 30005 1535 30039
rect 1535 30005 1544 30039
rect 1492 29996 1544 30005
rect 23848 29996 23900 30048
rect 27528 30209 27537 30243
rect 27537 30209 27571 30243
rect 27571 30209 27580 30243
rect 27528 30200 27580 30209
rect 30380 30200 30432 30252
rect 37924 30064 37976 30116
rect 26056 29996 26108 30048
rect 26976 30039 27028 30048
rect 26976 30005 26985 30039
rect 26985 30005 27019 30039
rect 27019 30005 27028 30039
rect 26976 29996 27028 30005
rect 30932 29996 30984 30048
rect 38016 30039 38068 30048
rect 38016 30005 38025 30039
rect 38025 30005 38059 30039
rect 38059 30005 38068 30039
rect 38016 29996 38068 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 21088 29792 21140 29844
rect 16948 29724 17000 29776
rect 23388 29792 23440 29844
rect 23664 29792 23716 29844
rect 27528 29835 27580 29844
rect 27528 29801 27537 29835
rect 27537 29801 27571 29835
rect 27571 29801 27580 29835
rect 27528 29792 27580 29801
rect 34612 29792 34664 29844
rect 22192 29724 22244 29776
rect 22284 29724 22336 29776
rect 23112 29724 23164 29776
rect 26976 29699 27028 29708
rect 4988 29588 5040 29640
rect 20444 29631 20496 29640
rect 20444 29597 20453 29631
rect 20453 29597 20487 29631
rect 20487 29597 20496 29631
rect 20444 29588 20496 29597
rect 22192 29588 22244 29640
rect 9036 29520 9088 29572
rect 20536 29520 20588 29572
rect 1492 29495 1544 29504
rect 1492 29461 1501 29495
rect 1501 29461 1535 29495
rect 1535 29461 1544 29495
rect 1492 29452 1544 29461
rect 22560 29452 22612 29504
rect 26976 29665 26985 29699
rect 26985 29665 27019 29699
rect 27019 29665 27028 29699
rect 26976 29656 27028 29665
rect 23848 29588 23900 29640
rect 36728 29656 36780 29708
rect 34244 29588 34296 29640
rect 38108 29631 38160 29640
rect 38108 29597 38117 29631
rect 38117 29597 38151 29631
rect 38151 29597 38160 29631
rect 38108 29588 38160 29597
rect 23112 29520 23164 29572
rect 24768 29563 24820 29572
rect 24768 29529 24777 29563
rect 24777 29529 24811 29563
rect 24811 29529 24820 29563
rect 24768 29520 24820 29529
rect 26056 29452 26108 29504
rect 27068 29495 27120 29504
rect 27068 29461 27077 29495
rect 27077 29461 27111 29495
rect 27111 29461 27120 29495
rect 27068 29452 27120 29461
rect 27988 29495 28040 29504
rect 27988 29461 27997 29495
rect 27997 29461 28031 29495
rect 28031 29461 28040 29495
rect 27988 29452 28040 29461
rect 37924 29495 37976 29504
rect 37924 29461 37933 29495
rect 37933 29461 37967 29495
rect 37967 29461 37976 29495
rect 37924 29452 37976 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 1400 29155 1452 29164
rect 1400 29121 1409 29155
rect 1409 29121 1443 29155
rect 1443 29121 1452 29155
rect 1400 29112 1452 29121
rect 19340 29248 19392 29300
rect 20352 29248 20404 29300
rect 22192 29291 22244 29300
rect 22192 29257 22201 29291
rect 22201 29257 22235 29291
rect 22235 29257 22244 29291
rect 22192 29248 22244 29257
rect 23296 29248 23348 29300
rect 23388 29248 23440 29300
rect 27068 29291 27120 29300
rect 27068 29257 27077 29291
rect 27077 29257 27111 29291
rect 27111 29257 27120 29291
rect 27068 29248 27120 29257
rect 34244 29291 34296 29300
rect 34244 29257 34253 29291
rect 34253 29257 34287 29291
rect 34287 29257 34296 29291
rect 34244 29248 34296 29257
rect 15200 29180 15252 29232
rect 22468 29180 22520 29232
rect 4620 29044 4672 29096
rect 5264 29044 5316 29096
rect 20812 29112 20864 29164
rect 37924 29180 37976 29232
rect 18604 29044 18656 29096
rect 20536 29087 20588 29096
rect 20536 29053 20545 29087
rect 20545 29053 20579 29087
rect 20579 29053 20588 29087
rect 20536 29044 20588 29053
rect 22560 28976 22612 29028
rect 23296 29044 23348 29096
rect 26976 29044 27028 29096
rect 33600 29087 33652 29096
rect 33600 29053 33609 29087
rect 33609 29053 33643 29087
rect 33643 29053 33652 29087
rect 33600 29044 33652 29053
rect 38108 29155 38160 29164
rect 38108 29121 38117 29155
rect 38117 29121 38151 29155
rect 38151 29121 38160 29155
rect 38108 29112 38160 29121
rect 23204 28976 23256 29028
rect 32956 29019 33008 29028
rect 32956 28985 32965 29019
rect 32965 28985 32999 29019
rect 32999 28985 33008 29019
rect 37556 29044 37608 29096
rect 32956 28976 33008 28985
rect 36636 28976 36688 29028
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 20812 28747 20864 28756
rect 20812 28713 20821 28747
rect 20821 28713 20855 28747
rect 20855 28713 20864 28747
rect 20812 28704 20864 28713
rect 33416 28747 33468 28756
rect 33416 28713 33425 28747
rect 33425 28713 33459 28747
rect 33459 28713 33468 28747
rect 33416 28704 33468 28713
rect 33600 28704 33652 28756
rect 4712 28636 4764 28688
rect 25964 28636 26016 28688
rect 19432 28568 19484 28620
rect 20168 28568 20220 28620
rect 22468 28568 22520 28620
rect 3240 28500 3292 28552
rect 20352 28432 20404 28484
rect 21916 28432 21968 28484
rect 4620 28364 4672 28416
rect 19432 28364 19484 28416
rect 20168 28407 20220 28416
rect 20168 28373 20177 28407
rect 20177 28373 20211 28407
rect 20211 28373 20220 28407
rect 20168 28364 20220 28373
rect 22100 28364 22152 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 5356 28203 5408 28212
rect 5356 28169 5365 28203
rect 5365 28169 5399 28203
rect 5399 28169 5408 28203
rect 5356 28160 5408 28169
rect 19340 28203 19392 28212
rect 19340 28169 19349 28203
rect 19349 28169 19383 28203
rect 19383 28169 19392 28203
rect 19340 28160 19392 28169
rect 20444 28160 20496 28212
rect 21916 28203 21968 28212
rect 21916 28169 21925 28203
rect 21925 28169 21959 28203
rect 21959 28169 21968 28203
rect 21916 28160 21968 28169
rect 23112 28160 23164 28212
rect 22008 28092 22060 28144
rect 1400 28067 1452 28076
rect 1400 28033 1409 28067
rect 1409 28033 1443 28067
rect 1443 28033 1452 28067
rect 1400 28024 1452 28033
rect 21272 28024 21324 28076
rect 4620 27956 4672 28008
rect 20168 27956 20220 28008
rect 25320 28024 25372 28076
rect 26056 28024 26108 28076
rect 22468 27999 22520 28008
rect 22468 27965 22477 27999
rect 22477 27965 22511 27999
rect 22511 27965 22520 27999
rect 22468 27956 22520 27965
rect 25964 27999 26016 28008
rect 25964 27965 25973 27999
rect 25973 27965 26007 27999
rect 26007 27965 26016 27999
rect 25964 27956 26016 27965
rect 4896 27863 4948 27872
rect 4896 27829 4905 27863
rect 4905 27829 4939 27863
rect 4939 27829 4948 27863
rect 4896 27820 4948 27829
rect 23480 27820 23532 27872
rect 26148 27820 26200 27872
rect 38016 27931 38068 27940
rect 38016 27897 38025 27931
rect 38025 27897 38059 27931
rect 38059 27897 38068 27931
rect 38016 27888 38068 27897
rect 37556 27820 37608 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 20352 27616 20404 27668
rect 1860 27548 1912 27600
rect 20996 27591 21048 27600
rect 20996 27557 21005 27591
rect 21005 27557 21039 27591
rect 21039 27557 21048 27591
rect 23112 27616 23164 27668
rect 20996 27548 21048 27557
rect 19432 27480 19484 27532
rect 1400 27455 1452 27464
rect 1400 27421 1409 27455
rect 1409 27421 1443 27455
rect 1443 27421 1452 27455
rect 1400 27412 1452 27421
rect 4896 27412 4948 27464
rect 5448 27387 5500 27396
rect 5448 27353 5457 27387
rect 5457 27353 5491 27387
rect 5491 27353 5500 27387
rect 5448 27344 5500 27353
rect 3240 27276 3292 27328
rect 20904 27412 20956 27464
rect 23112 27412 23164 27464
rect 17960 27344 18012 27396
rect 19984 27319 20036 27328
rect 19984 27285 19993 27319
rect 19993 27285 20027 27319
rect 20027 27285 20036 27319
rect 19984 27276 20036 27285
rect 20444 27319 20496 27328
rect 20444 27285 20453 27319
rect 20453 27285 20487 27319
rect 20487 27285 20496 27319
rect 20444 27276 20496 27285
rect 21916 27319 21968 27328
rect 21916 27285 21925 27319
rect 21925 27285 21959 27319
rect 21959 27285 21968 27319
rect 21916 27276 21968 27285
rect 37280 27319 37332 27328
rect 37280 27285 37289 27319
rect 37289 27285 37323 27319
rect 37323 27285 37332 27319
rect 37280 27276 37332 27285
rect 38016 27319 38068 27328
rect 38016 27285 38025 27319
rect 38025 27285 38059 27319
rect 38059 27285 38068 27319
rect 38016 27276 38068 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 14648 27072 14700 27124
rect 19984 27072 20036 27124
rect 5632 27004 5684 27056
rect 21180 27004 21232 27056
rect 14832 26936 14884 26988
rect 20444 26936 20496 26988
rect 22284 27072 22336 27124
rect 23112 27072 23164 27124
rect 38108 26979 38160 26988
rect 4068 26868 4120 26920
rect 6368 26868 6420 26920
rect 18604 26868 18656 26920
rect 38108 26945 38117 26979
rect 38117 26945 38151 26979
rect 38151 26945 38160 26979
rect 38108 26936 38160 26945
rect 20996 26911 21048 26920
rect 20996 26877 21005 26911
rect 21005 26877 21039 26911
rect 21039 26877 21048 26911
rect 20996 26868 21048 26877
rect 21640 26868 21692 26920
rect 1492 26775 1544 26784
rect 1492 26741 1501 26775
rect 1501 26741 1535 26775
rect 1535 26741 1544 26775
rect 1492 26732 1544 26741
rect 19432 26732 19484 26784
rect 23204 26775 23256 26784
rect 23204 26741 23213 26775
rect 23213 26741 23247 26775
rect 23247 26741 23256 26775
rect 23204 26732 23256 26741
rect 37280 26732 37332 26784
rect 37924 26775 37976 26784
rect 37924 26741 37933 26775
rect 37933 26741 37967 26775
rect 37967 26741 37976 26775
rect 37924 26732 37976 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 18604 26571 18656 26580
rect 18604 26537 18613 26571
rect 18613 26537 18647 26571
rect 18647 26537 18656 26571
rect 18604 26528 18656 26537
rect 20904 26571 20956 26580
rect 20904 26537 20913 26571
rect 20913 26537 20947 26571
rect 20947 26537 20956 26571
rect 20904 26528 20956 26537
rect 21456 26460 21508 26512
rect 23388 26528 23440 26580
rect 26424 26460 26476 26512
rect 38016 26503 38068 26512
rect 38016 26469 38025 26503
rect 38025 26469 38059 26503
rect 38059 26469 38068 26503
rect 38016 26460 38068 26469
rect 23204 26392 23256 26444
rect 37924 26392 37976 26444
rect 3332 26324 3384 26376
rect 21732 26324 21784 26376
rect 27712 26324 27764 26376
rect 38568 26324 38620 26376
rect 1492 26231 1544 26240
rect 1492 26197 1501 26231
rect 1501 26197 1535 26231
rect 1535 26197 1544 26231
rect 1492 26188 1544 26197
rect 23388 26231 23440 26240
rect 23388 26197 23397 26231
rect 23397 26197 23431 26231
rect 23431 26197 23440 26231
rect 23388 26188 23440 26197
rect 30380 26256 30432 26308
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 18972 25984 19024 26036
rect 20996 25984 21048 26036
rect 23848 26027 23900 26036
rect 23848 25993 23857 26027
rect 23857 25993 23891 26027
rect 23891 25993 23900 26027
rect 23848 25984 23900 25993
rect 26424 26027 26476 26036
rect 26424 25993 26433 26027
rect 26433 25993 26467 26027
rect 26467 25993 26476 26027
rect 26424 25984 26476 25993
rect 27712 26027 27764 26036
rect 27712 25993 27721 26027
rect 27721 25993 27755 26027
rect 27755 25993 27764 26027
rect 27712 25984 27764 25993
rect 18144 25891 18196 25900
rect 18144 25857 18153 25891
rect 18153 25857 18187 25891
rect 18187 25857 18196 25891
rect 18144 25848 18196 25857
rect 18604 25848 18656 25900
rect 22376 25848 22428 25900
rect 19432 25780 19484 25832
rect 20628 25780 20680 25832
rect 22468 25823 22520 25832
rect 22468 25789 22477 25823
rect 22477 25789 22511 25823
rect 22511 25789 22520 25823
rect 22468 25780 22520 25789
rect 22560 25823 22612 25832
rect 22560 25789 22569 25823
rect 22569 25789 22603 25823
rect 22603 25789 22612 25823
rect 27068 25823 27120 25832
rect 22560 25780 22612 25789
rect 27068 25789 27077 25823
rect 27077 25789 27111 25823
rect 27111 25789 27120 25823
rect 27068 25780 27120 25789
rect 37924 25780 37976 25832
rect 21640 25712 21692 25764
rect 36636 25712 36688 25764
rect 1860 25644 1912 25696
rect 2320 25644 2372 25696
rect 18052 25644 18104 25696
rect 20352 25687 20404 25696
rect 20352 25653 20361 25687
rect 20361 25653 20395 25687
rect 20395 25653 20404 25687
rect 20352 25644 20404 25653
rect 22652 25644 22704 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 25320 25440 25372 25492
rect 37924 25483 37976 25492
rect 37924 25449 37933 25483
rect 37933 25449 37967 25483
rect 37967 25449 37976 25483
rect 37924 25440 37976 25449
rect 20628 25372 20680 25424
rect 18972 25304 19024 25356
rect 20996 25304 21048 25356
rect 21640 25347 21692 25356
rect 21640 25313 21649 25347
rect 21649 25313 21683 25347
rect 21683 25313 21692 25347
rect 21640 25304 21692 25313
rect 22284 25372 22336 25424
rect 24400 25415 24452 25424
rect 24400 25381 24409 25415
rect 24409 25381 24443 25415
rect 24443 25381 24452 25415
rect 24400 25372 24452 25381
rect 22928 25347 22980 25356
rect 22928 25313 22937 25347
rect 22937 25313 22971 25347
rect 22971 25313 22980 25347
rect 22928 25304 22980 25313
rect 1860 25279 1912 25288
rect 1860 25245 1869 25279
rect 1869 25245 1903 25279
rect 1903 25245 1912 25279
rect 1860 25236 1912 25245
rect 18144 25236 18196 25288
rect 20352 25236 20404 25288
rect 23112 25236 23164 25288
rect 23664 25236 23716 25288
rect 2596 25168 2648 25220
rect 18236 25211 18288 25220
rect 18236 25177 18245 25211
rect 18245 25177 18279 25211
rect 18279 25177 18288 25211
rect 18236 25168 18288 25177
rect 19340 25168 19392 25220
rect 19248 25143 19300 25152
rect 19248 25109 19257 25143
rect 19257 25109 19291 25143
rect 19291 25109 19300 25143
rect 19248 25100 19300 25109
rect 20628 25100 20680 25152
rect 21180 25143 21232 25152
rect 21180 25109 21189 25143
rect 21189 25109 21223 25143
rect 21223 25109 21232 25143
rect 21180 25100 21232 25109
rect 35440 25236 35492 25288
rect 38108 25279 38160 25288
rect 38108 25245 38117 25279
rect 38117 25245 38151 25279
rect 38151 25245 38160 25279
rect 38108 25236 38160 25245
rect 25044 25211 25096 25220
rect 25044 25177 25053 25211
rect 25053 25177 25087 25211
rect 25087 25177 25096 25211
rect 25044 25168 25096 25177
rect 24400 25100 24452 25152
rect 26240 25100 26292 25152
rect 27068 25100 27120 25152
rect 37832 25100 37884 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 22008 24939 22060 24948
rect 22008 24905 22017 24939
rect 22017 24905 22051 24939
rect 22051 24905 22060 24939
rect 22008 24896 22060 24905
rect 23664 24939 23716 24948
rect 23664 24905 23673 24939
rect 23673 24905 23707 24939
rect 23707 24905 23716 24939
rect 23664 24896 23716 24905
rect 23388 24828 23440 24880
rect 25044 24828 25096 24880
rect 1400 24803 1452 24812
rect 1400 24769 1409 24803
rect 1409 24769 1443 24803
rect 1443 24769 1452 24803
rect 1400 24760 1452 24769
rect 17960 24803 18012 24812
rect 17960 24769 17969 24803
rect 17969 24769 18003 24803
rect 18003 24769 18012 24803
rect 17960 24760 18012 24769
rect 19248 24803 19300 24812
rect 19248 24769 19257 24803
rect 19257 24769 19291 24803
rect 19291 24769 19300 24803
rect 19248 24760 19300 24769
rect 21180 24760 21232 24812
rect 21824 24803 21876 24812
rect 21824 24769 21833 24803
rect 21833 24769 21867 24803
rect 21867 24769 21876 24803
rect 21824 24760 21876 24769
rect 18972 24735 19024 24744
rect 18972 24701 18981 24735
rect 18981 24701 19015 24735
rect 19015 24701 19024 24735
rect 18972 24692 19024 24701
rect 20996 24735 21048 24744
rect 20996 24701 21005 24735
rect 21005 24701 21039 24735
rect 21039 24701 21048 24735
rect 20996 24692 21048 24701
rect 21088 24692 21140 24744
rect 22284 24692 22336 24744
rect 23112 24556 23164 24608
rect 25320 24803 25372 24812
rect 25320 24769 25329 24803
rect 25329 24769 25363 24803
rect 25363 24769 25372 24803
rect 25320 24760 25372 24769
rect 24216 24735 24268 24744
rect 24216 24701 24225 24735
rect 24225 24701 24259 24735
rect 24259 24701 24268 24735
rect 24216 24692 24268 24701
rect 24768 24692 24820 24744
rect 25228 24624 25280 24676
rect 33416 24692 33468 24744
rect 38108 24803 38160 24812
rect 38108 24769 38117 24803
rect 38117 24769 38151 24803
rect 38151 24769 38160 24803
rect 38108 24760 38160 24769
rect 27896 24599 27948 24608
rect 27896 24565 27905 24599
rect 27905 24565 27939 24599
rect 27939 24565 27948 24599
rect 27896 24556 27948 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 19340 24395 19392 24404
rect 19340 24361 19349 24395
rect 19349 24361 19383 24395
rect 19383 24361 19392 24395
rect 19340 24352 19392 24361
rect 22560 24352 22612 24404
rect 24768 24395 24820 24404
rect 24768 24361 24777 24395
rect 24777 24361 24811 24395
rect 24811 24361 24820 24395
rect 24768 24352 24820 24361
rect 16212 24284 16264 24336
rect 21916 24284 21968 24336
rect 13636 24148 13688 24200
rect 18328 24191 18380 24200
rect 18328 24157 18337 24191
rect 18337 24157 18371 24191
rect 18371 24157 18380 24191
rect 18328 24148 18380 24157
rect 21456 24259 21508 24268
rect 21456 24225 21465 24259
rect 21465 24225 21499 24259
rect 21499 24225 21508 24259
rect 21456 24216 21508 24225
rect 23204 24216 23256 24268
rect 19432 24148 19484 24200
rect 20076 24148 20128 24200
rect 22468 24148 22520 24200
rect 22744 24191 22796 24200
rect 22744 24157 22753 24191
rect 22753 24157 22787 24191
rect 22787 24157 22796 24191
rect 22744 24148 22796 24157
rect 24492 24148 24544 24200
rect 24860 24191 24912 24200
rect 1860 24123 1912 24132
rect 1860 24089 1869 24123
rect 1869 24089 1903 24123
rect 1903 24089 1912 24123
rect 1860 24080 1912 24089
rect 2044 24123 2096 24132
rect 2044 24089 2053 24123
rect 2053 24089 2087 24123
rect 2087 24089 2096 24123
rect 2044 24080 2096 24089
rect 2228 24080 2280 24132
rect 17960 24080 18012 24132
rect 20904 24080 20956 24132
rect 21916 24080 21968 24132
rect 18696 24055 18748 24064
rect 18696 24021 18705 24055
rect 18705 24021 18739 24055
rect 18739 24021 18748 24055
rect 18696 24012 18748 24021
rect 22376 24080 22428 24132
rect 24860 24157 24869 24191
rect 24869 24157 24903 24191
rect 24903 24157 24912 24191
rect 24860 24148 24912 24157
rect 27896 24216 27948 24268
rect 36544 24352 36596 24404
rect 37648 24216 37700 24268
rect 29460 24148 29512 24200
rect 23296 24012 23348 24064
rect 24400 24055 24452 24064
rect 24400 24021 24409 24055
rect 24409 24021 24443 24055
rect 24443 24021 24452 24055
rect 24400 24012 24452 24021
rect 25228 24012 25280 24064
rect 28540 24012 28592 24064
rect 38016 24055 38068 24064
rect 38016 24021 38025 24055
rect 38025 24021 38059 24055
rect 38059 24021 38068 24055
rect 38016 24012 38068 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 13636 23851 13688 23860
rect 13636 23817 13645 23851
rect 13645 23817 13679 23851
rect 13679 23817 13688 23851
rect 13636 23808 13688 23817
rect 21548 23808 21600 23860
rect 21824 23851 21876 23860
rect 21824 23817 21833 23851
rect 21833 23817 21867 23851
rect 21867 23817 21876 23851
rect 21824 23808 21876 23817
rect 21916 23808 21968 23860
rect 24216 23808 24268 23860
rect 18144 23740 18196 23792
rect 8208 23604 8260 23656
rect 14556 23604 14608 23656
rect 1492 23511 1544 23520
rect 1492 23477 1501 23511
rect 1501 23477 1535 23511
rect 1535 23477 1544 23511
rect 1492 23468 1544 23477
rect 17960 23672 18012 23724
rect 18236 23672 18288 23724
rect 18696 23672 18748 23724
rect 24400 23740 24452 23792
rect 21732 23672 21784 23724
rect 23112 23715 23164 23724
rect 23112 23681 23121 23715
rect 23121 23681 23155 23715
rect 23155 23681 23164 23715
rect 23112 23672 23164 23681
rect 19432 23647 19484 23656
rect 15200 23468 15252 23520
rect 19432 23613 19441 23647
rect 19441 23613 19475 23647
rect 19475 23613 19484 23647
rect 19432 23604 19484 23613
rect 22284 23647 22336 23656
rect 19340 23536 19392 23588
rect 22284 23613 22293 23647
rect 22293 23613 22327 23647
rect 22327 23613 22336 23647
rect 22284 23604 22336 23613
rect 22376 23647 22428 23656
rect 22376 23613 22385 23647
rect 22385 23613 22419 23647
rect 22419 23613 22428 23647
rect 23388 23647 23440 23656
rect 22376 23604 22428 23613
rect 23388 23613 23397 23647
rect 23397 23613 23431 23647
rect 23431 23613 23440 23647
rect 23388 23604 23440 23613
rect 22560 23536 22612 23588
rect 23296 23536 23348 23588
rect 24860 23808 24912 23860
rect 29460 23851 29512 23860
rect 29460 23817 29469 23851
rect 29469 23817 29503 23851
rect 29503 23817 29512 23851
rect 29460 23808 29512 23817
rect 37372 23851 37424 23860
rect 37372 23817 37381 23851
rect 37381 23817 37415 23851
rect 37415 23817 37424 23851
rect 37372 23808 37424 23817
rect 27896 23604 27948 23656
rect 22376 23468 22428 23520
rect 24492 23468 24544 23520
rect 29920 23511 29972 23520
rect 29920 23477 29929 23511
rect 29929 23477 29963 23511
rect 29963 23477 29972 23511
rect 29920 23468 29972 23477
rect 38016 23511 38068 23520
rect 38016 23477 38025 23511
rect 38025 23477 38059 23511
rect 38059 23477 38068 23511
rect 38016 23468 38068 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 18328 23264 18380 23316
rect 18604 23307 18656 23316
rect 18604 23273 18613 23307
rect 18613 23273 18647 23307
rect 18647 23273 18656 23307
rect 18604 23264 18656 23273
rect 19432 23264 19484 23316
rect 20076 23264 20128 23316
rect 24860 23264 24912 23316
rect 27896 23307 27948 23316
rect 27896 23273 27905 23307
rect 27905 23273 27939 23307
rect 27939 23273 27948 23307
rect 27896 23264 27948 23273
rect 5080 23196 5132 23248
rect 10324 23171 10376 23180
rect 10324 23137 10333 23171
rect 10333 23137 10367 23171
rect 10367 23137 10376 23171
rect 10324 23128 10376 23137
rect 10232 23060 10284 23112
rect 20628 23196 20680 23248
rect 15200 23128 15252 23180
rect 16672 23060 16724 23112
rect 18512 23128 18564 23180
rect 19984 23128 20036 23180
rect 20904 23128 20956 23180
rect 22560 23196 22612 23248
rect 26240 23196 26292 23248
rect 26792 23196 26844 23248
rect 22376 23128 22428 23180
rect 23020 23128 23072 23180
rect 22928 23060 22980 23112
rect 28540 23103 28592 23112
rect 28540 23069 28549 23103
rect 28549 23069 28583 23103
rect 28583 23069 28592 23103
rect 28540 23060 28592 23069
rect 19524 22992 19576 23044
rect 20260 22992 20312 23044
rect 23664 22992 23716 23044
rect 14556 22967 14608 22976
rect 14556 22933 14565 22967
rect 14565 22933 14599 22967
rect 14599 22933 14608 22967
rect 14556 22924 14608 22933
rect 18604 22924 18656 22976
rect 20904 22967 20956 22976
rect 20904 22933 20913 22967
rect 20913 22933 20947 22967
rect 20947 22933 20956 22967
rect 20904 22924 20956 22933
rect 21640 22924 21692 22976
rect 22284 22924 22336 22976
rect 23296 22924 23348 22976
rect 30840 22924 30892 22976
rect 38108 22967 38160 22976
rect 38108 22933 38117 22967
rect 38117 22933 38151 22967
rect 38151 22933 38160 22967
rect 38108 22924 38160 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 10232 22763 10284 22772
rect 10232 22729 10241 22763
rect 10241 22729 10275 22763
rect 10275 22729 10284 22763
rect 10232 22720 10284 22729
rect 16672 22763 16724 22772
rect 16672 22729 16681 22763
rect 16681 22729 16715 22763
rect 16715 22729 16724 22763
rect 16672 22720 16724 22729
rect 18512 22720 18564 22772
rect 19984 22720 20036 22772
rect 20076 22720 20128 22772
rect 20260 22763 20312 22772
rect 20260 22729 20269 22763
rect 20269 22729 20303 22763
rect 20303 22729 20312 22763
rect 20260 22720 20312 22729
rect 20904 22720 20956 22772
rect 21272 22720 21324 22772
rect 21732 22720 21784 22772
rect 22468 22763 22520 22772
rect 22468 22729 22477 22763
rect 22477 22729 22511 22763
rect 22511 22729 22520 22763
rect 22468 22720 22520 22729
rect 23572 22763 23624 22772
rect 23572 22729 23581 22763
rect 23581 22729 23615 22763
rect 23615 22729 23624 22763
rect 23572 22720 23624 22729
rect 14556 22652 14608 22704
rect 20628 22652 20680 22704
rect 1400 22627 1452 22636
rect 1400 22593 1409 22627
rect 1409 22593 1443 22627
rect 1443 22593 1452 22627
rect 1400 22584 1452 22593
rect 10508 22584 10560 22636
rect 24584 22652 24636 22704
rect 11152 22516 11204 22568
rect 17132 22559 17184 22568
rect 17132 22525 17141 22559
rect 17141 22525 17175 22559
rect 17175 22525 17184 22559
rect 17132 22516 17184 22525
rect 17316 22559 17368 22568
rect 17316 22525 17325 22559
rect 17325 22525 17359 22559
rect 17359 22525 17368 22559
rect 17316 22516 17368 22525
rect 22928 22627 22980 22636
rect 21456 22516 21508 22568
rect 22928 22593 22937 22627
rect 22937 22593 22971 22627
rect 22971 22593 22980 22627
rect 22928 22584 22980 22593
rect 23296 22584 23348 22636
rect 22836 22516 22888 22568
rect 24676 22516 24728 22568
rect 38108 22559 38160 22568
rect 38108 22525 38117 22559
rect 38117 22525 38151 22559
rect 38151 22525 38160 22559
rect 38108 22516 38160 22525
rect 1584 22423 1636 22432
rect 1584 22389 1593 22423
rect 1593 22389 1627 22423
rect 1627 22389 1636 22423
rect 1584 22380 1636 22389
rect 23664 22380 23716 22432
rect 24768 22380 24820 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 1584 22176 1636 22228
rect 17132 22176 17184 22228
rect 23572 22176 23624 22228
rect 37372 22176 37424 22228
rect 11152 22083 11204 22092
rect 11152 22049 11161 22083
rect 11161 22049 11195 22083
rect 11195 22049 11204 22083
rect 11152 22040 11204 22049
rect 17960 22040 18012 22092
rect 21088 22040 21140 22092
rect 22376 22040 22428 22092
rect 22468 22083 22520 22092
rect 22468 22049 22477 22083
rect 22477 22049 22511 22083
rect 22511 22049 22520 22083
rect 22468 22040 22520 22049
rect 1400 22015 1452 22024
rect 1400 21981 1409 22015
rect 1409 21981 1443 22015
rect 1443 21981 1452 22015
rect 1400 21972 1452 21981
rect 38108 22015 38160 22024
rect 38108 21981 38117 22015
rect 38117 21981 38151 22015
rect 38151 21981 38160 22015
rect 38108 21972 38160 21981
rect 1676 21836 1728 21888
rect 3056 21836 3108 21888
rect 17316 21836 17368 21888
rect 17592 21879 17644 21888
rect 17592 21845 17601 21879
rect 17601 21845 17635 21879
rect 17635 21845 17644 21879
rect 17592 21836 17644 21845
rect 20352 21879 20404 21888
rect 20352 21845 20361 21879
rect 20361 21845 20395 21879
rect 20395 21845 20404 21879
rect 20352 21836 20404 21845
rect 22928 21879 22980 21888
rect 22928 21845 22937 21879
rect 22937 21845 22971 21879
rect 22971 21845 22980 21879
rect 22928 21836 22980 21845
rect 24768 21836 24820 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 5356 21632 5408 21684
rect 4068 21496 4120 21548
rect 20352 21496 20404 21548
rect 37924 21496 37976 21548
rect 2044 21428 2096 21480
rect 17592 21360 17644 21412
rect 21088 21360 21140 21412
rect 20536 21292 20588 21344
rect 24308 21360 24360 21412
rect 37280 21360 37332 21412
rect 21732 21292 21784 21344
rect 38016 21335 38068 21344
rect 38016 21301 38025 21335
rect 38025 21301 38059 21335
rect 38059 21301 38068 21335
rect 38016 21292 38068 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 2044 21131 2096 21140
rect 2044 21097 2053 21131
rect 2053 21097 2087 21131
rect 2087 21097 2096 21131
rect 2044 21088 2096 21097
rect 37832 21088 37884 21140
rect 5356 20952 5408 21004
rect 37280 20952 37332 21004
rect 37832 20952 37884 21004
rect 1400 20927 1452 20936
rect 1400 20893 1409 20927
rect 1409 20893 1443 20927
rect 1443 20893 1452 20927
rect 1400 20884 1452 20893
rect 6460 20927 6512 20936
rect 6460 20893 6469 20927
rect 6469 20893 6503 20927
rect 6503 20893 6512 20927
rect 6460 20884 6512 20893
rect 38108 20927 38160 20936
rect 38108 20893 38117 20927
rect 38117 20893 38151 20927
rect 38151 20893 38160 20927
rect 38108 20884 38160 20893
rect 7472 20791 7524 20800
rect 7472 20757 7481 20791
rect 7481 20757 7515 20791
rect 7515 20757 7524 20791
rect 7472 20748 7524 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 6460 20544 6512 20596
rect 33416 20544 33468 20596
rect 1400 20519 1452 20528
rect 1400 20485 1409 20519
rect 1409 20485 1443 20519
rect 1443 20485 1452 20519
rect 1400 20476 1452 20485
rect 1584 20408 1636 20460
rect 36268 20408 36320 20460
rect 3516 20383 3568 20392
rect 3516 20349 3525 20383
rect 3525 20349 3559 20383
rect 3559 20349 3568 20383
rect 3516 20340 3568 20349
rect 33784 20340 33836 20392
rect 32588 20272 32640 20324
rect 2228 20204 2280 20256
rect 2872 20247 2924 20256
rect 2872 20213 2881 20247
rect 2881 20213 2915 20247
rect 2915 20213 2924 20247
rect 2872 20204 2924 20213
rect 12808 20204 12860 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 3516 20000 3568 20052
rect 5356 20000 5408 20052
rect 12256 20043 12308 20052
rect 12256 20009 12265 20043
rect 12265 20009 12299 20043
rect 12299 20009 12308 20043
rect 12256 20000 12308 20009
rect 13176 20000 13228 20052
rect 14556 20000 14608 20052
rect 21916 20000 21968 20052
rect 5448 19932 5500 19984
rect 14556 19864 14608 19916
rect 1952 19839 2004 19848
rect 1952 19805 1961 19839
rect 1961 19805 1995 19839
rect 1995 19805 2004 19839
rect 1952 19796 2004 19805
rect 2228 19839 2280 19848
rect 2228 19805 2237 19839
rect 2237 19805 2271 19839
rect 2271 19805 2280 19839
rect 2228 19796 2280 19805
rect 2872 19839 2924 19848
rect 2872 19805 2881 19839
rect 2881 19805 2915 19839
rect 2915 19805 2924 19839
rect 2872 19796 2924 19805
rect 12808 19796 12860 19848
rect 2596 19728 2648 19780
rect 1676 19660 1728 19712
rect 12716 19660 12768 19712
rect 13176 19703 13228 19712
rect 13176 19669 13185 19703
rect 13185 19669 13219 19703
rect 13219 19669 13228 19703
rect 22928 19796 22980 19848
rect 33140 19864 33192 19916
rect 33416 19864 33468 19916
rect 35440 19796 35492 19848
rect 13176 19660 13228 19669
rect 34244 19660 34296 19712
rect 38016 19703 38068 19712
rect 38016 19669 38025 19703
rect 38025 19669 38059 19703
rect 38059 19669 38068 19703
rect 38016 19660 38068 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 3332 19499 3384 19508
rect 3332 19465 3341 19499
rect 3341 19465 3375 19499
rect 3375 19465 3384 19499
rect 3332 19456 3384 19465
rect 33784 19499 33836 19508
rect 33784 19465 33793 19499
rect 33793 19465 33827 19499
rect 33827 19465 33836 19499
rect 33784 19456 33836 19465
rect 1676 19363 1728 19372
rect 1676 19329 1685 19363
rect 1685 19329 1719 19363
rect 1719 19329 1728 19363
rect 1676 19320 1728 19329
rect 3516 19363 3568 19372
rect 3516 19329 3525 19363
rect 3525 19329 3559 19363
rect 3559 19329 3568 19363
rect 3516 19320 3568 19329
rect 12716 19363 12768 19372
rect 12716 19329 12725 19363
rect 12725 19329 12759 19363
rect 12759 19329 12768 19363
rect 12716 19320 12768 19329
rect 22284 19363 22336 19372
rect 22284 19329 22293 19363
rect 22293 19329 22327 19363
rect 22327 19329 22336 19363
rect 22284 19320 22336 19329
rect 23756 19320 23808 19372
rect 34244 19363 34296 19372
rect 21916 19252 21968 19304
rect 33140 19295 33192 19304
rect 33140 19261 33149 19295
rect 33149 19261 33183 19295
rect 33183 19261 33192 19295
rect 33140 19252 33192 19261
rect 33324 19295 33376 19304
rect 33324 19261 33333 19295
rect 33333 19261 33367 19295
rect 33367 19261 33376 19295
rect 33324 19252 33376 19261
rect 1492 19159 1544 19168
rect 1492 19125 1501 19159
rect 1501 19125 1535 19159
rect 1535 19125 1544 19159
rect 1492 19116 1544 19125
rect 1952 19116 2004 19168
rect 34244 19329 34253 19363
rect 34253 19329 34287 19363
rect 34287 19329 34296 19363
rect 34244 19320 34296 19329
rect 12532 19159 12584 19168
rect 12532 19125 12541 19159
rect 12541 19125 12575 19159
rect 12575 19125 12584 19159
rect 12532 19116 12584 19125
rect 21916 19159 21968 19168
rect 21916 19125 21925 19159
rect 21925 19125 21959 19159
rect 21959 19125 21968 19159
rect 21916 19116 21968 19125
rect 23756 19159 23808 19168
rect 23756 19125 23765 19159
rect 23765 19125 23799 19159
rect 23799 19125 23808 19159
rect 23756 19116 23808 19125
rect 35348 19116 35400 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 33140 18912 33192 18964
rect 10416 18776 10468 18828
rect 12532 18708 12584 18760
rect 21916 18776 21968 18828
rect 35348 18708 35400 18760
rect 1492 18615 1544 18624
rect 1492 18581 1501 18615
rect 1501 18581 1535 18615
rect 1535 18581 1544 18615
rect 1492 18572 1544 18581
rect 9128 18572 9180 18624
rect 26056 18572 26108 18624
rect 33324 18572 33376 18624
rect 38016 18615 38068 18624
rect 38016 18581 38025 18615
rect 38025 18581 38059 18615
rect 38059 18581 38068 18615
rect 38016 18572 38068 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 14280 18411 14332 18420
rect 14280 18377 14289 18411
rect 14289 18377 14323 18411
rect 14323 18377 14332 18411
rect 14280 18368 14332 18377
rect 22468 18368 22520 18420
rect 22652 18300 22704 18352
rect 12992 18275 13044 18284
rect 12992 18241 13001 18275
rect 13001 18241 13035 18275
rect 13035 18241 13044 18275
rect 12992 18232 13044 18241
rect 24584 18096 24636 18148
rect 38108 18275 38160 18284
rect 38108 18241 38117 18275
rect 38117 18241 38151 18275
rect 38151 18241 38160 18275
rect 38108 18232 38160 18241
rect 33784 18096 33836 18148
rect 1492 18071 1544 18080
rect 1492 18037 1501 18071
rect 1501 18037 1535 18071
rect 1535 18037 1544 18071
rect 1492 18028 1544 18037
rect 26516 18028 26568 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 3516 17824 3568 17876
rect 12992 17756 13044 17808
rect 4620 17688 4672 17740
rect 8024 17620 8076 17672
rect 21824 17620 21876 17672
rect 26516 17663 26568 17672
rect 26516 17629 26525 17663
rect 26525 17629 26559 17663
rect 26559 17629 26568 17663
rect 26516 17620 26568 17629
rect 38108 17663 38160 17672
rect 38108 17629 38117 17663
rect 38117 17629 38151 17663
rect 38151 17629 38160 17663
rect 38108 17620 38160 17629
rect 1584 17484 1636 17536
rect 4896 17484 4948 17536
rect 10324 17484 10376 17536
rect 33876 17484 33928 17536
rect 37280 17527 37332 17536
rect 37280 17493 37289 17527
rect 37289 17493 37323 17527
rect 37323 17493 37332 17527
rect 37280 17484 37332 17493
rect 37648 17484 37700 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 1584 17323 1636 17332
rect 1584 17289 1593 17323
rect 1593 17289 1627 17323
rect 1627 17289 1636 17323
rect 1584 17280 1636 17289
rect 4620 17323 4672 17332
rect 4620 17289 4629 17323
rect 4629 17289 4663 17323
rect 4663 17289 4672 17323
rect 4620 17280 4672 17289
rect 21180 17280 21232 17332
rect 35808 17280 35860 17332
rect 37648 17323 37700 17332
rect 37648 17289 37657 17323
rect 37657 17289 37691 17323
rect 37691 17289 37700 17323
rect 37648 17280 37700 17289
rect 37740 17323 37792 17332
rect 37740 17289 37749 17323
rect 37749 17289 37783 17323
rect 37783 17289 37792 17323
rect 37740 17280 37792 17289
rect 21272 17212 21324 17264
rect 1400 17187 1452 17196
rect 1400 17153 1409 17187
rect 1409 17153 1443 17187
rect 1443 17153 1452 17187
rect 1400 17144 1452 17153
rect 37648 17144 37700 17196
rect 26976 17076 27028 17128
rect 37280 17076 37332 17128
rect 1952 16940 2004 16992
rect 8208 16940 8260 16992
rect 38016 16940 38068 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 18052 16668 18104 16720
rect 4068 16600 4120 16652
rect 2044 16532 2096 16584
rect 26148 16532 26200 16584
rect 26332 16396 26384 16448
rect 37188 16532 37240 16584
rect 38016 16575 38068 16584
rect 38016 16541 38025 16575
rect 38025 16541 38059 16575
rect 38059 16541 38068 16575
rect 38016 16532 38068 16541
rect 27068 16439 27120 16448
rect 27068 16405 27077 16439
rect 27077 16405 27111 16439
rect 27111 16405 27120 16439
rect 27068 16396 27120 16405
rect 35440 16396 35492 16448
rect 37740 16396 37792 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 2044 16235 2096 16244
rect 2044 16201 2053 16235
rect 2053 16201 2087 16235
rect 2087 16201 2096 16235
rect 2044 16192 2096 16201
rect 13820 16192 13872 16244
rect 21640 16192 21692 16244
rect 26148 16192 26200 16244
rect 37372 16235 37424 16244
rect 37372 16201 37381 16235
rect 37381 16201 37415 16235
rect 37415 16201 37424 16235
rect 37372 16192 37424 16201
rect 1400 16099 1452 16108
rect 1400 16065 1409 16099
rect 1409 16065 1443 16099
rect 1443 16065 1452 16099
rect 1400 16056 1452 16065
rect 1768 15852 1820 15904
rect 15476 15895 15528 15904
rect 15476 15861 15485 15895
rect 15485 15861 15519 15895
rect 15519 15861 15528 15895
rect 15476 15852 15528 15861
rect 27068 15988 27120 16040
rect 38476 15988 38528 16040
rect 21732 15852 21784 15904
rect 38016 15895 38068 15904
rect 38016 15861 38025 15895
rect 38025 15861 38059 15895
rect 38059 15861 38068 15895
rect 38016 15852 38068 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 1400 15691 1452 15700
rect 1400 15657 1409 15691
rect 1409 15657 1443 15691
rect 1443 15657 1452 15691
rect 1400 15648 1452 15657
rect 15476 15555 15528 15564
rect 15476 15521 15485 15555
rect 15485 15521 15519 15555
rect 15519 15521 15528 15555
rect 15476 15512 15528 15521
rect 16304 15444 16356 15496
rect 38108 15487 38160 15496
rect 38108 15453 38117 15487
rect 38117 15453 38151 15487
rect 38151 15453 38160 15487
rect 38108 15444 38160 15453
rect 26332 15308 26384 15360
rect 26976 15308 27028 15360
rect 37924 15351 37976 15360
rect 37924 15317 37933 15351
rect 37933 15317 37967 15351
rect 37967 15317 37976 15351
rect 37924 15308 37976 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 1768 15104 1820 15156
rect 4804 15104 4856 15156
rect 27068 15104 27120 15156
rect 4804 15011 4856 15020
rect 4804 14977 4813 15011
rect 4813 14977 4847 15011
rect 4847 14977 4856 15011
rect 4804 14968 4856 14977
rect 38016 15104 38068 15156
rect 37924 15036 37976 15088
rect 34612 15011 34664 15020
rect 28356 14943 28408 14952
rect 28356 14909 28365 14943
rect 28365 14909 28399 14943
rect 28399 14909 28408 14943
rect 28356 14900 28408 14909
rect 34612 14977 34621 15011
rect 34621 14977 34655 15011
rect 34655 14977 34664 15011
rect 34612 14968 34664 14977
rect 38568 14832 38620 14884
rect 27896 14807 27948 14816
rect 27896 14773 27905 14807
rect 27905 14773 27939 14807
rect 27939 14773 27948 14807
rect 27896 14764 27948 14773
rect 38108 14807 38160 14816
rect 38108 14773 38117 14807
rect 38117 14773 38151 14807
rect 38151 14773 38160 14807
rect 38108 14764 38160 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 26700 14560 26752 14612
rect 27896 14424 27948 14476
rect 37832 14467 37884 14476
rect 37832 14433 37841 14467
rect 37841 14433 37875 14467
rect 37875 14433 37884 14467
rect 37832 14424 37884 14433
rect 18972 14356 19024 14408
rect 27620 14399 27672 14408
rect 27620 14365 27629 14399
rect 27629 14365 27663 14399
rect 27663 14365 27672 14399
rect 27620 14356 27672 14365
rect 38108 14399 38160 14408
rect 38108 14365 38117 14399
rect 38117 14365 38151 14399
rect 38151 14365 38160 14399
rect 38108 14356 38160 14365
rect 1492 14263 1544 14272
rect 1492 14229 1501 14263
rect 1501 14229 1535 14263
rect 1535 14229 1544 14263
rect 1492 14220 1544 14229
rect 24124 14220 24176 14272
rect 26424 14220 26476 14272
rect 34428 14220 34480 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 24124 14016 24176 14068
rect 9220 13948 9272 14000
rect 14464 13948 14516 14000
rect 4620 13923 4672 13932
rect 2044 13812 2096 13864
rect 4620 13889 4629 13923
rect 4629 13889 4663 13923
rect 4663 13889 4672 13923
rect 4620 13880 4672 13889
rect 34520 14016 34572 14068
rect 26424 13948 26476 14000
rect 38292 13948 38344 14000
rect 14464 13812 14516 13864
rect 36820 13880 36872 13932
rect 27436 13855 27488 13864
rect 27436 13821 27445 13855
rect 27445 13821 27479 13855
rect 27479 13821 27488 13855
rect 27436 13812 27488 13821
rect 34428 13855 34480 13864
rect 26240 13744 26292 13796
rect 26700 13744 26752 13796
rect 34428 13821 34437 13855
rect 34437 13821 34471 13855
rect 34471 13821 34480 13855
rect 34428 13812 34480 13821
rect 26884 13676 26936 13728
rect 33968 13676 34020 13728
rect 38016 13719 38068 13728
rect 38016 13685 38025 13719
rect 38025 13685 38059 13719
rect 38059 13685 38068 13719
rect 38016 13676 38068 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 2044 13515 2096 13524
rect 2044 13481 2053 13515
rect 2053 13481 2087 13515
rect 2087 13481 2096 13515
rect 2044 13472 2096 13481
rect 4620 13472 4672 13524
rect 34612 13472 34664 13524
rect 4712 13336 4764 13388
rect 7472 13336 7524 13388
rect 34428 13336 34480 13388
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 5080 13268 5132 13320
rect 26884 13311 26936 13320
rect 26884 13277 26893 13311
rect 26893 13277 26927 13311
rect 26927 13277 26936 13311
rect 26884 13268 26936 13277
rect 33968 13311 34020 13320
rect 33968 13277 33977 13311
rect 33977 13277 34011 13311
rect 34011 13277 34020 13311
rect 33968 13268 34020 13277
rect 4712 13132 4764 13184
rect 35072 13268 35124 13320
rect 34980 13200 35032 13252
rect 35348 13268 35400 13320
rect 36820 13268 36872 13320
rect 37924 13200 37976 13252
rect 34612 13132 34664 13184
rect 35348 13132 35400 13184
rect 37832 13132 37884 13184
rect 38016 13175 38068 13184
rect 38016 13141 38025 13175
rect 38025 13141 38059 13175
rect 38059 13141 38068 13175
rect 38016 13132 38068 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 12992 12903 13044 12912
rect 12992 12869 13001 12903
rect 13001 12869 13035 12903
rect 13035 12869 13044 12903
rect 12992 12860 13044 12869
rect 10600 12792 10652 12844
rect 37648 12792 37700 12844
rect 38108 12767 38160 12776
rect 38108 12733 38117 12767
rect 38117 12733 38151 12767
rect 38151 12733 38160 12767
rect 38108 12724 38160 12733
rect 1492 12631 1544 12640
rect 1492 12597 1501 12631
rect 1501 12597 1535 12631
rect 1535 12597 1544 12631
rect 1492 12588 1544 12597
rect 13912 12588 13964 12640
rect 34428 12588 34480 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 10600 12427 10652 12436
rect 10600 12393 10609 12427
rect 10609 12393 10643 12427
rect 10643 12393 10652 12427
rect 10600 12384 10652 12393
rect 14648 12384 14700 12436
rect 20168 12384 20220 12436
rect 34428 12384 34480 12436
rect 38108 12359 38160 12368
rect 38108 12325 38117 12359
rect 38117 12325 38151 12359
rect 38151 12325 38160 12359
rect 38108 12316 38160 12325
rect 11796 12291 11848 12300
rect 11796 12257 11805 12291
rect 11805 12257 11839 12291
rect 11839 12257 11848 12291
rect 11796 12248 11848 12257
rect 1492 12087 1544 12096
rect 1492 12053 1501 12087
rect 1501 12053 1535 12087
rect 1535 12053 1544 12087
rect 1492 12044 1544 12053
rect 11612 12087 11664 12096
rect 11612 12053 11621 12087
rect 11621 12053 11655 12087
rect 11655 12053 11664 12087
rect 11612 12044 11664 12053
rect 17776 12044 17828 12096
rect 37280 12044 37332 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 3976 11840 4028 11892
rect 4804 11840 4856 11892
rect 22100 11840 22152 11892
rect 29736 11840 29788 11892
rect 8300 11772 8352 11824
rect 11796 11772 11848 11824
rect 14648 11772 14700 11824
rect 26792 11772 26844 11824
rect 37096 11772 37148 11824
rect 1492 11747 1544 11756
rect 1492 11713 1501 11747
rect 1501 11713 1535 11747
rect 1535 11713 1544 11747
rect 1492 11704 1544 11713
rect 1860 11704 1912 11756
rect 4620 11704 4672 11756
rect 14832 11747 14884 11756
rect 14832 11713 14841 11747
rect 14841 11713 14875 11747
rect 14875 11713 14884 11747
rect 14832 11704 14884 11713
rect 23480 11704 23532 11756
rect 37648 11704 37700 11756
rect 11612 11636 11664 11688
rect 15016 11636 15068 11688
rect 37280 11679 37332 11688
rect 37280 11645 37289 11679
rect 37289 11645 37323 11679
rect 37323 11645 37332 11679
rect 37280 11636 37332 11645
rect 9772 11568 9824 11620
rect 20996 11568 21048 11620
rect 29828 11568 29880 11620
rect 4712 11500 4764 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 1676 11296 1728 11348
rect 37924 11339 37976 11348
rect 37924 11305 37933 11339
rect 37933 11305 37967 11339
rect 37967 11305 37976 11339
rect 37924 11296 37976 11305
rect 1400 11135 1452 11144
rect 1400 11101 1409 11135
rect 1409 11101 1443 11135
rect 1443 11101 1452 11135
rect 1400 11092 1452 11101
rect 38108 11135 38160 11144
rect 38108 11101 38117 11135
rect 38117 11101 38151 11135
rect 38151 11101 38160 11135
rect 38108 11092 38160 11101
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 2412 10752 2464 10804
rect 8300 10795 8352 10804
rect 8300 10761 8309 10795
rect 8309 10761 8343 10795
rect 8343 10761 8352 10795
rect 8300 10752 8352 10761
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 6184 10616 6236 10668
rect 14740 10659 14792 10668
rect 14740 10625 14749 10659
rect 14749 10625 14783 10659
rect 14783 10625 14792 10659
rect 14740 10616 14792 10625
rect 38108 10659 38160 10668
rect 38108 10625 38117 10659
rect 38117 10625 38151 10659
rect 38151 10625 38160 10659
rect 38108 10616 38160 10625
rect 8300 10548 8352 10600
rect 14556 10591 14608 10600
rect 14556 10557 14565 10591
rect 14565 10557 14599 10591
rect 14599 10557 14608 10591
rect 14556 10548 14608 10557
rect 2504 10480 2556 10532
rect 23388 10480 23440 10532
rect 37280 10548 37332 10600
rect 1584 10455 1636 10464
rect 1584 10421 1593 10455
rect 1593 10421 1627 10455
rect 1627 10421 1636 10455
rect 1584 10412 1636 10421
rect 12164 10412 12216 10464
rect 15108 10455 15160 10464
rect 15108 10421 15117 10455
rect 15117 10421 15151 10455
rect 15151 10421 15160 10455
rect 15108 10412 15160 10421
rect 23756 10412 23808 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 1584 10208 1636 10260
rect 14740 10208 14792 10260
rect 37556 10208 37608 10260
rect 17224 10140 17276 10192
rect 1400 10047 1452 10056
rect 1400 10013 1409 10047
rect 1409 10013 1443 10047
rect 1443 10013 1452 10047
rect 1400 10004 1452 10013
rect 12164 10047 12216 10056
rect 12164 10013 12173 10047
rect 12173 10013 12207 10047
rect 12207 10013 12216 10047
rect 12164 10004 12216 10013
rect 15108 10004 15160 10056
rect 38108 10047 38160 10056
rect 38108 10013 38117 10047
rect 38117 10013 38151 10047
rect 38151 10013 38160 10047
rect 38108 10004 38160 10013
rect 14924 9936 14976 9988
rect 18144 9868 18196 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 14648 9596 14700 9648
rect 15476 9571 15528 9580
rect 15476 9537 15485 9571
rect 15485 9537 15519 9571
rect 15519 9537 15528 9571
rect 15476 9528 15528 9537
rect 14648 9503 14700 9512
rect 14648 9469 14657 9503
rect 14657 9469 14691 9503
rect 14691 9469 14700 9503
rect 14648 9460 14700 9469
rect 15016 9392 15068 9444
rect 30932 9324 30984 9376
rect 38108 9367 38160 9376
rect 38108 9333 38117 9367
rect 38117 9333 38151 9367
rect 38151 9333 38160 9367
rect 38108 9324 38160 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 33784 8984 33836 9036
rect 38108 8959 38160 8968
rect 38108 8925 38117 8959
rect 38117 8925 38151 8959
rect 38151 8925 38160 8959
rect 38108 8916 38160 8925
rect 19340 8848 19392 8900
rect 1492 8823 1544 8832
rect 1492 8789 1501 8823
rect 1501 8789 1535 8823
rect 1535 8789 1544 8823
rect 1492 8780 1544 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 14924 8576 14976 8628
rect 3700 8440 3752 8492
rect 15936 8440 15988 8492
rect 16304 8440 16356 8492
rect 2228 8415 2280 8424
rect 2228 8381 2237 8415
rect 2237 8381 2271 8415
rect 2271 8381 2280 8415
rect 2228 8372 2280 8381
rect 17960 8304 18012 8356
rect 38016 8347 38068 8356
rect 38016 8313 38025 8347
rect 38025 8313 38059 8347
rect 38059 8313 38068 8347
rect 38016 8304 38068 8313
rect 16120 8279 16172 8288
rect 16120 8245 16129 8279
rect 16129 8245 16163 8279
rect 16163 8245 16172 8279
rect 16120 8236 16172 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 13820 7896 13872 7948
rect 16120 7896 16172 7948
rect 2044 7828 2096 7880
rect 31024 7828 31076 7880
rect 36176 7760 36228 7812
rect 38016 7735 38068 7744
rect 38016 7701 38025 7735
rect 38025 7701 38059 7735
rect 38059 7701 38068 7735
rect 38016 7692 38068 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 2044 7531 2096 7540
rect 2044 7497 2053 7531
rect 2053 7497 2087 7531
rect 2087 7497 2096 7531
rect 2044 7488 2096 7497
rect 1400 7395 1452 7404
rect 1400 7361 1409 7395
rect 1409 7361 1443 7395
rect 1443 7361 1452 7395
rect 1400 7352 1452 7361
rect 22560 7395 22612 7404
rect 22560 7361 22569 7395
rect 22569 7361 22603 7395
rect 22603 7361 22612 7395
rect 22560 7352 22612 7361
rect 38016 7395 38068 7404
rect 38016 7361 38025 7395
rect 38025 7361 38059 7395
rect 38059 7361 38068 7395
rect 38016 7352 38068 7361
rect 4896 7284 4948 7336
rect 4620 7216 4672 7268
rect 31024 7216 31076 7268
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 1400 6919 1452 6928
rect 1400 6885 1409 6919
rect 1409 6885 1443 6919
rect 1443 6885 1452 6919
rect 1400 6876 1452 6885
rect 10692 6808 10744 6860
rect 12164 6808 12216 6860
rect 17960 6808 18012 6860
rect 22560 6808 22612 6860
rect 21732 6783 21784 6792
rect 21732 6749 21741 6783
rect 21741 6749 21775 6783
rect 21775 6749 21784 6783
rect 21732 6740 21784 6749
rect 11520 6672 11572 6724
rect 21548 6715 21600 6724
rect 21548 6681 21557 6715
rect 21557 6681 21591 6715
rect 21591 6681 21600 6715
rect 21548 6672 21600 6681
rect 30472 6604 30524 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 11520 6443 11572 6452
rect 11520 6409 11529 6443
rect 11529 6409 11563 6443
rect 11563 6409 11572 6443
rect 11520 6400 11572 6409
rect 17960 6400 18012 6452
rect 24952 6400 25004 6452
rect 37280 6443 37332 6452
rect 37280 6409 37289 6443
rect 37289 6409 37323 6443
rect 37323 6409 37332 6443
rect 37280 6400 37332 6409
rect 2320 6332 2372 6384
rect 20720 6332 20772 6384
rect 1768 6264 1820 6316
rect 1492 6171 1544 6180
rect 1492 6137 1501 6171
rect 1501 6137 1535 6171
rect 1535 6137 1544 6171
rect 1492 6128 1544 6137
rect 11980 6239 12032 6248
rect 11980 6205 11989 6239
rect 11989 6205 12023 6239
rect 12023 6205 12032 6239
rect 12164 6239 12216 6248
rect 11980 6196 12032 6205
rect 12164 6205 12173 6239
rect 12173 6205 12207 6239
rect 12207 6205 12216 6239
rect 12164 6196 12216 6205
rect 12256 6196 12308 6248
rect 14556 6196 14608 6248
rect 38384 6196 38436 6248
rect 38016 6171 38068 6180
rect 38016 6137 38025 6171
rect 38025 6137 38059 6171
rect 38059 6137 38068 6171
rect 38016 6128 38068 6137
rect 12808 6103 12860 6112
rect 12808 6069 12817 6103
rect 12817 6069 12851 6103
rect 12851 6069 12860 6103
rect 12808 6060 12860 6069
rect 12992 6060 13044 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 14556 5856 14608 5908
rect 17316 5856 17368 5908
rect 25412 5856 25464 5908
rect 4620 5788 4672 5840
rect 6368 5695 6420 5704
rect 6368 5661 6377 5695
rect 6377 5661 6411 5695
rect 6411 5661 6420 5695
rect 6368 5652 6420 5661
rect 8484 5584 8536 5636
rect 27620 5788 27672 5840
rect 12808 5720 12860 5772
rect 24952 5763 25004 5772
rect 12992 5695 13044 5704
rect 12992 5661 13001 5695
rect 13001 5661 13035 5695
rect 13035 5661 13044 5695
rect 12992 5652 13044 5661
rect 24952 5729 24961 5763
rect 24961 5729 24995 5763
rect 24995 5729 25004 5763
rect 24952 5720 25004 5729
rect 26332 5720 26384 5772
rect 26700 5652 26752 5704
rect 27620 5652 27672 5704
rect 37832 5695 37884 5704
rect 37832 5661 37841 5695
rect 37841 5661 37875 5695
rect 37875 5661 37884 5695
rect 37832 5652 37884 5661
rect 1492 5559 1544 5568
rect 1492 5525 1501 5559
rect 1501 5525 1535 5559
rect 1535 5525 1544 5559
rect 1492 5516 1544 5525
rect 2964 5516 3016 5568
rect 5816 5516 5868 5568
rect 9588 5516 9640 5568
rect 23756 5559 23808 5568
rect 23756 5525 23765 5559
rect 23765 5525 23799 5559
rect 23799 5525 23808 5559
rect 23756 5516 23808 5525
rect 24400 5559 24452 5568
rect 24400 5525 24409 5559
rect 24409 5525 24443 5559
rect 24443 5525 24452 5559
rect 24400 5516 24452 5525
rect 25412 5584 25464 5636
rect 38200 5584 38252 5636
rect 27068 5516 27120 5568
rect 37372 5559 37424 5568
rect 37372 5525 37381 5559
rect 37381 5525 37415 5559
rect 37415 5525 37424 5559
rect 37372 5516 37424 5525
rect 38016 5559 38068 5568
rect 38016 5525 38025 5559
rect 38025 5525 38059 5559
rect 38059 5525 38068 5559
rect 38016 5516 38068 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 6184 5312 6236 5364
rect 26332 5355 26384 5364
rect 26332 5321 26341 5355
rect 26341 5321 26375 5355
rect 26375 5321 26384 5355
rect 26332 5312 26384 5321
rect 37832 5312 37884 5364
rect 38476 5312 38528 5364
rect 1400 5219 1452 5228
rect 1400 5185 1409 5219
rect 1409 5185 1443 5219
rect 1443 5185 1452 5219
rect 1400 5176 1452 5185
rect 5816 5219 5868 5228
rect 5816 5185 5825 5219
rect 5825 5185 5859 5219
rect 5859 5185 5868 5219
rect 5816 5176 5868 5185
rect 24400 5176 24452 5228
rect 27068 5219 27120 5228
rect 27068 5185 27077 5219
rect 27077 5185 27111 5219
rect 27111 5185 27120 5219
rect 27068 5176 27120 5185
rect 37740 5176 37792 5228
rect 1676 4972 1728 5024
rect 2872 4972 2924 5024
rect 4804 4972 4856 5024
rect 25596 4972 25648 5024
rect 28908 4972 28960 5024
rect 36636 5015 36688 5024
rect 36636 4981 36645 5015
rect 36645 4981 36679 5015
rect 36679 4981 36688 5015
rect 36636 4972 36688 4981
rect 38016 5015 38068 5024
rect 38016 4981 38025 5015
rect 38025 4981 38059 5015
rect 38059 4981 38068 5015
rect 38016 4972 38068 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 2136 4811 2188 4820
rect 2136 4777 2145 4811
rect 2145 4777 2179 4811
rect 2179 4777 2188 4811
rect 2136 4768 2188 4777
rect 36176 4811 36228 4820
rect 36176 4777 36185 4811
rect 36185 4777 36219 4811
rect 36219 4777 36228 4811
rect 36176 4768 36228 4777
rect 37648 4700 37700 4752
rect 2136 4564 2188 4616
rect 17960 4564 18012 4616
rect 38016 4539 38068 4548
rect 38016 4505 38025 4539
rect 38025 4505 38059 4539
rect 38059 4505 38068 4539
rect 38016 4496 38068 4505
rect 1492 4471 1544 4480
rect 1492 4437 1501 4471
rect 1501 4437 1535 4471
rect 1535 4437 1544 4471
rect 1492 4428 1544 4437
rect 2780 4471 2832 4480
rect 2780 4437 2789 4471
rect 2789 4437 2823 4471
rect 2823 4437 2832 4471
rect 2780 4428 2832 4437
rect 3884 4471 3936 4480
rect 3884 4437 3893 4471
rect 3893 4437 3927 4471
rect 3927 4437 3936 4471
rect 3884 4428 3936 4437
rect 15568 4471 15620 4480
rect 15568 4437 15577 4471
rect 15577 4437 15611 4471
rect 15611 4437 15620 4471
rect 15568 4428 15620 4437
rect 34796 4428 34848 4480
rect 35716 4471 35768 4480
rect 35716 4437 35725 4471
rect 35725 4437 35759 4471
rect 35759 4437 35768 4471
rect 35716 4428 35768 4437
rect 36728 4471 36780 4480
rect 36728 4437 36737 4471
rect 36737 4437 36771 4471
rect 36771 4437 36780 4471
rect 36728 4428 36780 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 37372 4156 37424 4208
rect 39304 4156 39356 4208
rect 664 4088 716 4140
rect 1676 4088 1728 4140
rect 2780 4088 2832 4140
rect 3332 4088 3384 4140
rect 10324 4088 10376 4140
rect 13452 4088 13504 4140
rect 18052 4088 18104 4140
rect 24676 4088 24728 4140
rect 26240 4088 26292 4140
rect 30840 4131 30892 4140
rect 30840 4097 30849 4131
rect 30849 4097 30883 4131
rect 30883 4097 30892 4131
rect 30840 4088 30892 4097
rect 37096 4088 37148 4140
rect 9680 3952 9732 4004
rect 15292 4020 15344 4072
rect 17500 3952 17552 4004
rect 25228 3952 25280 4004
rect 2688 3927 2740 3936
rect 2688 3893 2697 3927
rect 2697 3893 2731 3927
rect 2731 3893 2740 3927
rect 2688 3884 2740 3893
rect 3700 3927 3752 3936
rect 3700 3893 3709 3927
rect 3709 3893 3743 3927
rect 3743 3893 3752 3927
rect 3700 3884 3752 3893
rect 4068 3884 4120 3936
rect 4712 3927 4764 3936
rect 4712 3893 4721 3927
rect 4721 3893 4755 3927
rect 4755 3893 4764 3927
rect 4712 3884 4764 3893
rect 16120 3927 16172 3936
rect 16120 3893 16129 3927
rect 16129 3893 16163 3927
rect 16163 3893 16172 3927
rect 16120 3884 16172 3893
rect 35440 3927 35492 3936
rect 35440 3893 35449 3927
rect 35449 3893 35483 3927
rect 35483 3893 35492 3927
rect 35440 3884 35492 3893
rect 36084 3927 36136 3936
rect 36084 3893 36093 3927
rect 36093 3893 36127 3927
rect 36127 3893 36136 3927
rect 36084 3884 36136 3893
rect 36452 3884 36504 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 3976 3723 4028 3732
rect 3976 3689 3985 3723
rect 3985 3689 4019 3723
rect 4019 3689 4028 3723
rect 3976 3680 4028 3689
rect 5632 3723 5684 3732
rect 5632 3689 5641 3723
rect 5641 3689 5675 3723
rect 5675 3689 5684 3723
rect 5632 3680 5684 3689
rect 13452 3723 13504 3732
rect 13452 3689 13461 3723
rect 13461 3689 13495 3723
rect 13495 3689 13504 3723
rect 13452 3680 13504 3689
rect 14464 3680 14516 3732
rect 17960 3723 18012 3732
rect 4620 3612 4672 3664
rect 17960 3689 17969 3723
rect 17969 3689 18003 3723
rect 18003 3689 18012 3723
rect 17960 3680 18012 3689
rect 18052 3680 18104 3732
rect 26608 3680 26660 3732
rect 30472 3723 30524 3732
rect 30472 3689 30481 3723
rect 30481 3689 30515 3723
rect 30515 3689 30524 3723
rect 30472 3680 30524 3689
rect 31024 3723 31076 3732
rect 31024 3689 31033 3723
rect 31033 3689 31067 3723
rect 31067 3689 31076 3723
rect 31024 3680 31076 3689
rect 33876 3723 33928 3732
rect 33876 3689 33885 3723
rect 33885 3689 33919 3723
rect 33919 3689 33928 3723
rect 33876 3680 33928 3689
rect 1952 3587 2004 3596
rect 1952 3553 1961 3587
rect 1961 3553 1995 3587
rect 1995 3553 2004 3587
rect 1952 3544 2004 3553
rect 2228 3587 2280 3596
rect 2228 3553 2237 3587
rect 2237 3553 2271 3587
rect 2271 3553 2280 3587
rect 2228 3544 2280 3553
rect 4712 3544 4764 3596
rect 13912 3544 13964 3596
rect 17316 3587 17368 3596
rect 17316 3553 17325 3587
rect 17325 3553 17359 3587
rect 17359 3553 17368 3587
rect 17316 3544 17368 3553
rect 17500 3587 17552 3596
rect 17500 3553 17509 3587
rect 17509 3553 17543 3587
rect 17543 3553 17552 3587
rect 17500 3544 17552 3553
rect 18420 3612 18472 3664
rect 24676 3612 24728 3664
rect 33324 3612 33376 3664
rect 38660 3612 38712 3664
rect 22744 3544 22796 3596
rect 24768 3544 24820 3596
rect 36544 3544 36596 3596
rect 2688 3519 2740 3528
rect 2688 3485 2697 3519
rect 2697 3485 2731 3519
rect 2731 3485 2740 3519
rect 2688 3476 2740 3485
rect 3700 3476 3752 3528
rect 1952 3408 2004 3460
rect 2596 3408 2648 3460
rect 9496 3476 9548 3528
rect 14372 3476 14424 3528
rect 16120 3476 16172 3528
rect 4620 3340 4672 3392
rect 6184 3383 6236 3392
rect 6184 3349 6193 3383
rect 6193 3349 6227 3383
rect 6227 3349 6236 3383
rect 6184 3340 6236 3349
rect 11612 3383 11664 3392
rect 11612 3349 11621 3383
rect 11621 3349 11655 3383
rect 11655 3349 11664 3383
rect 11612 3340 11664 3349
rect 14924 3383 14976 3392
rect 14924 3349 14933 3383
rect 14933 3349 14967 3383
rect 14967 3349 14976 3383
rect 14924 3340 14976 3349
rect 27712 3476 27764 3528
rect 30932 3476 30984 3528
rect 36084 3476 36136 3528
rect 37096 3519 37148 3528
rect 17500 3408 17552 3460
rect 18420 3451 18472 3460
rect 18420 3417 18429 3451
rect 18429 3417 18463 3451
rect 18463 3417 18472 3451
rect 18420 3408 18472 3417
rect 25964 3408 26016 3460
rect 37096 3485 37105 3519
rect 37105 3485 37139 3519
rect 37139 3485 37148 3519
rect 37096 3476 37148 3485
rect 37832 3519 37884 3528
rect 37832 3485 37841 3519
rect 37841 3485 37875 3519
rect 37875 3485 37884 3519
rect 37832 3476 37884 3485
rect 17592 3383 17644 3392
rect 17592 3349 17601 3383
rect 17601 3349 17635 3383
rect 17635 3349 17644 3383
rect 17592 3340 17644 3349
rect 21088 3340 21140 3392
rect 23204 3383 23256 3392
rect 23204 3349 23213 3383
rect 23213 3349 23247 3383
rect 23247 3349 23256 3383
rect 23204 3340 23256 3349
rect 23664 3383 23716 3392
rect 23664 3349 23673 3383
rect 23673 3349 23707 3383
rect 23707 3349 23716 3383
rect 23664 3340 23716 3349
rect 24492 3340 24544 3392
rect 26424 3340 26476 3392
rect 27160 3340 27212 3392
rect 27528 3340 27580 3392
rect 28908 3340 28960 3392
rect 32036 3340 32088 3392
rect 32220 3383 32272 3392
rect 32220 3349 32229 3383
rect 32229 3349 32263 3383
rect 32263 3349 32272 3383
rect 32220 3340 32272 3349
rect 32772 3383 32824 3392
rect 32772 3349 32781 3383
rect 32781 3349 32815 3383
rect 32815 3349 32824 3383
rect 32772 3340 32824 3349
rect 32864 3340 32916 3392
rect 34152 3340 34204 3392
rect 36820 3340 36872 3392
rect 38016 3383 38068 3392
rect 38016 3349 38025 3383
rect 38025 3349 38059 3383
rect 38059 3349 38068 3383
rect 38016 3340 38068 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 2320 3179 2372 3188
rect 2320 3145 2329 3179
rect 2329 3145 2363 3179
rect 2363 3145 2372 3179
rect 2320 3136 2372 3145
rect 8484 3179 8536 3188
rect 8484 3145 8493 3179
rect 8493 3145 8527 3179
rect 8527 3145 8536 3179
rect 8484 3136 8536 3145
rect 9772 3179 9824 3188
rect 9772 3145 9781 3179
rect 9781 3145 9815 3179
rect 9815 3145 9824 3179
rect 9772 3136 9824 3145
rect 10416 3179 10468 3188
rect 10416 3145 10425 3179
rect 10425 3145 10459 3179
rect 10459 3145 10468 3179
rect 10416 3136 10468 3145
rect 12716 3136 12768 3188
rect 15292 3179 15344 3188
rect 20 3068 72 3120
rect 2872 3000 2924 3052
rect 3240 3068 3292 3120
rect 9496 3068 9548 3120
rect 9680 3068 9732 3120
rect 15292 3145 15301 3179
rect 15301 3145 15335 3179
rect 15335 3145 15344 3179
rect 15292 3136 15344 3145
rect 17592 3136 17644 3188
rect 17776 3136 17828 3188
rect 20536 3179 20588 3188
rect 20536 3145 20545 3179
rect 20545 3145 20579 3179
rect 20579 3145 20588 3179
rect 20536 3136 20588 3145
rect 25964 3179 26016 3188
rect 25964 3145 25973 3179
rect 25973 3145 26007 3179
rect 26007 3145 26016 3179
rect 25964 3136 26016 3145
rect 26976 3179 27028 3188
rect 26976 3145 26985 3179
rect 26985 3145 27019 3179
rect 27019 3145 27028 3179
rect 26976 3136 27028 3145
rect 27436 3136 27488 3188
rect 28356 3136 28408 3188
rect 4068 3000 4120 3052
rect 4620 3043 4672 3052
rect 4620 3009 4629 3043
rect 4629 3009 4663 3043
rect 4663 3009 4672 3043
rect 4620 3000 4672 3009
rect 5632 3000 5684 3052
rect 7104 3000 7156 3052
rect 8392 3000 8444 3052
rect 10968 3000 11020 3052
rect 12900 3000 12952 3052
rect 13912 3043 13964 3052
rect 13912 3009 13921 3043
rect 13921 3009 13955 3043
rect 13955 3009 13964 3043
rect 13912 3000 13964 3009
rect 14924 3000 14976 3052
rect 17408 3000 17460 3052
rect 18696 3000 18748 3052
rect 21088 3043 21140 3052
rect 21088 3009 21097 3043
rect 21097 3009 21131 3043
rect 21131 3009 21140 3043
rect 21088 3000 21140 3009
rect 24400 3000 24452 3052
rect 1308 2796 1360 2848
rect 12256 2932 12308 2984
rect 21456 2932 21508 2984
rect 11980 2864 12032 2916
rect 21548 2864 21600 2916
rect 23204 2932 23256 2984
rect 24676 2975 24728 2984
rect 24676 2941 24685 2975
rect 24685 2941 24719 2975
rect 24719 2941 24728 2975
rect 24676 2932 24728 2941
rect 5172 2796 5224 2848
rect 8392 2796 8444 2848
rect 9036 2796 9088 2848
rect 10968 2839 11020 2848
rect 10968 2805 10977 2839
rect 10977 2805 11011 2839
rect 11011 2805 11020 2839
rect 10968 2796 11020 2805
rect 16120 2796 16172 2848
rect 21916 2839 21968 2848
rect 21916 2805 21925 2839
rect 21925 2805 21959 2839
rect 21959 2805 21968 2839
rect 21916 2796 21968 2805
rect 22008 2796 22060 2848
rect 26424 3000 26476 3052
rect 27068 2932 27120 2984
rect 27528 2932 27580 2984
rect 28540 3000 28592 3052
rect 31668 3136 31720 3188
rect 34612 3136 34664 3188
rect 36544 3179 36596 3188
rect 36544 3145 36553 3179
rect 36553 3145 36587 3179
rect 36587 3145 36596 3179
rect 36544 3136 36596 3145
rect 32036 3068 32088 3120
rect 32312 3000 32364 3052
rect 32772 3000 32824 3052
rect 30472 2932 30524 2984
rect 27804 2796 27856 2848
rect 29644 2839 29696 2848
rect 29644 2805 29653 2839
rect 29653 2805 29687 2839
rect 29687 2805 29696 2839
rect 29644 2796 29696 2805
rect 32864 2932 32916 2984
rect 34152 3000 34204 3052
rect 35440 3000 35492 3052
rect 36176 3068 36228 3120
rect 36728 2932 36780 2984
rect 37924 2932 37976 2984
rect 34796 2864 34848 2916
rect 34520 2796 34572 2848
rect 35900 2839 35952 2848
rect 35900 2805 35909 2839
rect 35909 2805 35943 2839
rect 35943 2805 35952 2839
rect 35900 2796 35952 2805
rect 37372 2796 37424 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 8024 2635 8076 2644
rect 8024 2601 8033 2635
rect 8033 2601 8067 2635
rect 8067 2601 8076 2635
rect 8024 2592 8076 2601
rect 9128 2635 9180 2644
rect 9128 2601 9137 2635
rect 9137 2601 9171 2635
rect 9171 2601 9180 2635
rect 9128 2592 9180 2601
rect 15476 2635 15528 2644
rect 15476 2601 15485 2635
rect 15485 2601 15519 2635
rect 15519 2601 15528 2635
rect 15476 2592 15528 2601
rect 15936 2635 15988 2644
rect 15936 2601 15945 2635
rect 15945 2601 15979 2635
rect 15979 2601 15988 2635
rect 15936 2592 15988 2601
rect 23756 2592 23808 2644
rect 24400 2635 24452 2644
rect 24400 2601 24409 2635
rect 24409 2601 24443 2635
rect 24443 2601 24452 2635
rect 24400 2592 24452 2601
rect 26700 2592 26752 2644
rect 27620 2635 27672 2644
rect 27620 2601 27629 2635
rect 27629 2601 27663 2635
rect 27663 2601 27672 2635
rect 27620 2592 27672 2601
rect 27804 2592 27856 2644
rect 28448 2592 28500 2644
rect 34520 2592 34572 2644
rect 35808 2635 35860 2644
rect 35808 2601 35817 2635
rect 35817 2601 35851 2635
rect 35851 2601 35860 2635
rect 35808 2592 35860 2601
rect 3884 2456 3936 2508
rect 10508 2456 10560 2508
rect 18604 2524 18656 2576
rect 23848 2524 23900 2576
rect 17224 2456 17276 2508
rect 2964 2388 3016 2440
rect 4804 2388 4856 2440
rect 5816 2388 5868 2440
rect 6184 2388 6236 2440
rect 9588 2388 9640 2440
rect 9772 2388 9824 2440
rect 10416 2388 10468 2440
rect 11612 2388 11664 2440
rect 13268 2431 13320 2440
rect 13268 2397 13277 2431
rect 13277 2397 13311 2431
rect 13311 2397 13320 2431
rect 13268 2388 13320 2397
rect 14464 2388 14516 2440
rect 15568 2388 15620 2440
rect 16120 2431 16172 2440
rect 16120 2397 16129 2431
rect 16129 2397 16163 2431
rect 16163 2397 16172 2431
rect 16120 2388 16172 2397
rect 17684 2431 17736 2440
rect 17684 2397 17693 2431
rect 17693 2397 17727 2431
rect 17727 2397 17736 2431
rect 17684 2388 17736 2397
rect 18144 2431 18196 2440
rect 18144 2397 18153 2431
rect 18153 2397 18187 2431
rect 18187 2397 18196 2431
rect 18144 2388 18196 2397
rect 21916 2456 21968 2508
rect 22284 2499 22336 2508
rect 22284 2465 22293 2499
rect 22293 2465 22327 2499
rect 22327 2465 22336 2499
rect 22284 2456 22336 2465
rect 26148 2456 26200 2508
rect 20536 2388 20588 2440
rect 25596 2431 25648 2440
rect 7748 2320 7800 2372
rect 9036 2363 9088 2372
rect 9036 2329 9045 2363
rect 9045 2329 9079 2363
rect 9079 2329 9088 2363
rect 9036 2320 9088 2329
rect 3240 2252 3292 2304
rect 5724 2295 5776 2304
rect 5724 2261 5733 2295
rect 5733 2261 5767 2295
rect 5767 2261 5776 2295
rect 5724 2252 5776 2261
rect 6460 2252 6512 2304
rect 8760 2252 8812 2304
rect 9680 2252 9732 2304
rect 10324 2252 10376 2304
rect 12256 2252 12308 2304
rect 13544 2252 13596 2304
rect 16764 2252 16816 2304
rect 18052 2252 18104 2304
rect 19340 2252 19392 2304
rect 19984 2252 20036 2304
rect 20628 2252 20680 2304
rect 21916 2320 21968 2372
rect 25596 2397 25605 2431
rect 25605 2397 25639 2431
rect 25639 2397 25648 2431
rect 25596 2388 25648 2397
rect 27160 2431 27212 2440
rect 27160 2397 27169 2431
rect 27169 2397 27203 2431
rect 27203 2397 27212 2431
rect 27160 2388 27212 2397
rect 29736 2524 29788 2576
rect 27988 2456 28040 2508
rect 35716 2456 35768 2508
rect 37648 2456 37700 2508
rect 23664 2320 23716 2372
rect 24860 2295 24912 2304
rect 24860 2261 24869 2295
rect 24869 2261 24903 2295
rect 24903 2261 24912 2295
rect 24860 2252 24912 2261
rect 25780 2320 25832 2372
rect 27712 2320 27764 2372
rect 29644 2388 29696 2440
rect 30012 2431 30064 2440
rect 30012 2397 30021 2431
rect 30021 2397 30055 2431
rect 30055 2397 30064 2431
rect 30012 2388 30064 2397
rect 30840 2388 30892 2440
rect 31760 2388 31812 2440
rect 32220 2388 32272 2440
rect 33876 2431 33928 2440
rect 33876 2397 33885 2431
rect 33885 2397 33919 2431
rect 33919 2397 33928 2431
rect 33876 2388 33928 2397
rect 34796 2388 34848 2440
rect 36636 2431 36688 2440
rect 36636 2397 36645 2431
rect 36645 2397 36679 2431
rect 36679 2397 36688 2431
rect 36636 2388 36688 2397
rect 36452 2320 36504 2372
rect 28448 2252 28500 2304
rect 30288 2252 30340 2304
rect 33508 2252 33560 2304
rect 34796 2252 34848 2304
rect 35164 2252 35216 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 20076 2048 20128 2100
rect 30012 2048 30064 2100
rect 5724 1980 5776 2032
rect 24308 1980 24360 2032
rect 29920 1980 29972 2032
rect 35164 1980 35216 2032
rect 24860 1912 24912 1964
rect 31484 1912 31536 1964
rect 25136 1844 25188 1896
rect 27160 1844 27212 1896
rect 22560 1708 22612 1760
rect 23664 1708 23716 1760
<< metal2 >>
rect 18 49314 74 50000
rect 18 49286 152 49314
rect 18 49200 74 49286
rect 20 47456 72 47462
rect 20 47398 72 47404
rect 32 45558 60 47398
rect 20 45552 72 45558
rect 20 45494 72 45500
rect 124 45490 152 49286
rect 662 49200 718 50000
rect 1306 49314 1362 50000
rect 952 49286 1362 49314
rect 676 46714 704 49200
rect 952 47462 980 49286
rect 1306 49200 1362 49286
rect 1950 49314 2006 50000
rect 2594 49314 2650 50000
rect 2870 49736 2926 49745
rect 2926 49694 3004 49722
rect 2870 49671 2926 49680
rect 1950 49286 2084 49314
rect 1950 49200 2006 49286
rect 940 47456 992 47462
rect 940 47398 992 47404
rect 2056 47054 2084 49286
rect 2594 49286 2728 49314
rect 2594 49200 2650 49286
rect 2044 47048 2096 47054
rect 2044 46990 2096 46996
rect 2596 47048 2648 47054
rect 2596 46990 2648 46996
rect 664 46708 716 46714
rect 664 46650 716 46656
rect 2504 46436 2556 46442
rect 2504 46378 2556 46384
rect 2320 46368 2372 46374
rect 2320 46310 2372 46316
rect 2332 45966 2360 46310
rect 2320 45960 2372 45966
rect 2320 45902 2372 45908
rect 1492 45824 1544 45830
rect 1492 45766 1544 45772
rect 1504 45665 1532 45766
rect 1490 45656 1546 45665
rect 1490 45591 1546 45600
rect 112 45484 164 45490
rect 112 45426 164 45432
rect 1308 45484 1360 45490
rect 1308 45426 1360 45432
rect 1320 44470 1348 45426
rect 2412 45348 2464 45354
rect 2412 45290 2464 45296
rect 1952 44736 2004 44742
rect 1952 44678 2004 44684
rect 1308 44464 1360 44470
rect 1308 44406 1360 44412
rect 1400 44396 1452 44402
rect 1400 44338 1452 44344
rect 1412 44305 1440 44338
rect 1398 44296 1454 44305
rect 1398 44231 1454 44240
rect 1768 44192 1820 44198
rect 1768 44134 1820 44140
rect 1400 43784 1452 43790
rect 1400 43726 1452 43732
rect 1412 43625 1440 43726
rect 1398 43616 1454 43625
rect 1398 43551 1454 43560
rect 1400 43308 1452 43314
rect 1400 43250 1452 43256
rect 1412 42945 1440 43250
rect 1398 42936 1454 42945
rect 1398 42871 1454 42880
rect 1400 42696 1452 42702
rect 1400 42638 1452 42644
rect 1412 42265 1440 42638
rect 1398 42256 1454 42265
rect 1398 42191 1454 42200
rect 1400 39976 1452 39982
rect 1400 39918 1452 39924
rect 1584 39976 1636 39982
rect 1584 39918 1636 39924
rect 1412 39574 1440 39918
rect 1400 39568 1452 39574
rect 1398 39536 1400 39545
rect 1452 39536 1454 39545
rect 1398 39471 1454 39480
rect 1490 38856 1546 38865
rect 1490 38791 1492 38800
rect 1544 38791 1546 38800
rect 1492 38762 1544 38768
rect 1492 37120 1544 37126
rect 1492 37062 1544 37068
rect 1504 36825 1532 37062
rect 1490 36816 1546 36825
rect 1490 36751 1546 36760
rect 1490 36136 1546 36145
rect 1490 36071 1546 36080
rect 1504 36038 1532 36071
rect 1492 36032 1544 36038
rect 1492 35974 1544 35980
rect 1492 35488 1544 35494
rect 1490 35456 1492 35465
rect 1544 35456 1546 35465
rect 1490 35391 1546 35400
rect 1492 34944 1544 34950
rect 1492 34886 1544 34892
rect 1504 34785 1532 34886
rect 1490 34776 1546 34785
rect 1490 34711 1546 34720
rect 1400 33516 1452 33522
rect 1400 33458 1452 33464
rect 1412 33425 1440 33458
rect 1398 33416 1454 33425
rect 1398 33351 1454 33360
rect 1400 32904 1452 32910
rect 1400 32846 1452 32852
rect 1412 32745 1440 32846
rect 1398 32736 1454 32745
rect 1398 32671 1454 32680
rect 1492 32224 1544 32230
rect 1492 32166 1544 32172
rect 1504 32065 1532 32166
rect 1490 32056 1546 32065
rect 1490 31991 1546 32000
rect 1400 31816 1452 31822
rect 1400 31758 1452 31764
rect 1412 31385 1440 31758
rect 1398 31376 1454 31385
rect 1398 31311 1454 31320
rect 1412 30938 1440 31311
rect 1596 31142 1624 39918
rect 1676 36168 1728 36174
rect 1676 36110 1728 36116
rect 1688 35290 1716 36110
rect 1676 35284 1728 35290
rect 1676 35226 1728 35232
rect 1780 33998 1808 44134
rect 1860 42016 1912 42022
rect 1860 41958 1912 41964
rect 1872 41614 1900 41958
rect 1860 41608 1912 41614
rect 1858 41576 1860 41585
rect 1912 41576 1914 41585
rect 1858 41511 1914 41520
rect 1860 40452 1912 40458
rect 1860 40394 1912 40400
rect 1872 40225 1900 40394
rect 1858 40216 1914 40225
rect 1858 40151 1914 40160
rect 1964 39370 1992 44678
rect 2228 41064 2280 41070
rect 2228 41006 2280 41012
rect 2240 40905 2268 41006
rect 2226 40896 2282 40905
rect 2226 40831 2282 40840
rect 2044 40452 2096 40458
rect 2044 40394 2096 40400
rect 1952 39364 2004 39370
rect 1952 39306 2004 39312
rect 1768 33992 1820 33998
rect 1768 33934 1820 33940
rect 1676 33856 1728 33862
rect 1676 33798 1728 33804
rect 1584 31136 1636 31142
rect 1584 31078 1636 31084
rect 1400 30932 1452 30938
rect 1400 30874 1452 30880
rect 1492 30048 1544 30054
rect 1490 30016 1492 30025
rect 1544 30016 1546 30025
rect 1490 29951 1546 29960
rect 1492 29504 1544 29510
rect 1492 29446 1544 29452
rect 1504 29345 1532 29446
rect 1490 29336 1546 29345
rect 1490 29271 1546 29280
rect 1400 29164 1452 29170
rect 1400 29106 1452 29112
rect 1412 28665 1440 29106
rect 1398 28656 1454 28665
rect 1398 28591 1454 28600
rect 1400 28076 1452 28082
rect 1400 28018 1452 28024
rect 1412 27985 1440 28018
rect 1398 27976 1454 27985
rect 1398 27911 1454 27920
rect 1400 27464 1452 27470
rect 1400 27406 1452 27412
rect 1412 27305 1440 27406
rect 1398 27296 1454 27305
rect 1398 27231 1454 27240
rect 1492 26784 1544 26790
rect 1492 26726 1544 26732
rect 1504 26625 1532 26726
rect 1490 26616 1546 26625
rect 1490 26551 1546 26560
rect 1492 26240 1544 26246
rect 1492 26182 1544 26188
rect 1504 25945 1532 26182
rect 1490 25936 1546 25945
rect 1490 25871 1546 25880
rect 1400 24812 1452 24818
rect 1400 24754 1452 24760
rect 1412 24585 1440 24754
rect 1398 24576 1454 24585
rect 1398 24511 1454 24520
rect 1492 23520 1544 23526
rect 1492 23462 1544 23468
rect 1504 23225 1532 23462
rect 1490 23216 1546 23225
rect 1490 23151 1546 23160
rect 1400 22636 1452 22642
rect 1400 22578 1452 22584
rect 1412 22545 1440 22578
rect 1398 22536 1454 22545
rect 1398 22471 1454 22480
rect 1584 22432 1636 22438
rect 1584 22374 1636 22380
rect 1596 22234 1624 22374
rect 1584 22228 1636 22234
rect 1584 22170 1636 22176
rect 1400 22024 1452 22030
rect 1400 21966 1452 21972
rect 1412 21865 1440 21966
rect 1688 21894 1716 33798
rect 1860 31272 1912 31278
rect 1860 31214 1912 31220
rect 1768 31136 1820 31142
rect 1768 31078 1820 31084
rect 1676 21888 1728 21894
rect 1398 21856 1454 21865
rect 1676 21830 1728 21836
rect 1398 21791 1454 21800
rect 1400 20936 1452 20942
rect 1400 20878 1452 20884
rect 1412 20534 1440 20878
rect 1400 20528 1452 20534
rect 1398 20496 1400 20505
rect 1452 20496 1454 20505
rect 1398 20431 1454 20440
rect 1584 20460 1636 20466
rect 1584 20402 1636 20408
rect 1492 19168 1544 19174
rect 1490 19136 1492 19145
rect 1544 19136 1546 19145
rect 1490 19071 1546 19080
rect 1492 18624 1544 18630
rect 1492 18566 1544 18572
rect 1596 18578 1624 20402
rect 1676 19712 1728 19718
rect 1676 19654 1728 19660
rect 1688 19378 1716 19654
rect 1676 19372 1728 19378
rect 1676 19314 1728 19320
rect 1504 18465 1532 18566
rect 1596 18550 1716 18578
rect 1490 18456 1546 18465
rect 1490 18391 1546 18400
rect 1492 18080 1544 18086
rect 1492 18022 1544 18028
rect 1504 17785 1532 18022
rect 1490 17776 1546 17785
rect 1490 17711 1546 17720
rect 1584 17536 1636 17542
rect 1584 17478 1636 17484
rect 1596 17338 1624 17478
rect 1584 17332 1636 17338
rect 1584 17274 1636 17280
rect 1400 17196 1452 17202
rect 1400 17138 1452 17144
rect 1412 17105 1440 17138
rect 1398 17096 1454 17105
rect 1398 17031 1454 17040
rect 1400 16108 1452 16114
rect 1400 16050 1452 16056
rect 1412 15745 1440 16050
rect 1398 15736 1454 15745
rect 1398 15671 1400 15680
rect 1452 15671 1454 15680
rect 1400 15642 1452 15648
rect 1490 14376 1546 14385
rect 1490 14311 1546 14320
rect 1504 14278 1532 14311
rect 1492 14272 1544 14278
rect 1492 14214 1544 14220
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1412 13025 1440 13262
rect 1398 13016 1454 13025
rect 1398 12951 1454 12960
rect 1492 12640 1544 12646
rect 1492 12582 1544 12588
rect 1504 12345 1532 12582
rect 1490 12336 1546 12345
rect 1490 12271 1546 12280
rect 1492 12096 1544 12102
rect 1492 12038 1544 12044
rect 1504 11762 1532 12038
rect 1492 11756 1544 11762
rect 1492 11698 1544 11704
rect 1504 11665 1532 11698
rect 1490 11656 1546 11665
rect 1490 11591 1546 11600
rect 1688 11354 1716 18550
rect 1780 15910 1808 31078
rect 1872 27606 1900 31214
rect 1860 27600 1912 27606
rect 1860 27542 1912 27548
rect 2056 26234 2084 40394
rect 2228 38344 2280 38350
rect 2228 38286 2280 38292
rect 2240 38185 2268 38286
rect 2226 38176 2282 38185
rect 2226 38111 2282 38120
rect 2228 37800 2280 37806
rect 2228 37742 2280 37748
rect 2240 37505 2268 37742
rect 2226 37496 2282 37505
rect 2226 37431 2282 37440
rect 2136 37120 2188 37126
rect 2136 37062 2188 37068
rect 2148 31090 2176 37062
rect 2228 35488 2280 35494
rect 2228 35430 2280 35436
rect 2240 35154 2268 35430
rect 2228 35148 2280 35154
rect 2228 35090 2280 35096
rect 2320 35080 2372 35086
rect 2320 35022 2372 35028
rect 2228 34536 2280 34542
rect 2228 34478 2280 34484
rect 2240 34105 2268 34478
rect 2332 34202 2360 35022
rect 2320 34196 2372 34202
rect 2320 34138 2372 34144
rect 2226 34096 2282 34105
rect 2226 34031 2282 34040
rect 2148 31062 2268 31090
rect 2056 26206 2176 26234
rect 1860 25696 1912 25702
rect 1860 25638 1912 25644
rect 1872 25294 1900 25638
rect 1860 25288 1912 25294
rect 1858 25256 1860 25265
rect 1912 25256 1914 25265
rect 1858 25191 1914 25200
rect 2042 24168 2098 24177
rect 1860 24132 1912 24138
rect 2042 24103 2044 24112
rect 1860 24074 1912 24080
rect 2096 24103 2098 24112
rect 2044 24074 2096 24080
rect 1872 23905 1900 24074
rect 1858 23896 1914 23905
rect 1858 23831 1914 23840
rect 2044 21480 2096 21486
rect 2044 21422 2096 21428
rect 2056 21185 2084 21422
rect 2042 21176 2098 21185
rect 2042 21111 2044 21120
rect 2096 21111 2098 21120
rect 2044 21082 2096 21088
rect 2148 19938 2176 26206
rect 2240 24138 2268 31062
rect 2320 25696 2372 25702
rect 2320 25638 2372 25644
rect 2228 24132 2280 24138
rect 2228 24074 2280 24080
rect 2228 20256 2280 20262
rect 2228 20198 2280 20204
rect 1872 19910 2176 19938
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1768 15156 1820 15162
rect 1768 15098 1820 15104
rect 1676 11348 1728 11354
rect 1676 11290 1728 11296
rect 1400 11144 1452 11150
rect 1400 11086 1452 11092
rect 1412 10985 1440 11086
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1412 10305 1440 10610
rect 1584 10464 1636 10470
rect 1584 10406 1636 10412
rect 1398 10296 1454 10305
rect 1596 10266 1624 10406
rect 1398 10231 1454 10240
rect 1584 10260 1636 10266
rect 1584 10202 1636 10208
rect 1400 10056 1452 10062
rect 1400 9998 1452 10004
rect 1412 9625 1440 9998
rect 1398 9616 1454 9625
rect 1398 9551 1454 9560
rect 1490 8936 1546 8945
rect 1490 8871 1546 8880
rect 1504 8838 1532 8871
rect 1492 8832 1544 8838
rect 1492 8774 1544 8780
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1412 6934 1440 7346
rect 1400 6928 1452 6934
rect 1398 6896 1400 6905
rect 1452 6896 1454 6905
rect 1398 6831 1454 6840
rect 1780 6322 1808 15098
rect 1872 11762 1900 19910
rect 2240 19854 2268 20198
rect 1952 19848 2004 19854
rect 2228 19848 2280 19854
rect 1952 19790 2004 19796
rect 2226 19816 2228 19825
rect 2280 19816 2282 19825
rect 1964 19174 1992 19790
rect 2226 19751 2282 19760
rect 1952 19168 2004 19174
rect 1952 19110 2004 19116
rect 1952 16992 2004 16998
rect 1952 16934 2004 16940
rect 1860 11756 1912 11762
rect 1860 11698 1912 11704
rect 1768 6316 1820 6322
rect 1768 6258 1820 6264
rect 1490 6216 1546 6225
rect 1490 6151 1492 6160
rect 1544 6151 1546 6160
rect 1492 6122 1544 6128
rect 1492 5568 1544 5574
rect 1490 5536 1492 5545
rect 1544 5536 1546 5545
rect 1490 5471 1546 5480
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1412 4865 1440 5170
rect 1676 5024 1728 5030
rect 1676 4966 1728 4972
rect 1398 4856 1454 4865
rect 1398 4791 1454 4800
rect 1492 4480 1544 4486
rect 1492 4422 1544 4428
rect 1504 4185 1532 4422
rect 1490 4176 1546 4185
rect 664 4140 716 4146
rect 1688 4146 1716 4966
rect 1490 4111 1546 4120
rect 1676 4140 1728 4146
rect 664 4082 716 4088
rect 1676 4082 1728 4088
rect 20 3120 72 3126
rect 20 3062 72 3068
rect 32 800 60 3062
rect 676 800 704 4082
rect 1964 3602 1992 16934
rect 2044 16584 2096 16590
rect 2044 16526 2096 16532
rect 2056 16425 2084 16526
rect 2042 16416 2098 16425
rect 2042 16351 2098 16360
rect 2056 16250 2084 16351
rect 2044 16244 2096 16250
rect 2044 16186 2096 16192
rect 2044 13864 2096 13870
rect 2044 13806 2096 13812
rect 2056 13705 2084 13806
rect 2042 13696 2098 13705
rect 2042 13631 2098 13640
rect 2056 13530 2084 13631
rect 2044 13524 2096 13530
rect 2044 13466 2096 13472
rect 2228 8424 2280 8430
rect 2228 8366 2280 8372
rect 2240 8265 2268 8366
rect 2226 8256 2282 8265
rect 2226 8191 2282 8200
rect 2044 7880 2096 7886
rect 2044 7822 2096 7828
rect 2056 7585 2084 7822
rect 2042 7576 2098 7585
rect 2042 7511 2044 7520
rect 2096 7511 2098 7520
rect 2044 7482 2096 7488
rect 2332 6914 2360 25638
rect 2424 10810 2452 45290
rect 2412 10804 2464 10810
rect 2412 10746 2464 10752
rect 2516 10538 2544 46378
rect 2608 45490 2636 46990
rect 2700 46918 2728 49286
rect 2778 47696 2834 47705
rect 2778 47631 2834 47640
rect 2688 46912 2740 46918
rect 2688 46854 2740 46860
rect 2792 46170 2820 47631
rect 2870 47016 2926 47025
rect 2870 46951 2926 46960
rect 2780 46164 2832 46170
rect 2780 46106 2832 46112
rect 2688 45960 2740 45966
rect 2688 45902 2740 45908
rect 2596 45484 2648 45490
rect 2596 45426 2648 45432
rect 2596 43648 2648 43654
rect 2596 43590 2648 43596
rect 2608 31414 2636 43590
rect 2700 39438 2728 45902
rect 2778 44976 2834 44985
rect 2778 44911 2834 44920
rect 2792 44878 2820 44911
rect 2780 44872 2832 44878
rect 2780 44814 2832 44820
rect 2884 44810 2912 46951
rect 2976 46170 3004 49694
rect 3238 49200 3294 50000
rect 3882 49200 3938 50000
rect 4526 49314 4582 50000
rect 5170 49314 5226 50000
rect 4526 49286 4660 49314
rect 4526 49200 4582 49286
rect 3054 49056 3110 49065
rect 3054 48991 3110 49000
rect 3068 46646 3096 48991
rect 3146 48376 3202 48385
rect 3146 48311 3202 48320
rect 3056 46640 3108 46646
rect 3056 46582 3108 46588
rect 3160 46594 3188 48311
rect 3252 47054 3280 49200
rect 3240 47048 3292 47054
rect 3240 46990 3292 46996
rect 3792 46912 3844 46918
rect 3792 46854 3844 46860
rect 3068 46458 3096 46582
rect 3160 46578 3280 46594
rect 3148 46572 3280 46578
rect 3200 46566 3280 46572
rect 3148 46514 3200 46520
rect 3068 46430 3188 46458
rect 3056 46368 3108 46374
rect 3056 46310 3108 46316
rect 2964 46164 3016 46170
rect 2964 46106 3016 46112
rect 2964 45824 3016 45830
rect 2964 45766 3016 45772
rect 2976 45558 3004 45766
rect 2964 45552 3016 45558
rect 2964 45494 3016 45500
rect 2872 44804 2924 44810
rect 2872 44746 2924 44752
rect 2884 44538 2912 44746
rect 2872 44532 2924 44538
rect 2872 44474 2924 44480
rect 2688 39432 2740 39438
rect 2688 39374 2740 39380
rect 2688 32428 2740 32434
rect 2688 32370 2740 32376
rect 2700 32026 2728 32370
rect 2688 32020 2740 32026
rect 2688 31962 2740 31968
rect 2872 31816 2924 31822
rect 2872 31758 2924 31764
rect 2884 31482 2912 31758
rect 2872 31476 2924 31482
rect 2872 31418 2924 31424
rect 2596 31408 2648 31414
rect 2596 31350 2648 31356
rect 2596 25220 2648 25226
rect 2596 25162 2648 25168
rect 2608 19786 2636 25162
rect 3068 21894 3096 46310
rect 3160 45830 3188 46430
rect 3252 46102 3280 46566
rect 3240 46096 3292 46102
rect 3240 46038 3292 46044
rect 3240 45960 3292 45966
rect 3240 45902 3292 45908
rect 3148 45824 3200 45830
rect 3148 45766 3200 45772
rect 3252 45286 3280 45902
rect 3240 45280 3292 45286
rect 3240 45222 3292 45228
rect 3252 28558 3280 45222
rect 3804 45082 3832 46854
rect 3896 46714 3924 49200
rect 4214 47356 4522 47365
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47291 4522 47300
rect 4632 47258 4660 49286
rect 5170 49286 5396 49314
rect 5170 49200 5226 49286
rect 4620 47252 4672 47258
rect 4620 47194 4672 47200
rect 5368 47054 5396 49286
rect 5814 49200 5870 50000
rect 6458 49314 6514 50000
rect 7102 49314 7158 50000
rect 7746 49314 7802 50000
rect 6458 49286 6592 49314
rect 6458 49200 6514 49286
rect 4804 47048 4856 47054
rect 4804 46990 4856 46996
rect 5356 47048 5408 47054
rect 5356 46990 5408 46996
rect 3976 46980 4028 46986
rect 3976 46922 4028 46928
rect 3884 46708 3936 46714
rect 3884 46650 3936 46656
rect 3896 46170 3924 46650
rect 3884 46164 3936 46170
rect 3884 46106 3936 46112
rect 3792 45076 3844 45082
rect 3792 45018 3844 45024
rect 3700 42628 3752 42634
rect 3700 42570 3752 42576
rect 3712 42022 3740 42570
rect 3700 42016 3752 42022
rect 3700 41958 3752 41964
rect 3240 28552 3292 28558
rect 3240 28494 3292 28500
rect 3240 27328 3292 27334
rect 3240 27270 3292 27276
rect 3056 21888 3108 21894
rect 3056 21830 3108 21836
rect 2872 20256 2924 20262
rect 2872 20198 2924 20204
rect 2884 19854 2912 20198
rect 2872 19848 2924 19854
rect 2872 19790 2924 19796
rect 2596 19780 2648 19786
rect 2596 19722 2648 19728
rect 2504 10532 2556 10538
rect 2504 10474 2556 10480
rect 2148 6886 2360 6914
rect 2148 4826 2176 6886
rect 2320 6384 2372 6390
rect 2320 6326 2372 6332
rect 2136 4820 2188 4826
rect 2136 4762 2188 4768
rect 2148 4622 2176 4762
rect 2136 4616 2188 4622
rect 2136 4558 2188 4564
rect 1952 3596 2004 3602
rect 1952 3538 2004 3544
rect 2228 3596 2280 3602
rect 2228 3538 2280 3544
rect 2240 3505 2268 3538
rect 2226 3496 2282 3505
rect 1952 3460 2004 3466
rect 2226 3431 2282 3440
rect 1952 3402 2004 3408
rect 1308 2848 1360 2854
rect 1308 2790 1360 2796
rect 1320 800 1348 2790
rect 1964 800 1992 3402
rect 2332 3194 2360 6326
rect 2964 5568 3016 5574
rect 2964 5510 3016 5516
rect 2872 5024 2924 5030
rect 2872 4966 2924 4972
rect 2780 4480 2832 4486
rect 2780 4422 2832 4428
rect 2792 4146 2820 4422
rect 2780 4140 2832 4146
rect 2780 4082 2832 4088
rect 2688 3936 2740 3942
rect 2688 3878 2740 3884
rect 2700 3534 2728 3878
rect 2688 3528 2740 3534
rect 2688 3470 2740 3476
rect 2596 3460 2648 3466
rect 2596 3402 2648 3408
rect 2320 3188 2372 3194
rect 2320 3130 2372 3136
rect 2608 800 2636 3402
rect 2792 1465 2820 4082
rect 2884 3058 2912 4966
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2884 2145 2912 2994
rect 2976 2446 3004 5510
rect 3252 3126 3280 27270
rect 3332 26376 3384 26382
rect 3332 26318 3384 26324
rect 3344 19514 3372 26318
rect 3516 20392 3568 20398
rect 3516 20334 3568 20340
rect 3528 20058 3556 20334
rect 3516 20052 3568 20058
rect 3516 19994 3568 20000
rect 3332 19508 3384 19514
rect 3332 19450 3384 19456
rect 3516 19372 3568 19378
rect 3516 19314 3568 19320
rect 3528 17882 3556 19314
rect 3516 17876 3568 17882
rect 3516 17818 3568 17824
rect 3712 8498 3740 41958
rect 3988 31482 4016 46922
rect 4214 46268 4522 46277
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46203 4522 46212
rect 4816 46170 4844 46990
rect 5368 46714 5396 46990
rect 5540 46980 5592 46986
rect 5540 46922 5592 46928
rect 5356 46708 5408 46714
rect 5356 46650 5408 46656
rect 5356 46368 5408 46374
rect 5356 46310 5408 46316
rect 4804 46164 4856 46170
rect 4804 46106 4856 46112
rect 5080 46164 5132 46170
rect 5080 46106 5132 46112
rect 4214 45180 4522 45189
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45115 4522 45124
rect 4620 44736 4672 44742
rect 4620 44678 4672 44684
rect 4214 44092 4522 44101
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44027 4522 44036
rect 4214 43004 4522 43013
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42939 4522 42948
rect 4632 42770 4660 44678
rect 4896 43240 4948 43246
rect 4896 43182 4948 43188
rect 4908 42906 4936 43182
rect 4988 43172 5040 43178
rect 4988 43114 5040 43120
rect 5000 42906 5028 43114
rect 4896 42900 4948 42906
rect 4896 42842 4948 42848
rect 4988 42900 5040 42906
rect 4988 42842 5040 42848
rect 4620 42764 4672 42770
rect 4620 42706 4672 42712
rect 4712 42696 4764 42702
rect 4712 42638 4764 42644
rect 4724 42566 4752 42638
rect 4712 42560 4764 42566
rect 4712 42502 4764 42508
rect 4214 41916 4522 41925
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41851 4522 41860
rect 4068 41540 4120 41546
rect 4068 41482 4120 41488
rect 4080 37942 4108 41482
rect 4214 40828 4522 40837
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40763 4522 40772
rect 4214 39740 4522 39749
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39675 4522 39684
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 4068 37936 4120 37942
rect 4068 37878 4120 37884
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4620 33856 4672 33862
rect 4620 33798 4672 33804
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4068 31884 4120 31890
rect 4068 31826 4120 31832
rect 3976 31476 4028 31482
rect 3976 31418 4028 31424
rect 4080 26926 4108 31826
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4632 29102 4660 33798
rect 4620 29096 4672 29102
rect 4620 29038 4672 29044
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4724 28694 4752 42502
rect 4804 34536 4856 34542
rect 4804 34478 4856 34484
rect 4712 28688 4764 28694
rect 4712 28630 4764 28636
rect 4724 28506 4752 28630
rect 4632 28478 4752 28506
rect 4632 28422 4660 28478
rect 4620 28416 4672 28422
rect 4620 28358 4672 28364
rect 4632 28014 4660 28358
rect 4620 28008 4672 28014
rect 4620 27950 4672 27956
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4068 26920 4120 26926
rect 4068 26862 4120 26868
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4068 21548 4120 21554
rect 4068 21490 4120 21496
rect 4080 16658 4108 21490
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4632 17746 4660 27950
rect 4620 17740 4672 17746
rect 4620 17682 4672 17688
rect 4632 17338 4660 17682
rect 4620 17332 4672 17338
rect 4620 17274 4672 17280
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4068 16652 4120 16658
rect 4068 16594 4120 16600
rect 4632 16574 4660 17274
rect 4632 16546 4752 16574
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4620 13932 4672 13938
rect 4620 13874 4672 13880
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4632 13530 4660 13874
rect 4620 13524 4672 13530
rect 4620 13466 4672 13472
rect 4724 13394 4752 16546
rect 4816 15162 4844 34478
rect 4988 31136 5040 31142
rect 4988 31078 5040 31084
rect 5000 29646 5028 31078
rect 4988 29640 5040 29646
rect 4988 29582 5040 29588
rect 4896 27872 4948 27878
rect 4896 27814 4948 27820
rect 4908 27470 4936 27814
rect 4896 27464 4948 27470
rect 4896 27406 4948 27412
rect 5092 23254 5120 46106
rect 5172 33312 5224 33318
rect 5172 33254 5224 33260
rect 5184 31346 5212 33254
rect 5172 31340 5224 31346
rect 5172 31282 5224 31288
rect 5264 29096 5316 29102
rect 5264 29038 5316 29044
rect 5080 23248 5132 23254
rect 5080 23190 5132 23196
rect 5276 22094 5304 29038
rect 5368 28218 5396 46310
rect 5448 35556 5500 35562
rect 5448 35498 5500 35504
rect 5460 33454 5488 35498
rect 5448 33448 5500 33454
rect 5448 33390 5500 33396
rect 5460 33114 5488 33390
rect 5448 33108 5500 33114
rect 5448 33050 5500 33056
rect 5460 31414 5488 33050
rect 5552 31958 5580 46922
rect 5828 46714 5856 49200
rect 6460 47184 6512 47190
rect 6460 47126 6512 47132
rect 5816 46708 5868 46714
rect 5816 46650 5868 46656
rect 5540 31952 5592 31958
rect 5540 31894 5592 31900
rect 5448 31408 5500 31414
rect 5448 31350 5500 31356
rect 5356 28212 5408 28218
rect 5356 28154 5408 28160
rect 5448 27396 5500 27402
rect 5448 27338 5500 27344
rect 5276 22066 5396 22094
rect 5368 21690 5396 22066
rect 5356 21684 5408 21690
rect 5356 21626 5408 21632
rect 5368 21010 5396 21626
rect 5356 21004 5408 21010
rect 5356 20946 5408 20952
rect 5368 20058 5396 20946
rect 5356 20052 5408 20058
rect 5356 19994 5408 20000
rect 5460 19990 5488 27338
rect 5632 27056 5684 27062
rect 5632 26998 5684 27004
rect 5448 19984 5500 19990
rect 5448 19926 5500 19932
rect 4896 17536 4948 17542
rect 4896 17478 4948 17484
rect 4804 15156 4856 15162
rect 4804 15098 4856 15104
rect 4804 15020 4856 15026
rect 4804 14962 4856 14968
rect 4712 13388 4764 13394
rect 4712 13330 4764 13336
rect 4724 13190 4752 13330
rect 4712 13184 4764 13190
rect 4712 13126 4764 13132
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 3976 11892 4028 11898
rect 3976 11834 4028 11840
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3884 4480 3936 4486
rect 3884 4422 3936 4428
rect 3332 4140 3384 4146
rect 3332 4082 3384 4088
rect 3240 3120 3292 3126
rect 3240 3062 3292 3068
rect 3344 2825 3372 4082
rect 3700 3936 3752 3942
rect 3700 3878 3752 3884
rect 3712 3534 3740 3878
rect 3700 3528 3752 3534
rect 3700 3470 3752 3476
rect 3330 2816 3386 2825
rect 3330 2751 3386 2760
rect 3896 2514 3924 4422
rect 3988 3738 4016 11834
rect 4620 11756 4672 11762
rect 4620 11698 4672 11704
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7274 4660 11698
rect 4724 11558 4752 13126
rect 4816 11898 4844 14962
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 4712 11552 4764 11558
rect 4712 11494 4764 11500
rect 4620 7268 4672 7274
rect 4620 7210 4672 7216
rect 4724 7154 4752 11494
rect 4908 7342 4936 17478
rect 5080 13320 5132 13326
rect 5080 13262 5132 13268
rect 4896 7336 4948 7342
rect 4896 7278 4948 7284
rect 4632 7126 4752 7154
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4632 5846 4660 7126
rect 5092 7018 5120 13262
rect 4724 6990 5120 7018
rect 4620 5840 4672 5846
rect 4620 5782 4672 5788
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4724 4026 4752 6990
rect 4804 5024 4856 5030
rect 4804 4966 4856 4972
rect 4632 3998 4752 4026
rect 4068 3936 4120 3942
rect 4068 3878 4120 3884
rect 3976 3732 4028 3738
rect 3976 3674 4028 3680
rect 4080 3058 4108 3878
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4632 3670 4660 3998
rect 4712 3936 4764 3942
rect 4712 3878 4764 3884
rect 4620 3664 4672 3670
rect 4620 3606 4672 3612
rect 4724 3602 4752 3878
rect 4712 3596 4764 3602
rect 4712 3538 4764 3544
rect 4620 3392 4672 3398
rect 4620 3334 4672 3340
rect 4632 3058 4660 3334
rect 4068 3052 4120 3058
rect 4068 2994 4120 3000
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 3884 2508 3936 2514
rect 3884 2450 3936 2456
rect 2964 2440 3016 2446
rect 2964 2382 3016 2388
rect 2870 2136 2926 2145
rect 2870 2071 2926 2080
rect 2778 1456 2834 1465
rect 2778 1391 2834 1400
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 2976 785 3004 2382
rect 3240 2304 3292 2310
rect 3240 2246 3292 2252
rect 3252 800 3280 2246
rect 3896 800 3924 2450
rect 4632 2122 4660 2994
rect 4816 2446 4844 4966
rect 5644 3738 5672 26998
rect 6368 26920 6420 26926
rect 6368 26862 6420 26868
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 5816 5568 5868 5574
rect 5816 5510 5868 5516
rect 5828 5234 5856 5510
rect 6196 5370 6224 10610
rect 6380 5710 6408 26862
rect 6472 20942 6500 47126
rect 6564 47054 6592 49286
rect 7102 49286 7236 49314
rect 7102 49200 7158 49286
rect 7208 47122 7236 49286
rect 7746 49286 7972 49314
rect 7746 49200 7802 49286
rect 7196 47116 7248 47122
rect 7196 47058 7248 47064
rect 6552 47048 6604 47054
rect 6552 46990 6604 46996
rect 6564 46458 6592 46990
rect 7208 46714 7236 47058
rect 7472 47048 7524 47054
rect 7472 46990 7524 46996
rect 7196 46708 7248 46714
rect 7196 46650 7248 46656
rect 6564 46430 6684 46458
rect 6552 46368 6604 46374
rect 6552 46310 6604 46316
rect 6564 35630 6592 46310
rect 6656 46170 6684 46430
rect 6644 46164 6696 46170
rect 6644 46106 6696 46112
rect 7484 44810 7512 46990
rect 7944 46714 7972 49286
rect 8390 49200 8446 50000
rect 9034 49314 9090 50000
rect 9678 49314 9734 50000
rect 10966 49314 11022 50000
rect 9034 49286 9168 49314
rect 9034 49200 9090 49286
rect 8404 47054 8432 49200
rect 8392 47048 8444 47054
rect 8392 46990 8444 46996
rect 8944 47048 8996 47054
rect 8944 46990 8996 46996
rect 7932 46708 7984 46714
rect 7932 46650 7984 46656
rect 8300 46572 8352 46578
rect 8300 46514 8352 46520
rect 8312 45898 8340 46514
rect 8392 46504 8444 46510
rect 8392 46446 8444 46452
rect 8300 45892 8352 45898
rect 8300 45834 8352 45840
rect 7472 44804 7524 44810
rect 7472 44746 7524 44752
rect 8404 38010 8432 46446
rect 8956 46170 8984 46990
rect 9140 46578 9168 49286
rect 9678 49286 9904 49314
rect 9678 49200 9734 49286
rect 9876 47258 9904 49286
rect 10796 49286 11022 49314
rect 9864 47252 9916 47258
rect 9864 47194 9916 47200
rect 10796 47054 10824 49286
rect 10966 49200 11022 49286
rect 11610 49314 11666 50000
rect 12254 49314 12310 50000
rect 12898 49314 12954 50000
rect 13542 49314 13598 50000
rect 11610 49286 11744 49314
rect 11610 49200 11666 49286
rect 10968 47456 11020 47462
rect 10968 47398 11020 47404
rect 10980 47258 11008 47398
rect 10968 47252 11020 47258
rect 10968 47194 11020 47200
rect 10048 47048 10100 47054
rect 10048 46990 10100 46996
rect 10784 47048 10836 47054
rect 10784 46990 10836 46996
rect 9220 46980 9272 46986
rect 9220 46922 9272 46928
rect 9128 46572 9180 46578
rect 9128 46514 9180 46520
rect 8944 46164 8996 46170
rect 8944 46106 8996 46112
rect 9036 45892 9088 45898
rect 9036 45834 9088 45840
rect 8392 38004 8444 38010
rect 8392 37946 8444 37952
rect 8576 37868 8628 37874
rect 8576 37810 8628 37816
rect 8588 37466 8616 37810
rect 8576 37460 8628 37466
rect 8576 37402 8628 37408
rect 8760 35692 8812 35698
rect 8760 35634 8812 35640
rect 6552 35624 6604 35630
rect 6552 35566 6604 35572
rect 8772 35494 8800 35634
rect 8760 35488 8812 35494
rect 8760 35430 8812 35436
rect 8208 23656 8260 23662
rect 8208 23598 8260 23604
rect 6460 20936 6512 20942
rect 6460 20878 6512 20884
rect 6472 20602 6500 20878
rect 7472 20800 7524 20806
rect 7472 20742 7524 20748
rect 6460 20596 6512 20602
rect 6460 20538 6512 20544
rect 7484 13394 7512 20742
rect 8024 17672 8076 17678
rect 8024 17614 8076 17620
rect 7472 13388 7524 13394
rect 7472 13330 7524 13336
rect 6368 5704 6420 5710
rect 6368 5646 6420 5652
rect 6184 5364 6236 5370
rect 6184 5306 6236 5312
rect 5816 5228 5868 5234
rect 5816 5170 5868 5176
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5644 3058 5672 3674
rect 6184 3392 6236 3398
rect 6184 3334 6236 3340
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 5172 2848 5224 2854
rect 5172 2790 5224 2796
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 4540 2094 4660 2122
rect 4540 800 4568 2094
rect 5184 800 5212 2790
rect 6196 2446 6224 3334
rect 7104 3052 7156 3058
rect 7104 2994 7156 3000
rect 5816 2440 5868 2446
rect 5816 2382 5868 2388
rect 6184 2440 6236 2446
rect 6184 2382 6236 2388
rect 5724 2304 5776 2310
rect 5724 2246 5776 2252
rect 5736 2038 5764 2246
rect 5724 2032 5776 2038
rect 5724 1974 5776 1980
rect 5828 800 5856 2382
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 6472 800 6500 2246
rect 7116 800 7144 2994
rect 8036 2650 8064 17614
rect 8220 16998 8248 23598
rect 8208 16992 8260 16998
rect 8208 16934 8260 16940
rect 8300 11824 8352 11830
rect 8300 11766 8352 11772
rect 8312 10810 8340 11766
rect 8300 10804 8352 10810
rect 8300 10746 8352 10752
rect 8312 10606 8340 10746
rect 8300 10600 8352 10606
rect 8300 10542 8352 10548
rect 8484 5636 8536 5642
rect 8484 5578 8536 5584
rect 8496 3194 8524 5578
rect 8484 3188 8536 3194
rect 8484 3130 8536 3136
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 8404 2854 8432 2994
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 8024 2644 8076 2650
rect 8024 2586 8076 2592
rect 7748 2372 7800 2378
rect 7748 2314 7800 2320
rect 7760 800 7788 2314
rect 8404 800 8432 2790
rect 8772 2310 8800 35430
rect 9048 29578 9076 45834
rect 9036 29572 9088 29578
rect 9036 29514 9088 29520
rect 9128 18624 9180 18630
rect 9128 18566 9180 18572
rect 9036 2848 9088 2854
rect 9036 2790 9088 2796
rect 9048 2378 9076 2790
rect 9140 2650 9168 18566
rect 9232 14006 9260 46922
rect 10060 46374 10088 46990
rect 10796 46714 10824 46990
rect 10784 46708 10836 46714
rect 10784 46650 10836 46656
rect 11716 46578 11744 49286
rect 11992 49286 12310 49314
rect 11992 47054 12020 49286
rect 12254 49200 12310 49286
rect 12636 49286 12954 49314
rect 12636 47054 12664 49286
rect 12898 49200 12954 49286
rect 13280 49286 13598 49314
rect 13280 47054 13308 49286
rect 13542 49200 13598 49286
rect 14186 49314 14242 50000
rect 14830 49314 14886 50000
rect 14186 49286 14320 49314
rect 14186 49200 14242 49286
rect 13820 47524 13872 47530
rect 13820 47466 13872 47472
rect 11980 47048 12032 47054
rect 11980 46990 12032 46996
rect 12440 47048 12492 47054
rect 12440 46990 12492 46996
rect 12624 47048 12676 47054
rect 12624 46990 12676 46996
rect 13268 47048 13320 47054
rect 13268 46990 13320 46996
rect 11704 46572 11756 46578
rect 11704 46514 11756 46520
rect 10048 46368 10100 46374
rect 10048 46310 10100 46316
rect 10692 46368 10744 46374
rect 10692 46310 10744 46316
rect 9496 42628 9548 42634
rect 9496 42570 9548 42576
rect 9508 37262 9536 42570
rect 10324 39432 10376 39438
rect 10324 39374 10376 39380
rect 9956 37324 10008 37330
rect 9956 37266 10008 37272
rect 9496 37256 9548 37262
rect 9496 37198 9548 37204
rect 9968 36582 9996 37266
rect 9956 36576 10008 36582
rect 9956 36518 10008 36524
rect 10336 23186 10364 39374
rect 10324 23180 10376 23186
rect 10324 23122 10376 23128
rect 10232 23112 10284 23118
rect 10232 23054 10284 23060
rect 10244 22778 10272 23054
rect 10232 22772 10284 22778
rect 10232 22714 10284 22720
rect 10508 22636 10560 22642
rect 10508 22578 10560 22584
rect 10416 18828 10468 18834
rect 10416 18770 10468 18776
rect 10324 17536 10376 17542
rect 10324 17478 10376 17484
rect 9220 14000 9272 14006
rect 9220 13942 9272 13948
rect 9772 11620 9824 11626
rect 9772 11562 9824 11568
rect 9588 5568 9640 5574
rect 9588 5510 9640 5516
rect 9496 3528 9548 3534
rect 9496 3470 9548 3476
rect 9508 3126 9536 3470
rect 9496 3120 9548 3126
rect 9496 3062 9548 3068
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 9600 2446 9628 5510
rect 9680 4004 9732 4010
rect 9680 3946 9732 3952
rect 9692 3126 9720 3946
rect 9784 3194 9812 11562
rect 10336 4146 10364 17478
rect 10324 4140 10376 4146
rect 10324 4082 10376 4088
rect 10428 3194 10456 18770
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 9680 3120 9732 3126
rect 9680 3062 9732 3068
rect 9784 2446 9812 3130
rect 10428 2446 10456 3130
rect 10520 2514 10548 22578
rect 10600 12844 10652 12850
rect 10600 12786 10652 12792
rect 10612 12442 10640 12786
rect 10600 12436 10652 12442
rect 10600 12378 10652 12384
rect 10704 6866 10732 46310
rect 11716 46170 11744 46514
rect 11992 46170 12020 46990
rect 11704 46164 11756 46170
rect 11704 46106 11756 46112
rect 11980 46164 12032 46170
rect 11980 46106 12032 46112
rect 12452 42770 12480 46990
rect 12636 45558 12664 46990
rect 12716 46368 12768 46374
rect 12716 46310 12768 46316
rect 12728 46170 12756 46310
rect 12716 46164 12768 46170
rect 12716 46106 12768 46112
rect 13280 45966 13308 46990
rect 13832 46714 13860 47466
rect 14292 47122 14320 49286
rect 14830 49286 15148 49314
rect 14830 49200 14886 49286
rect 14464 47252 14516 47258
rect 14464 47194 14516 47200
rect 13912 47116 13964 47122
rect 13912 47058 13964 47064
rect 14280 47116 14332 47122
rect 14280 47058 14332 47064
rect 13820 46708 13872 46714
rect 13820 46650 13872 46656
rect 13728 46572 13780 46578
rect 13728 46514 13780 46520
rect 13452 46368 13504 46374
rect 13452 46310 13504 46316
rect 13464 45966 13492 46310
rect 13268 45960 13320 45966
rect 13268 45902 13320 45908
rect 13452 45960 13504 45966
rect 13452 45902 13504 45908
rect 12624 45552 12676 45558
rect 12624 45494 12676 45500
rect 13740 45354 13768 46514
rect 13924 45558 13952 47058
rect 14372 46640 14424 46646
rect 14372 46582 14424 46588
rect 14280 46368 14332 46374
rect 14280 46310 14332 46316
rect 14292 45966 14320 46310
rect 14280 45960 14332 45966
rect 14280 45902 14332 45908
rect 13912 45552 13964 45558
rect 13912 45494 13964 45500
rect 13728 45348 13780 45354
rect 13728 45290 13780 45296
rect 14384 45286 14412 46582
rect 14372 45280 14424 45286
rect 14372 45222 14424 45228
rect 12440 42764 12492 42770
rect 12440 42706 12492 42712
rect 12256 39364 12308 39370
rect 12256 39306 12308 39312
rect 11152 22568 11204 22574
rect 11152 22510 11204 22516
rect 11164 22098 11192 22510
rect 11152 22092 11204 22098
rect 11152 22034 11204 22040
rect 12268 20058 12296 39306
rect 14280 31340 14332 31346
rect 14280 31282 14332 31288
rect 14292 30802 14320 31282
rect 14280 30796 14332 30802
rect 14280 30738 14332 30744
rect 13636 24200 13688 24206
rect 13636 24142 13688 24148
rect 13648 23866 13676 24142
rect 13636 23860 13688 23866
rect 13636 23802 13688 23808
rect 12808 20256 12860 20262
rect 12808 20198 12860 20204
rect 12256 20052 12308 20058
rect 12256 19994 12308 20000
rect 12820 19854 12848 20198
rect 13176 20052 13228 20058
rect 13176 19994 13228 20000
rect 12808 19848 12860 19854
rect 12808 19790 12860 19796
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 12728 19378 12756 19654
rect 12716 19372 12768 19378
rect 12716 19314 12768 19320
rect 12532 19168 12584 19174
rect 12532 19110 12584 19116
rect 12544 18766 12572 19110
rect 12532 18760 12584 18766
rect 12532 18702 12584 18708
rect 12820 12434 12848 19790
rect 13188 19718 13216 19994
rect 13176 19712 13228 19718
rect 13176 19654 13228 19660
rect 14292 18426 14320 30738
rect 14280 18420 14332 18426
rect 14280 18362 14332 18368
rect 12992 18284 13044 18290
rect 12992 18226 13044 18232
rect 13004 17814 13032 18226
rect 12992 17808 13044 17814
rect 12992 17750 13044 17756
rect 13004 12918 13032 17750
rect 13820 16244 13872 16250
rect 13820 16186 13872 16192
rect 12992 12912 13044 12918
rect 12992 12854 13044 12860
rect 12728 12406 12848 12434
rect 11796 12300 11848 12306
rect 11796 12242 11848 12248
rect 11612 12096 11664 12102
rect 11612 12038 11664 12044
rect 11624 11694 11652 12038
rect 11808 11830 11836 12242
rect 11796 11824 11848 11830
rect 11796 11766 11848 11772
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 12164 10464 12216 10470
rect 12164 10406 12216 10412
rect 12176 10062 12204 10406
rect 12164 10056 12216 10062
rect 12164 9998 12216 10004
rect 10692 6860 10744 6866
rect 10692 6802 10744 6808
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 11520 6724 11572 6730
rect 11520 6666 11572 6672
rect 11532 6458 11560 6666
rect 11520 6452 11572 6458
rect 11520 6394 11572 6400
rect 12176 6254 12204 6802
rect 11980 6248 12032 6254
rect 11980 6190 12032 6196
rect 12164 6248 12216 6254
rect 12164 6190 12216 6196
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 10968 3052 11020 3058
rect 10968 2994 11020 3000
rect 10980 2854 11008 2994
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 10508 2508 10560 2514
rect 10508 2450 10560 2456
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 9772 2440 9824 2446
rect 9772 2382 9824 2388
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 9036 2372 9088 2378
rect 9036 2314 9088 2320
rect 8760 2304 8812 2310
rect 8760 2246 8812 2252
rect 9048 800 9076 2314
rect 9680 2304 9732 2310
rect 9680 2246 9732 2252
rect 10324 2304 10376 2310
rect 10324 2246 10376 2252
rect 9692 800 9720 2246
rect 10336 800 10364 2246
rect 10980 800 11008 2790
rect 11624 2446 11652 3334
rect 11992 2922 12020 6190
rect 12268 2990 12296 6190
rect 12728 3194 12756 12406
rect 13832 7954 13860 16186
rect 13912 12640 13964 12646
rect 13912 12582 13964 12588
rect 13820 7948 13872 7954
rect 13820 7890 13872 7896
rect 12808 6112 12860 6118
rect 12808 6054 12860 6060
rect 12992 6112 13044 6118
rect 12992 6054 13044 6060
rect 12820 5778 12848 6054
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 13004 5710 13032 6054
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 13452 4140 13504 4146
rect 13452 4082 13504 4088
rect 13464 3738 13492 4082
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 12716 3188 12768 3194
rect 12716 3130 12768 3136
rect 12900 3052 12952 3058
rect 12900 2994 12952 3000
rect 12256 2984 12308 2990
rect 12256 2926 12308 2932
rect 11980 2916 12032 2922
rect 11980 2858 12032 2864
rect 11612 2440 11664 2446
rect 11612 2382 11664 2388
rect 11624 800 11652 2382
rect 12256 2304 12308 2310
rect 12256 2246 12308 2252
rect 12268 800 12296 2246
rect 12912 800 12940 2994
rect 13464 2774 13492 3674
rect 13924 3602 13952 12582
rect 13912 3596 13964 3602
rect 13912 3538 13964 3544
rect 13924 3058 13952 3538
rect 14384 3534 14412 45222
rect 14476 38350 14504 47194
rect 14648 47048 14700 47054
rect 14648 46990 14700 46996
rect 14464 38344 14516 38350
rect 14464 38286 14516 38292
rect 14556 31272 14608 31278
rect 14556 31214 14608 31220
rect 14568 30938 14596 31214
rect 14556 30932 14608 30938
rect 14556 30874 14608 30880
rect 14660 27130 14688 46990
rect 15120 46170 15148 49286
rect 15474 49200 15530 50000
rect 16118 49200 16174 50000
rect 16762 49200 16818 50000
rect 17406 49314 17462 50000
rect 18050 49314 18106 50000
rect 18694 49314 18750 50000
rect 19338 49314 19394 50000
rect 19982 49314 20038 50000
rect 17406 49286 17908 49314
rect 17406 49200 17462 49286
rect 15384 47116 15436 47122
rect 15384 47058 15436 47064
rect 15292 46504 15344 46510
rect 15292 46446 15344 46452
rect 15200 46368 15252 46374
rect 15200 46310 15252 46316
rect 15212 46170 15240 46310
rect 15108 46164 15160 46170
rect 15108 46106 15160 46112
rect 15200 46164 15252 46170
rect 15200 46106 15252 46112
rect 15304 45554 15332 46446
rect 15396 45966 15424 47058
rect 15488 46714 15516 49200
rect 16132 46918 16160 49200
rect 16776 47258 16804 49200
rect 17880 47274 17908 49286
rect 18050 49286 18368 49314
rect 18050 49200 18106 49286
rect 17880 47258 18000 47274
rect 16764 47252 16816 47258
rect 17880 47252 18012 47258
rect 17880 47246 17960 47252
rect 16764 47194 16816 47200
rect 17960 47194 18012 47200
rect 18052 47184 18104 47190
rect 18052 47126 18104 47132
rect 16672 47048 16724 47054
rect 16672 46990 16724 46996
rect 16948 47048 17000 47054
rect 16948 46990 17000 46996
rect 17960 47048 18012 47054
rect 17960 46990 18012 46996
rect 16684 46918 16712 46990
rect 16120 46912 16172 46918
rect 16120 46854 16172 46860
rect 16672 46912 16724 46918
rect 16672 46854 16724 46860
rect 15476 46708 15528 46714
rect 15476 46650 15528 46656
rect 16212 46572 16264 46578
rect 16212 46514 16264 46520
rect 16028 46028 16080 46034
rect 16028 45970 16080 45976
rect 15384 45960 15436 45966
rect 15384 45902 15436 45908
rect 16040 45830 16068 45970
rect 16028 45824 16080 45830
rect 16028 45766 16080 45772
rect 15212 45526 15332 45554
rect 15212 45286 15240 45526
rect 16040 45286 16068 45766
rect 15200 45280 15252 45286
rect 15200 45222 15252 45228
rect 16028 45280 16080 45286
rect 16028 45222 16080 45228
rect 15016 38344 15068 38350
rect 15016 38286 15068 38292
rect 15028 31958 15056 38286
rect 15212 35494 15240 45222
rect 16224 44742 16252 46514
rect 16488 46504 16540 46510
rect 16488 46446 16540 46452
rect 16500 46034 16528 46446
rect 16488 46028 16540 46034
rect 16488 45970 16540 45976
rect 16684 45082 16712 46854
rect 16672 45076 16724 45082
rect 16672 45018 16724 45024
rect 16212 44736 16264 44742
rect 16212 44678 16264 44684
rect 15476 38956 15528 38962
rect 15476 38898 15528 38904
rect 15488 38010 15516 38898
rect 15476 38004 15528 38010
rect 15476 37946 15528 37952
rect 15200 35488 15252 35494
rect 15200 35430 15252 35436
rect 15108 33380 15160 33386
rect 15108 33322 15160 33328
rect 15120 32842 15148 33322
rect 15108 32836 15160 32842
rect 15108 32778 15160 32784
rect 15016 31952 15068 31958
rect 15016 31894 15068 31900
rect 15212 29238 15240 35430
rect 15292 31816 15344 31822
rect 15292 31758 15344 31764
rect 15304 31414 15332 31758
rect 15292 31408 15344 31414
rect 15292 31350 15344 31356
rect 15752 31136 15804 31142
rect 15752 31078 15804 31084
rect 15764 30802 15792 31078
rect 15752 30796 15804 30802
rect 15752 30738 15804 30744
rect 15200 29232 15252 29238
rect 15200 29174 15252 29180
rect 14648 27124 14700 27130
rect 14648 27066 14700 27072
rect 14832 26988 14884 26994
rect 14832 26930 14884 26936
rect 14556 23656 14608 23662
rect 14556 23598 14608 23604
rect 14568 22982 14596 23598
rect 14556 22976 14608 22982
rect 14556 22918 14608 22924
rect 14568 22710 14596 22918
rect 14556 22704 14608 22710
rect 14556 22646 14608 22652
rect 14568 20058 14596 22646
rect 14556 20052 14608 20058
rect 14556 19994 14608 20000
rect 14568 19922 14596 19994
rect 14556 19916 14608 19922
rect 14556 19858 14608 19864
rect 14464 14000 14516 14006
rect 14464 13942 14516 13948
rect 14476 13870 14504 13942
rect 14464 13864 14516 13870
rect 14464 13806 14516 13812
rect 14648 12436 14700 12442
rect 14648 12378 14700 12384
rect 14660 11830 14688 12378
rect 14648 11824 14700 11830
rect 14648 11766 14700 11772
rect 14556 10600 14608 10606
rect 14556 10542 14608 10548
rect 14568 6254 14596 10542
rect 14660 9654 14688 11766
rect 14844 11762 14872 26930
rect 16224 24342 16252 44678
rect 16764 31680 16816 31686
rect 16764 31622 16816 31628
rect 16776 30666 16804 31622
rect 16764 30660 16816 30666
rect 16764 30602 16816 30608
rect 16960 29782 16988 46990
rect 17408 46980 17460 46986
rect 17408 46922 17460 46928
rect 17420 46714 17448 46922
rect 17408 46708 17460 46714
rect 17408 46650 17460 46656
rect 17776 46368 17828 46374
rect 17776 46310 17828 46316
rect 17132 46164 17184 46170
rect 17132 46106 17184 46112
rect 17144 33522 17172 46106
rect 17316 45824 17368 45830
rect 17316 45766 17368 45772
rect 17328 45558 17356 45766
rect 17316 45552 17368 45558
rect 17316 45494 17368 45500
rect 17788 45490 17816 46310
rect 17868 45824 17920 45830
rect 17868 45766 17920 45772
rect 17776 45484 17828 45490
rect 17776 45426 17828 45432
rect 17592 45348 17644 45354
rect 17592 45290 17644 45296
rect 17224 36032 17276 36038
rect 17224 35974 17276 35980
rect 17132 33516 17184 33522
rect 17132 33458 17184 33464
rect 17144 33114 17172 33458
rect 17132 33108 17184 33114
rect 17132 33050 17184 33056
rect 17236 30870 17264 35974
rect 17604 31754 17632 45290
rect 17880 33658 17908 45766
rect 17972 45354 18000 46990
rect 18064 46034 18092 47126
rect 18052 46028 18104 46034
rect 18052 45970 18104 45976
rect 18340 45966 18368 49286
rect 18694 49286 18828 49314
rect 18694 49200 18750 49286
rect 18800 46578 18828 49286
rect 19338 49286 19656 49314
rect 19338 49200 19394 49286
rect 19628 47054 19656 49286
rect 19982 49286 20300 49314
rect 19982 49200 20038 49286
rect 20076 47524 20128 47530
rect 20076 47466 20128 47472
rect 20088 47258 20116 47466
rect 20076 47252 20128 47258
rect 20076 47194 20128 47200
rect 20272 47054 20300 49286
rect 20626 49200 20682 50000
rect 21270 49200 21326 50000
rect 21914 49200 21970 50000
rect 22558 49314 22614 50000
rect 23202 49314 23258 50000
rect 22480 49286 22614 49314
rect 20640 47274 20668 49200
rect 20640 47258 20760 47274
rect 20640 47252 20772 47258
rect 20640 47246 20720 47252
rect 20720 47194 20772 47200
rect 20444 47116 20496 47122
rect 20444 47058 20496 47064
rect 19340 47048 19392 47054
rect 19340 46990 19392 46996
rect 19616 47048 19668 47054
rect 19616 46990 19668 46996
rect 20260 47048 20312 47054
rect 20260 46990 20312 46996
rect 18788 46572 18840 46578
rect 18788 46514 18840 46520
rect 18328 45960 18380 45966
rect 18328 45902 18380 45908
rect 17960 45348 18012 45354
rect 17960 45290 18012 45296
rect 18340 45082 18368 45902
rect 18800 45626 18828 46514
rect 18972 46368 19024 46374
rect 18972 46310 19024 46316
rect 18788 45620 18840 45626
rect 18788 45562 18840 45568
rect 18328 45076 18380 45082
rect 18328 45018 18380 45024
rect 18512 42764 18564 42770
rect 18512 42706 18564 42712
rect 17868 33652 17920 33658
rect 17868 33594 17920 33600
rect 18236 33312 18288 33318
rect 18236 33254 18288 33260
rect 18248 31890 18276 33254
rect 18236 31884 18288 31890
rect 18236 31826 18288 31832
rect 17604 31726 17724 31754
rect 17224 30864 17276 30870
rect 17224 30806 17276 30812
rect 17236 30258 17264 30806
rect 17224 30252 17276 30258
rect 17224 30194 17276 30200
rect 16948 29776 17000 29782
rect 16948 29718 17000 29724
rect 16212 24336 16264 24342
rect 16212 24278 16264 24284
rect 15200 23520 15252 23526
rect 15200 23462 15252 23468
rect 15212 23186 15240 23462
rect 15200 23180 15252 23186
rect 15200 23122 15252 23128
rect 16672 23112 16724 23118
rect 16672 23054 16724 23060
rect 16684 22778 16712 23054
rect 16672 22772 16724 22778
rect 16672 22714 16724 22720
rect 17132 22568 17184 22574
rect 17132 22510 17184 22516
rect 17316 22568 17368 22574
rect 17316 22510 17368 22516
rect 17144 22234 17172 22510
rect 17132 22228 17184 22234
rect 17132 22170 17184 22176
rect 17328 21894 17356 22510
rect 17316 21888 17368 21894
rect 17316 21830 17368 21836
rect 17592 21888 17644 21894
rect 17592 21830 17644 21836
rect 17604 21418 17632 21830
rect 17592 21412 17644 21418
rect 17592 21354 17644 21360
rect 15476 15904 15528 15910
rect 15476 15846 15528 15852
rect 15488 15570 15516 15846
rect 15476 15564 15528 15570
rect 15476 15506 15528 15512
rect 16304 15496 16356 15502
rect 16304 15438 16356 15444
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 15016 11688 15068 11694
rect 15016 11630 15068 11636
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14752 10266 14780 10610
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 14924 9988 14976 9994
rect 14924 9930 14976 9936
rect 14648 9648 14700 9654
rect 14648 9590 14700 9596
rect 14660 9518 14688 9590
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14936 8634 14964 9930
rect 15028 9450 15056 11630
rect 15108 10464 15160 10470
rect 15108 10406 15160 10412
rect 15120 10062 15148 10406
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15476 9580 15528 9586
rect 15476 9522 15528 9528
rect 15016 9444 15068 9450
rect 15016 9386 15068 9392
rect 14924 8628 14976 8634
rect 14924 8570 14976 8576
rect 14556 6248 14608 6254
rect 14556 6190 14608 6196
rect 14568 5914 14596 6190
rect 14556 5908 14608 5914
rect 14556 5850 14608 5856
rect 15292 4072 15344 4078
rect 15292 4014 15344 4020
rect 14464 3732 14516 3738
rect 14464 3674 14516 3680
rect 14372 3528 14424 3534
rect 14372 3470 14424 3476
rect 13912 3052 13964 3058
rect 13912 2994 13964 3000
rect 13280 2746 13492 2774
rect 13280 2446 13308 2746
rect 14476 2446 14504 3674
rect 14924 3392 14976 3398
rect 14924 3334 14976 3340
rect 14936 3058 14964 3334
rect 15304 3194 15332 4014
rect 15292 3188 15344 3194
rect 15292 3130 15344 3136
rect 14924 3052 14976 3058
rect 14924 2994 14976 3000
rect 14936 2774 14964 2994
rect 14844 2746 14964 2774
rect 13268 2440 13320 2446
rect 13268 2382 13320 2388
rect 14464 2440 14516 2446
rect 14464 2382 14516 2388
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 13556 800 13584 2246
rect 14844 800 14872 2746
rect 15488 2650 15516 9522
rect 16316 8498 16344 15438
rect 17224 10192 17276 10198
rect 17224 10134 17276 10140
rect 15936 8492 15988 8498
rect 15936 8434 15988 8440
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 15568 4480 15620 4486
rect 15568 4422 15620 4428
rect 15476 2644 15528 2650
rect 15476 2586 15528 2592
rect 15580 2446 15608 4422
rect 15948 2650 15976 8434
rect 16120 8288 16172 8294
rect 16120 8230 16172 8236
rect 16132 7954 16160 8230
rect 16120 7948 16172 7954
rect 16120 7890 16172 7896
rect 16120 3936 16172 3942
rect 16120 3878 16172 3884
rect 16132 3534 16160 3878
rect 16120 3528 16172 3534
rect 16120 3470 16172 3476
rect 16120 2848 16172 2854
rect 16120 2790 16172 2796
rect 15936 2644 15988 2650
rect 15936 2586 15988 2592
rect 16132 2446 16160 2790
rect 17236 2514 17264 10134
rect 17316 5908 17368 5914
rect 17316 5850 17368 5856
rect 17328 3602 17356 5850
rect 17500 4004 17552 4010
rect 17500 3946 17552 3952
rect 17512 3602 17540 3946
rect 17316 3596 17368 3602
rect 17500 3596 17552 3602
rect 17368 3556 17448 3584
rect 17316 3538 17368 3544
rect 17420 3448 17448 3556
rect 17500 3538 17552 3544
rect 17500 3460 17552 3466
rect 17420 3420 17500 3448
rect 17500 3402 17552 3408
rect 17592 3392 17644 3398
rect 17592 3334 17644 3340
rect 17604 3194 17632 3334
rect 17592 3188 17644 3194
rect 17592 3130 17644 3136
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17224 2508 17276 2514
rect 17224 2450 17276 2456
rect 15568 2440 15620 2446
rect 15568 2382 15620 2388
rect 16120 2440 16172 2446
rect 16120 2382 16172 2388
rect 15580 2292 15608 2382
rect 15488 2264 15608 2292
rect 15488 800 15516 2264
rect 16132 800 16160 2382
rect 16764 2304 16816 2310
rect 16764 2246 16816 2252
rect 16776 800 16804 2246
rect 17420 800 17448 2994
rect 17696 2446 17724 31726
rect 18052 31272 18104 31278
rect 18052 31214 18104 31220
rect 17960 27396 18012 27402
rect 17960 27338 18012 27344
rect 17972 24818 18000 27338
rect 18064 25702 18092 31214
rect 18236 31136 18288 31142
rect 18236 31078 18288 31084
rect 18144 25900 18196 25906
rect 18144 25842 18196 25848
rect 18052 25696 18104 25702
rect 18052 25638 18104 25644
rect 18156 25294 18184 25842
rect 18144 25288 18196 25294
rect 18144 25230 18196 25236
rect 17960 24812 18012 24818
rect 17960 24754 18012 24760
rect 17972 24138 18000 24754
rect 17960 24132 18012 24138
rect 18012 24092 18092 24120
rect 17960 24074 18012 24080
rect 17960 23724 18012 23730
rect 17960 23666 18012 23672
rect 17972 22098 18000 23666
rect 17960 22092 18012 22098
rect 17960 22034 18012 22040
rect 17776 12096 17828 12102
rect 17776 12038 17828 12044
rect 17788 3194 17816 12038
rect 17972 8362 18000 22034
rect 18064 16726 18092 24092
rect 18156 23798 18184 25230
rect 18248 25226 18276 31078
rect 18236 25220 18288 25226
rect 18236 25162 18288 25168
rect 18144 23792 18196 23798
rect 18144 23734 18196 23740
rect 18248 23730 18276 25162
rect 18328 24200 18380 24206
rect 18328 24142 18380 24148
rect 18236 23724 18288 23730
rect 18236 23666 18288 23672
rect 18340 23322 18368 24142
rect 18328 23316 18380 23322
rect 18328 23258 18380 23264
rect 18524 23186 18552 42706
rect 18604 29096 18656 29102
rect 18604 29038 18656 29044
rect 18616 26926 18644 29038
rect 18604 26920 18656 26926
rect 18604 26862 18656 26868
rect 18616 26586 18644 26862
rect 18604 26580 18656 26586
rect 18604 26522 18656 26528
rect 18616 25906 18644 26522
rect 18984 26042 19012 46310
rect 19352 46170 19380 46990
rect 19574 46812 19882 46821
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46747 19882 46756
rect 20272 46714 20300 46990
rect 20260 46708 20312 46714
rect 20260 46650 20312 46656
rect 19340 46164 19392 46170
rect 19340 46106 19392 46112
rect 19574 45724 19882 45733
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45659 19882 45668
rect 19574 44636 19882 44645
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44571 19882 44580
rect 19574 43548 19882 43557
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43483 19882 43492
rect 19574 42460 19882 42469
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42395 19882 42404
rect 19574 41372 19882 41381
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41307 19882 41316
rect 19248 40996 19300 41002
rect 19248 40938 19300 40944
rect 19260 32570 19288 40938
rect 19574 40284 19882 40293
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40219 19882 40228
rect 19432 39432 19484 39438
rect 19432 39374 19484 39380
rect 19444 38962 19472 39374
rect 19574 39196 19882 39205
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39131 19882 39140
rect 19432 38956 19484 38962
rect 19432 38898 19484 38904
rect 19574 38108 19882 38117
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38043 19882 38052
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 20260 33448 20312 33454
rect 20260 33390 20312 33396
rect 20272 33318 20300 33390
rect 20260 33312 20312 33318
rect 20260 33254 20312 33260
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19248 32564 19300 32570
rect 19248 32506 19300 32512
rect 19260 31958 19288 32506
rect 19248 31952 19300 31958
rect 19248 31894 19300 31900
rect 20168 31884 20220 31890
rect 20168 31826 20220 31832
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19340 29300 19392 29306
rect 19340 29242 19392 29248
rect 19352 28218 19380 29242
rect 20180 28626 20208 31826
rect 19432 28620 19484 28626
rect 19432 28562 19484 28568
rect 20168 28620 20220 28626
rect 20168 28562 20220 28568
rect 19444 28422 19472 28562
rect 19432 28416 19484 28422
rect 19432 28358 19484 28364
rect 20168 28416 20220 28422
rect 20272 28404 20300 33254
rect 20456 31754 20484 47058
rect 21088 47048 21140 47054
rect 21088 46990 21140 46996
rect 20812 46096 20864 46102
rect 20812 46038 20864 46044
rect 20628 42900 20680 42906
rect 20628 42842 20680 42848
rect 20640 42362 20668 42842
rect 20628 42356 20680 42362
rect 20628 42298 20680 42304
rect 20640 41614 20668 42298
rect 20628 41608 20680 41614
rect 20628 41550 20680 41556
rect 20824 41414 20852 46038
rect 20824 41386 20944 41414
rect 20916 40934 20944 41386
rect 20904 40928 20956 40934
rect 20904 40870 20956 40876
rect 20812 39500 20864 39506
rect 20812 39442 20864 39448
rect 20628 39432 20680 39438
rect 20628 39374 20680 39380
rect 20640 39098 20668 39374
rect 20628 39092 20680 39098
rect 20628 39034 20680 39040
rect 20824 38894 20852 39442
rect 20812 38888 20864 38894
rect 20812 38830 20864 38836
rect 20916 35086 20944 40870
rect 20996 39364 21048 39370
rect 20996 39306 21048 39312
rect 21008 38554 21036 39306
rect 20996 38548 21048 38554
rect 20996 38490 21048 38496
rect 20996 38276 21048 38282
rect 20996 38218 21048 38224
rect 20812 35080 20864 35086
rect 20812 35022 20864 35028
rect 20904 35080 20956 35086
rect 20904 35022 20956 35028
rect 20720 32768 20772 32774
rect 20720 32710 20772 32716
rect 20732 32502 20760 32710
rect 20720 32496 20772 32502
rect 20720 32438 20772 32444
rect 20364 31726 20484 31754
rect 20364 29306 20392 31726
rect 20444 29640 20496 29646
rect 20444 29582 20496 29588
rect 20352 29300 20404 29306
rect 20352 29242 20404 29248
rect 20364 28490 20392 29242
rect 20352 28484 20404 28490
rect 20352 28426 20404 28432
rect 20220 28376 20300 28404
rect 20168 28358 20220 28364
rect 19340 28212 19392 28218
rect 19340 28154 19392 28160
rect 19444 27538 19472 28358
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 20180 28014 20208 28358
rect 20168 28008 20220 28014
rect 20168 27950 20220 27956
rect 19432 27532 19484 27538
rect 19432 27474 19484 27480
rect 19444 26790 19472 27474
rect 19984 27328 20036 27334
rect 19984 27270 20036 27276
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19996 27130 20024 27270
rect 19984 27124 20036 27130
rect 19984 27066 20036 27072
rect 19432 26784 19484 26790
rect 19432 26726 19484 26732
rect 18972 26036 19024 26042
rect 18972 25978 19024 25984
rect 18604 25900 18656 25906
rect 18604 25842 18656 25848
rect 18984 25362 19012 25978
rect 19444 25838 19472 26726
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19432 25832 19484 25838
rect 19432 25774 19484 25780
rect 18972 25356 19024 25362
rect 18972 25298 19024 25304
rect 19340 25220 19392 25226
rect 19340 25162 19392 25168
rect 19248 25152 19300 25158
rect 19248 25094 19300 25100
rect 19260 24818 19288 25094
rect 19248 24812 19300 24818
rect 19248 24754 19300 24760
rect 18972 24744 19024 24750
rect 18972 24686 19024 24692
rect 18696 24064 18748 24070
rect 18696 24006 18748 24012
rect 18708 23730 18736 24006
rect 18696 23724 18748 23730
rect 18696 23666 18748 23672
rect 18604 23316 18656 23322
rect 18604 23258 18656 23264
rect 18512 23180 18564 23186
rect 18512 23122 18564 23128
rect 18524 22778 18552 23122
rect 18616 22982 18644 23258
rect 18604 22976 18656 22982
rect 18604 22918 18656 22924
rect 18512 22772 18564 22778
rect 18512 22714 18564 22720
rect 18052 16720 18104 16726
rect 18052 16662 18104 16668
rect 18144 9920 18196 9926
rect 18144 9862 18196 9868
rect 17960 8356 18012 8362
rect 17960 8298 18012 8304
rect 17972 6866 18000 8298
rect 17960 6860 18012 6866
rect 17960 6802 18012 6808
rect 17972 6458 18000 6802
rect 17960 6452 18012 6458
rect 17960 6394 18012 6400
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 17972 3738 18000 4558
rect 18052 4140 18104 4146
rect 18052 4082 18104 4088
rect 18064 3738 18092 4082
rect 17960 3732 18012 3738
rect 17960 3674 18012 3680
rect 18052 3732 18104 3738
rect 18052 3674 18104 3680
rect 17776 3188 17828 3194
rect 17776 3130 17828 3136
rect 18156 2446 18184 9862
rect 18420 3664 18472 3670
rect 18420 3606 18472 3612
rect 18432 3466 18460 3606
rect 18420 3460 18472 3466
rect 18420 3402 18472 3408
rect 18616 2582 18644 22918
rect 18984 14414 19012 24686
rect 19352 24410 19380 25162
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19340 24404 19392 24410
rect 19340 24346 19392 24352
rect 19432 24200 19484 24206
rect 19432 24142 19484 24148
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 19444 23746 19472 24142
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19444 23718 19564 23746
rect 19432 23656 19484 23662
rect 19432 23598 19484 23604
rect 19340 23588 19392 23594
rect 19340 23530 19392 23536
rect 18972 14408 19024 14414
rect 18972 14350 19024 14356
rect 19352 8906 19380 23530
rect 19444 23322 19472 23598
rect 19432 23316 19484 23322
rect 19432 23258 19484 23264
rect 19536 23050 19564 23718
rect 20088 23322 20116 24142
rect 20076 23316 20128 23322
rect 20076 23258 20128 23264
rect 19984 23180 20036 23186
rect 19984 23122 20036 23128
rect 19524 23044 19576 23050
rect 19524 22986 19576 22992
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19996 22778 20024 23122
rect 19984 22772 20036 22778
rect 19984 22714 20036 22720
rect 20076 22772 20128 22778
rect 20076 22714 20128 22720
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19340 8900 19392 8906
rect 19340 8842 19392 8848
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 18696 3052 18748 3058
rect 18696 2994 18748 3000
rect 18604 2576 18656 2582
rect 18604 2518 18656 2524
rect 17684 2440 17736 2446
rect 17684 2382 17736 2388
rect 18144 2440 18196 2446
rect 18144 2382 18196 2388
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 18064 800 18092 2246
rect 18708 800 18736 2994
rect 19340 2304 19392 2310
rect 19340 2246 19392 2252
rect 19984 2304 20036 2310
rect 19984 2246 20036 2252
rect 19352 800 19380 2246
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 800 20024 2246
rect 20088 2106 20116 22714
rect 20180 12442 20208 27950
rect 20364 27674 20392 28426
rect 20456 28218 20484 29582
rect 20536 29572 20588 29578
rect 20536 29514 20588 29520
rect 20548 29102 20576 29514
rect 20536 29096 20588 29102
rect 20536 29038 20588 29044
rect 20444 28212 20496 28218
rect 20444 28154 20496 28160
rect 20352 27668 20404 27674
rect 20352 27610 20404 27616
rect 20444 27328 20496 27334
rect 20444 27270 20496 27276
rect 20456 26994 20484 27270
rect 20444 26988 20496 26994
rect 20444 26930 20496 26936
rect 20628 25832 20680 25838
rect 20628 25774 20680 25780
rect 20352 25696 20404 25702
rect 20352 25638 20404 25644
rect 20364 25294 20392 25638
rect 20640 25430 20668 25774
rect 20628 25424 20680 25430
rect 20628 25366 20680 25372
rect 20352 25288 20404 25294
rect 20352 25230 20404 25236
rect 20640 25158 20668 25366
rect 20628 25152 20680 25158
rect 20628 25094 20680 25100
rect 20640 23254 20668 25094
rect 20628 23248 20680 23254
rect 20628 23190 20680 23196
rect 20260 23044 20312 23050
rect 20260 22986 20312 22992
rect 20272 22778 20300 22986
rect 20260 22772 20312 22778
rect 20260 22714 20312 22720
rect 20640 22710 20668 23190
rect 20628 22704 20680 22710
rect 20628 22646 20680 22652
rect 20352 21888 20404 21894
rect 20352 21830 20404 21836
rect 20364 21554 20392 21830
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 20536 21344 20588 21350
rect 20536 21286 20588 21292
rect 20168 12436 20220 12442
rect 20168 12378 20220 12384
rect 20548 3194 20576 21286
rect 20732 6390 20760 32438
rect 20824 31346 20852 35022
rect 21008 32570 21036 38218
rect 20996 32564 21048 32570
rect 20996 32506 21048 32512
rect 20996 31816 21048 31822
rect 20916 31764 20996 31770
rect 20916 31758 21048 31764
rect 20916 31742 21036 31758
rect 20812 31340 20864 31346
rect 20812 31282 20864 31288
rect 20916 31210 20944 31742
rect 20996 31680 21048 31686
rect 20996 31622 21048 31628
rect 21008 31482 21036 31622
rect 20996 31476 21048 31482
rect 20996 31418 21048 31424
rect 20904 31204 20956 31210
rect 20904 31146 20956 31152
rect 20812 29164 20864 29170
rect 20812 29106 20864 29112
rect 20824 28762 20852 29106
rect 20812 28756 20864 28762
rect 20812 28698 20864 28704
rect 21008 27606 21036 31418
rect 21100 29850 21128 46990
rect 21284 46714 21312 49200
rect 21272 46708 21324 46714
rect 21272 46650 21324 46656
rect 21928 46578 21956 49200
rect 22480 47258 22508 49286
rect 22558 49200 22614 49286
rect 23032 49286 23258 49314
rect 22468 47252 22520 47258
rect 22468 47194 22520 47200
rect 23032 47122 23060 49286
rect 23202 49200 23258 49286
rect 23846 49200 23902 50000
rect 24490 49314 24546 50000
rect 25778 49314 25834 50000
rect 24490 49286 24808 49314
rect 24490 49200 24546 49286
rect 23860 47122 23888 49200
rect 24308 47456 24360 47462
rect 24308 47398 24360 47404
rect 23020 47116 23072 47122
rect 23020 47058 23072 47064
rect 23848 47116 23900 47122
rect 23848 47058 23900 47064
rect 22836 47048 22888 47054
rect 22836 46990 22888 46996
rect 21916 46572 21968 46578
rect 21916 46514 21968 46520
rect 22100 46368 22152 46374
rect 22100 46310 22152 46316
rect 22192 46368 22244 46374
rect 22192 46310 22244 46316
rect 22008 45348 22060 45354
rect 22008 45290 22060 45296
rect 21640 41676 21692 41682
rect 21640 41618 21692 41624
rect 21652 41070 21680 41618
rect 21732 41472 21784 41478
rect 21732 41414 21784 41420
rect 21640 41064 21692 41070
rect 21640 41006 21692 41012
rect 21272 38956 21324 38962
rect 21272 38898 21324 38904
rect 21284 38350 21312 38898
rect 21272 38344 21324 38350
rect 21272 38286 21324 38292
rect 21652 35630 21680 41006
rect 21744 40934 21772 41414
rect 21732 40928 21784 40934
rect 21732 40870 21784 40876
rect 21916 39636 21968 39642
rect 21916 39578 21968 39584
rect 21928 39506 21956 39578
rect 21916 39500 21968 39506
rect 21916 39442 21968 39448
rect 21928 38554 21956 39442
rect 22020 39438 22048 45290
rect 22112 44266 22140 46310
rect 22100 44260 22152 44266
rect 22100 44202 22152 44208
rect 22008 39432 22060 39438
rect 22008 39374 22060 39380
rect 21916 38548 21968 38554
rect 21916 38490 21968 38496
rect 21732 36712 21784 36718
rect 21732 36654 21784 36660
rect 21640 35624 21692 35630
rect 21640 35566 21692 35572
rect 21548 33992 21600 33998
rect 21548 33934 21600 33940
rect 21364 32428 21416 32434
rect 21364 32370 21416 32376
rect 21376 32026 21404 32370
rect 21364 32020 21416 32026
rect 21364 31962 21416 31968
rect 21180 30116 21232 30122
rect 21180 30058 21232 30064
rect 21088 29844 21140 29850
rect 21088 29786 21140 29792
rect 20996 27600 21048 27606
rect 20996 27542 21048 27548
rect 20904 27464 20956 27470
rect 20904 27406 20956 27412
rect 20916 26586 20944 27406
rect 21192 27062 21220 30058
rect 21272 28076 21324 28082
rect 21272 28018 21324 28024
rect 21180 27056 21232 27062
rect 21180 26998 21232 27004
rect 20996 26920 21048 26926
rect 20996 26862 21048 26868
rect 20904 26580 20956 26586
rect 20904 26522 20956 26528
rect 21008 26042 21036 26862
rect 20996 26036 21048 26042
rect 20996 25978 21048 25984
rect 21008 25362 21036 25978
rect 20996 25356 21048 25362
rect 20996 25298 21048 25304
rect 21008 24834 21036 25298
rect 21180 25152 21232 25158
rect 21180 25094 21232 25100
rect 20916 24806 21036 24834
rect 21192 24818 21220 25094
rect 21180 24812 21232 24818
rect 20916 24138 20944 24806
rect 21180 24754 21232 24760
rect 20996 24744 21048 24750
rect 20996 24686 21048 24692
rect 21088 24744 21140 24750
rect 21284 24698 21312 28018
rect 21456 26512 21508 26518
rect 21456 26454 21508 26460
rect 21088 24686 21140 24692
rect 20904 24132 20956 24138
rect 20904 24074 20956 24080
rect 20916 23186 20944 24074
rect 20904 23180 20956 23186
rect 20904 23122 20956 23128
rect 20904 22976 20956 22982
rect 20904 22918 20956 22924
rect 20916 22778 20944 22918
rect 20904 22772 20956 22778
rect 20904 22714 20956 22720
rect 21008 11626 21036 24686
rect 21100 22098 21128 24686
rect 21192 24670 21312 24698
rect 21088 22092 21140 22098
rect 21088 22034 21140 22040
rect 21100 21418 21128 22034
rect 21088 21412 21140 21418
rect 21088 21354 21140 21360
rect 21192 17338 21220 24670
rect 21468 24274 21496 26454
rect 21456 24268 21508 24274
rect 21456 24210 21508 24216
rect 21560 23866 21588 33934
rect 21744 32842 21772 36654
rect 21824 36576 21876 36582
rect 21824 36518 21876 36524
rect 21836 34066 21864 36518
rect 22020 36310 22048 39374
rect 22100 37256 22152 37262
rect 22100 37198 22152 37204
rect 22112 36378 22140 37198
rect 22204 36922 22232 46310
rect 22468 44192 22520 44198
rect 22468 44134 22520 44140
rect 22480 43994 22508 44134
rect 22468 43988 22520 43994
rect 22468 43930 22520 43936
rect 22848 41414 22876 46990
rect 23032 46714 23060 47058
rect 23296 47048 23348 47054
rect 23296 46990 23348 46996
rect 23020 46708 23072 46714
rect 23020 46650 23072 46656
rect 22664 41386 22876 41414
rect 22284 38004 22336 38010
rect 22284 37946 22336 37952
rect 22192 36916 22244 36922
rect 22192 36858 22244 36864
rect 22296 36802 22324 37946
rect 22560 37732 22612 37738
rect 22560 37674 22612 37680
rect 22204 36774 22324 36802
rect 22100 36372 22152 36378
rect 22100 36314 22152 36320
rect 22008 36304 22060 36310
rect 22008 36246 22060 36252
rect 22020 36174 22048 36246
rect 22008 36168 22060 36174
rect 22008 36110 22060 36116
rect 22008 35624 22060 35630
rect 22008 35566 22060 35572
rect 21824 34060 21876 34066
rect 21824 34002 21876 34008
rect 21732 32836 21784 32842
rect 21732 32778 21784 32784
rect 21744 32366 21772 32778
rect 21916 32564 21968 32570
rect 21916 32506 21968 32512
rect 21732 32360 21784 32366
rect 21732 32302 21784 32308
rect 21640 31884 21692 31890
rect 21640 31826 21692 31832
rect 21652 26926 21680 31826
rect 21744 31482 21772 32302
rect 21928 32026 21956 32506
rect 21916 32020 21968 32026
rect 21916 31962 21968 31968
rect 22020 31822 22048 35566
rect 22100 35012 22152 35018
rect 22100 34954 22152 34960
rect 22008 31816 22060 31822
rect 22008 31758 22060 31764
rect 21732 31476 21784 31482
rect 21732 31418 21784 31424
rect 21744 31142 21772 31418
rect 21732 31136 21784 31142
rect 21732 31078 21784 31084
rect 22112 29186 22140 34954
rect 22204 29782 22232 36774
rect 22376 35488 22428 35494
rect 22376 35430 22428 35436
rect 22388 34678 22416 35430
rect 22376 34672 22428 34678
rect 22376 34614 22428 34620
rect 22284 33992 22336 33998
rect 22284 33934 22336 33940
rect 22296 33658 22324 33934
rect 22284 33652 22336 33658
rect 22284 33594 22336 33600
rect 22572 33538 22600 37674
rect 22664 34202 22692 41386
rect 22744 40452 22796 40458
rect 22744 40394 22796 40400
rect 22756 37466 22784 40394
rect 22744 37460 22796 37466
rect 22744 37402 22796 37408
rect 22756 36922 22784 37402
rect 22744 36916 22796 36922
rect 22744 36858 22796 36864
rect 23020 36032 23072 36038
rect 23020 35974 23072 35980
rect 23032 35612 23060 35974
rect 23112 35624 23164 35630
rect 23032 35584 23112 35612
rect 22836 34944 22888 34950
rect 22836 34886 22888 34892
rect 22652 34196 22704 34202
rect 22652 34138 22704 34144
rect 22744 34128 22796 34134
rect 22744 34070 22796 34076
rect 22756 33658 22784 34070
rect 22744 33652 22796 33658
rect 22744 33594 22796 33600
rect 22572 33510 22784 33538
rect 22560 32904 22612 32910
rect 22560 32846 22612 32852
rect 22572 32570 22600 32846
rect 22652 32768 22704 32774
rect 22652 32710 22704 32716
rect 22560 32564 22612 32570
rect 22560 32506 22612 32512
rect 22468 30592 22520 30598
rect 22468 30534 22520 30540
rect 22192 29776 22244 29782
rect 22192 29718 22244 29724
rect 22284 29776 22336 29782
rect 22284 29718 22336 29724
rect 22192 29640 22244 29646
rect 22192 29582 22244 29588
rect 22204 29306 22232 29582
rect 22192 29300 22244 29306
rect 22192 29242 22244 29248
rect 22112 29158 22232 29186
rect 21916 28484 21968 28490
rect 21916 28426 21968 28432
rect 21928 28218 21956 28426
rect 22100 28416 22152 28422
rect 22100 28358 22152 28364
rect 21916 28212 21968 28218
rect 21916 28154 21968 28160
rect 22008 28144 22060 28150
rect 22008 28086 22060 28092
rect 21916 27328 21968 27334
rect 21916 27270 21968 27276
rect 21640 26920 21692 26926
rect 21640 26862 21692 26868
rect 21732 26376 21784 26382
rect 21732 26318 21784 26324
rect 21640 25764 21692 25770
rect 21640 25706 21692 25712
rect 21652 25362 21680 25706
rect 21640 25356 21692 25362
rect 21640 25298 21692 25304
rect 21548 23860 21600 23866
rect 21548 23802 21600 23808
rect 21744 23730 21772 26318
rect 21824 24812 21876 24818
rect 21824 24754 21876 24760
rect 21836 23866 21864 24754
rect 21928 24342 21956 27270
rect 22020 24954 22048 28086
rect 22008 24948 22060 24954
rect 22008 24890 22060 24896
rect 21916 24336 21968 24342
rect 21916 24278 21968 24284
rect 21916 24132 21968 24138
rect 21916 24074 21968 24080
rect 21928 23866 21956 24074
rect 21824 23860 21876 23866
rect 21824 23802 21876 23808
rect 21916 23860 21968 23866
rect 21916 23802 21968 23808
rect 21732 23724 21784 23730
rect 21732 23666 21784 23672
rect 21640 22976 21692 22982
rect 21640 22918 21692 22924
rect 21272 22772 21324 22778
rect 21272 22714 21324 22720
rect 21180 17332 21232 17338
rect 21180 17274 21232 17280
rect 21284 17270 21312 22714
rect 21456 22568 21508 22574
rect 21456 22510 21508 22516
rect 21272 17264 21324 17270
rect 21272 17206 21324 17212
rect 20996 11620 21048 11626
rect 20996 11562 21048 11568
rect 20720 6384 20772 6390
rect 20720 6326 20772 6332
rect 21088 3392 21140 3398
rect 21088 3334 21140 3340
rect 20536 3188 20588 3194
rect 20536 3130 20588 3136
rect 20548 2446 20576 3130
rect 21100 3058 21128 3334
rect 21088 3052 21140 3058
rect 21088 2994 21140 3000
rect 21100 2774 21128 2994
rect 21468 2990 21496 22510
rect 21652 16250 21680 22918
rect 21744 22778 21772 23666
rect 21732 22772 21784 22778
rect 21732 22714 21784 22720
rect 21744 22094 21772 22714
rect 21744 22066 21864 22094
rect 21732 21344 21784 21350
rect 21732 21286 21784 21292
rect 21640 16244 21692 16250
rect 21640 16186 21692 16192
rect 21744 15910 21772 21286
rect 21836 17678 21864 22066
rect 21928 20058 21956 23802
rect 21916 20052 21968 20058
rect 21916 19994 21968 20000
rect 21928 19310 21956 19994
rect 21916 19304 21968 19310
rect 21916 19246 21968 19252
rect 21916 19168 21968 19174
rect 21916 19110 21968 19116
rect 21928 18834 21956 19110
rect 21916 18828 21968 18834
rect 21916 18770 21968 18776
rect 21824 17672 21876 17678
rect 21824 17614 21876 17620
rect 21732 15904 21784 15910
rect 21732 15846 21784 15852
rect 21744 6798 21772 15846
rect 22112 11898 22140 28358
rect 22204 22094 22232 29158
rect 22296 27130 22324 29718
rect 22480 29238 22508 30534
rect 22560 29504 22612 29510
rect 22560 29446 22612 29452
rect 22468 29232 22520 29238
rect 22468 29174 22520 29180
rect 22572 29034 22600 29446
rect 22560 29028 22612 29034
rect 22560 28970 22612 28976
rect 22468 28620 22520 28626
rect 22468 28562 22520 28568
rect 22480 28014 22508 28562
rect 22468 28008 22520 28014
rect 22468 27950 22520 27956
rect 22284 27124 22336 27130
rect 22284 27066 22336 27072
rect 22572 26024 22600 28970
rect 22296 25996 22600 26024
rect 22296 25430 22324 25996
rect 22664 25922 22692 32710
rect 22756 30190 22784 33510
rect 22848 32978 22876 34886
rect 22836 32972 22888 32978
rect 22836 32914 22888 32920
rect 22928 31340 22980 31346
rect 22928 31282 22980 31288
rect 22744 30184 22796 30190
rect 22744 30126 22796 30132
rect 22376 25900 22428 25906
rect 22376 25842 22428 25848
rect 22572 25894 22692 25922
rect 22284 25424 22336 25430
rect 22284 25366 22336 25372
rect 22296 24750 22324 25366
rect 22284 24744 22336 24750
rect 22284 24686 22336 24692
rect 22296 24018 22324 24686
rect 22388 24138 22416 25842
rect 22572 25838 22600 25894
rect 22468 25832 22520 25838
rect 22468 25774 22520 25780
rect 22560 25832 22612 25838
rect 22560 25774 22612 25780
rect 22480 24290 22508 25774
rect 22572 24410 22600 25774
rect 22652 25696 22704 25702
rect 22652 25638 22704 25644
rect 22560 24404 22612 24410
rect 22560 24346 22612 24352
rect 22480 24262 22600 24290
rect 22468 24200 22520 24206
rect 22468 24142 22520 24148
rect 22376 24132 22428 24138
rect 22376 24074 22428 24080
rect 22296 23990 22416 24018
rect 22388 23662 22416 23990
rect 22284 23656 22336 23662
rect 22284 23598 22336 23604
rect 22376 23656 22428 23662
rect 22376 23598 22428 23604
rect 22296 22982 22324 23598
rect 22388 23526 22416 23598
rect 22376 23520 22428 23526
rect 22376 23462 22428 23468
rect 22376 23180 22428 23186
rect 22376 23122 22428 23128
rect 22284 22976 22336 22982
rect 22284 22918 22336 22924
rect 22388 22098 22416 23122
rect 22480 22778 22508 24142
rect 22572 23594 22600 24262
rect 22560 23588 22612 23594
rect 22560 23530 22612 23536
rect 22560 23248 22612 23254
rect 22560 23190 22612 23196
rect 22468 22772 22520 22778
rect 22468 22714 22520 22720
rect 22572 22658 22600 23190
rect 22480 22630 22600 22658
rect 22480 22098 22508 22630
rect 22204 22066 22324 22094
rect 22296 19378 22324 22066
rect 22376 22092 22428 22098
rect 22376 22034 22428 22040
rect 22468 22092 22520 22098
rect 22468 22034 22520 22040
rect 22284 19372 22336 19378
rect 22284 19314 22336 19320
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 21732 6792 21784 6798
rect 21732 6734 21784 6740
rect 21548 6724 21600 6730
rect 21548 6666 21600 6672
rect 21456 2984 21508 2990
rect 21456 2926 21508 2932
rect 21560 2922 21588 6666
rect 21548 2916 21600 2922
rect 21548 2858 21600 2864
rect 21916 2848 21968 2854
rect 21916 2790 21968 2796
rect 22008 2848 22060 2854
rect 22008 2790 22060 2796
rect 21100 2746 21312 2774
rect 20536 2440 20588 2446
rect 20536 2382 20588 2388
rect 20628 2304 20680 2310
rect 20628 2246 20680 2252
rect 20076 2100 20128 2106
rect 20076 2042 20128 2048
rect 20640 800 20668 2246
rect 21284 800 21312 2746
rect 21928 2514 21956 2790
rect 21916 2508 21968 2514
rect 21916 2450 21968 2456
rect 22020 2394 22048 2790
rect 22296 2514 22324 19314
rect 22480 18426 22508 22034
rect 22468 18420 22520 18426
rect 22468 18362 22520 18368
rect 22664 18358 22692 25638
rect 22940 25362 22968 31282
rect 23032 30682 23060 35584
rect 23112 35566 23164 35572
rect 23308 33590 23336 46990
rect 23480 46096 23532 46102
rect 23480 46038 23532 46044
rect 23492 36922 23520 46038
rect 23756 43716 23808 43722
rect 23756 43658 23808 43664
rect 23480 36916 23532 36922
rect 23480 36858 23532 36864
rect 23492 35834 23520 36858
rect 23768 36378 23796 43658
rect 24320 36378 24348 47398
rect 24400 47116 24452 47122
rect 24400 47058 24452 47064
rect 24412 46170 24440 47058
rect 24676 47048 24728 47054
rect 24676 46990 24728 46996
rect 24400 46164 24452 46170
rect 24400 46106 24452 46112
rect 23756 36372 23808 36378
rect 23756 36314 23808 36320
rect 24308 36372 24360 36378
rect 24308 36314 24360 36320
rect 23480 35828 23532 35834
rect 23480 35770 23532 35776
rect 23768 35766 23796 36314
rect 24320 35834 24348 36314
rect 24308 35828 24360 35834
rect 24308 35770 24360 35776
rect 23756 35760 23808 35766
rect 23756 35702 23808 35708
rect 23768 35154 23796 35702
rect 23756 35148 23808 35154
rect 23756 35090 23808 35096
rect 23768 34746 23796 35090
rect 23756 34740 23808 34746
rect 23756 34682 23808 34688
rect 23664 34672 23716 34678
rect 23664 34614 23716 34620
rect 23296 33584 23348 33590
rect 23296 33526 23348 33532
rect 23296 33380 23348 33386
rect 23296 33322 23348 33328
rect 23204 32224 23256 32230
rect 23204 32166 23256 32172
rect 23112 32020 23164 32026
rect 23112 31962 23164 31968
rect 23124 31890 23152 31962
rect 23112 31884 23164 31890
rect 23112 31826 23164 31832
rect 23124 31482 23152 31826
rect 23112 31476 23164 31482
rect 23112 31418 23164 31424
rect 23216 31414 23244 32166
rect 23204 31408 23256 31414
rect 23204 31350 23256 31356
rect 23032 30654 23152 30682
rect 23020 30592 23072 30598
rect 23020 30534 23072 30540
rect 23032 30326 23060 30534
rect 23020 30320 23072 30326
rect 23020 30262 23072 30268
rect 23020 30184 23072 30190
rect 23020 30126 23072 30132
rect 22928 25356 22980 25362
rect 22928 25298 22980 25304
rect 22744 24200 22796 24206
rect 22744 24142 22796 24148
rect 22652 18352 22704 18358
rect 22652 18294 22704 18300
rect 22560 7404 22612 7410
rect 22560 7346 22612 7352
rect 22572 6866 22600 7346
rect 22560 6860 22612 6866
rect 22560 6802 22612 6808
rect 22756 3602 22784 24142
rect 23032 23186 23060 30126
rect 23124 29782 23152 30654
rect 23112 29776 23164 29782
rect 23112 29718 23164 29724
rect 23124 29578 23152 29718
rect 23112 29572 23164 29578
rect 23112 29514 23164 29520
rect 23308 29458 23336 33322
rect 23388 33040 23440 33046
rect 23388 32982 23440 32988
rect 23400 32026 23428 32982
rect 23572 32496 23624 32502
rect 23572 32438 23624 32444
rect 23388 32020 23440 32026
rect 23388 31962 23440 31968
rect 23584 31890 23612 32438
rect 23572 31884 23624 31890
rect 23572 31826 23624 31832
rect 23676 30326 23704 34614
rect 23756 33856 23808 33862
rect 23756 33798 23808 33804
rect 23768 32842 23796 33798
rect 23756 32836 23808 32842
rect 23756 32778 23808 32784
rect 23768 32366 23796 32778
rect 23756 32360 23808 32366
rect 23756 32302 23808 32308
rect 23848 32292 23900 32298
rect 23848 32234 23900 32240
rect 23860 31686 23888 32234
rect 23848 31680 23900 31686
rect 23848 31622 23900 31628
rect 24308 31680 24360 31686
rect 24308 31622 24360 31628
rect 23860 31482 23888 31622
rect 23848 31476 23900 31482
rect 23848 31418 23900 31424
rect 24320 30598 24348 31622
rect 24492 31136 24544 31142
rect 24492 31078 24544 31084
rect 24504 30870 24532 31078
rect 24492 30864 24544 30870
rect 24492 30806 24544 30812
rect 24308 30592 24360 30598
rect 24308 30534 24360 30540
rect 23664 30320 23716 30326
rect 23664 30262 23716 30268
rect 23676 29850 23704 30262
rect 23848 30048 23900 30054
rect 23848 29990 23900 29996
rect 23388 29844 23440 29850
rect 23388 29786 23440 29792
rect 23664 29844 23716 29850
rect 23664 29786 23716 29792
rect 23124 29430 23336 29458
rect 23124 28218 23152 29430
rect 23400 29306 23428 29786
rect 23860 29646 23888 29990
rect 23848 29640 23900 29646
rect 23848 29582 23900 29588
rect 23296 29300 23348 29306
rect 23296 29242 23348 29248
rect 23388 29300 23440 29306
rect 23388 29242 23440 29248
rect 23308 29102 23336 29242
rect 23296 29096 23348 29102
rect 23296 29038 23348 29044
rect 23204 29028 23256 29034
rect 23204 28970 23256 28976
rect 23112 28212 23164 28218
rect 23112 28154 23164 28160
rect 23124 27674 23152 28154
rect 23112 27668 23164 27674
rect 23112 27610 23164 27616
rect 23124 27470 23152 27610
rect 23112 27464 23164 27470
rect 23112 27406 23164 27412
rect 23124 27130 23152 27406
rect 23112 27124 23164 27130
rect 23112 27066 23164 27072
rect 23216 26790 23244 28970
rect 23480 27872 23532 27878
rect 23480 27814 23532 27820
rect 23204 26784 23256 26790
rect 23204 26726 23256 26732
rect 23216 26450 23244 26726
rect 23388 26580 23440 26586
rect 23388 26522 23440 26528
rect 23204 26444 23256 26450
rect 23204 26386 23256 26392
rect 23400 26246 23428 26522
rect 23388 26240 23440 26246
rect 23388 26182 23440 26188
rect 23112 25288 23164 25294
rect 23112 25230 23164 25236
rect 23124 24698 23152 25230
rect 23400 24886 23428 26182
rect 23388 24880 23440 24886
rect 23388 24822 23440 24828
rect 23124 24670 23244 24698
rect 23112 24608 23164 24614
rect 23112 24550 23164 24556
rect 23124 23730 23152 24550
rect 23216 24274 23244 24670
rect 23204 24268 23256 24274
rect 23204 24210 23256 24216
rect 23296 24064 23348 24070
rect 23296 24006 23348 24012
rect 23112 23724 23164 23730
rect 23112 23666 23164 23672
rect 23308 23594 23336 24006
rect 23388 23656 23440 23662
rect 23388 23598 23440 23604
rect 23296 23588 23348 23594
rect 23296 23530 23348 23536
rect 23020 23180 23072 23186
rect 23020 23122 23072 23128
rect 22928 23112 22980 23118
rect 22928 23054 22980 23060
rect 22940 22642 22968 23054
rect 23296 22976 23348 22982
rect 23296 22918 23348 22924
rect 23308 22642 23336 22918
rect 22928 22636 22980 22642
rect 22928 22578 22980 22584
rect 23296 22636 23348 22642
rect 23296 22578 23348 22584
rect 22836 22568 22888 22574
rect 22888 22516 22968 22522
rect 22836 22510 22968 22516
rect 22848 22494 22968 22510
rect 22940 21894 22968 22494
rect 22928 21888 22980 21894
rect 22928 21830 22980 21836
rect 22940 19854 22968 21830
rect 22928 19848 22980 19854
rect 22928 19790 22980 19796
rect 23400 10538 23428 23598
rect 23492 11762 23520 27814
rect 23860 26042 23888 29582
rect 23848 26036 23900 26042
rect 23848 25978 23900 25984
rect 23664 25288 23716 25294
rect 23664 25230 23716 25236
rect 23676 24954 23704 25230
rect 23664 24948 23716 24954
rect 23664 24890 23716 24896
rect 24216 24744 24268 24750
rect 24216 24686 24268 24692
rect 24228 23866 24256 24686
rect 24216 23860 24268 23866
rect 24216 23802 24268 23808
rect 23664 23044 23716 23050
rect 23664 22986 23716 22992
rect 23572 22772 23624 22778
rect 23572 22714 23624 22720
rect 23584 22234 23612 22714
rect 23676 22438 23704 22986
rect 23664 22432 23716 22438
rect 23664 22374 23716 22380
rect 23572 22228 23624 22234
rect 23572 22170 23624 22176
rect 24320 21418 24348 30534
rect 24400 25424 24452 25430
rect 24400 25366 24452 25372
rect 24412 25158 24440 25366
rect 24400 25152 24452 25158
rect 24400 25094 24452 25100
rect 24492 24200 24544 24206
rect 24492 24142 24544 24148
rect 24400 24064 24452 24070
rect 24400 24006 24452 24012
rect 24412 23798 24440 24006
rect 24400 23792 24452 23798
rect 24400 23734 24452 23740
rect 24504 23526 24532 24142
rect 24492 23520 24544 23526
rect 24492 23462 24544 23468
rect 24308 21412 24360 21418
rect 24308 21354 24360 21360
rect 23756 19372 23808 19378
rect 23756 19314 23808 19320
rect 23768 19174 23796 19314
rect 23756 19168 23808 19174
rect 23756 19110 23808 19116
rect 23480 11756 23532 11762
rect 23480 11698 23532 11704
rect 23388 10532 23440 10538
rect 23388 10474 23440 10480
rect 23768 10470 23796 19110
rect 24124 14272 24176 14278
rect 24124 14214 24176 14220
rect 24136 14074 24164 14214
rect 24124 14068 24176 14074
rect 24124 14010 24176 14016
rect 23756 10464 23808 10470
rect 23756 10406 23808 10412
rect 24504 6914 24532 23462
rect 24584 22704 24636 22710
rect 24584 22646 24636 22652
rect 24596 18154 24624 22646
rect 24688 22574 24716 46990
rect 24780 46578 24808 49286
rect 25778 49286 26096 49314
rect 25778 49200 25834 49286
rect 24860 47116 24912 47122
rect 24860 47058 24912 47064
rect 24768 46572 24820 46578
rect 24768 46514 24820 46520
rect 24872 39642 24900 47058
rect 26068 47054 26096 49286
rect 26422 49200 26478 50000
rect 27066 49314 27122 50000
rect 27066 49286 27384 49314
rect 27066 49200 27122 49286
rect 26436 47258 26464 49200
rect 27356 47258 27384 49286
rect 27710 49200 27766 50000
rect 28354 49314 28410 50000
rect 28354 49286 28672 49314
rect 28354 49200 28410 49286
rect 26424 47252 26476 47258
rect 26424 47194 26476 47200
rect 27344 47252 27396 47258
rect 27344 47194 27396 47200
rect 27724 47190 27752 49200
rect 26148 47184 26200 47190
rect 26148 47126 26200 47132
rect 27712 47184 27764 47190
rect 27712 47126 27764 47132
rect 26056 47048 26108 47054
rect 26056 46990 26108 46996
rect 25412 46980 25464 46986
rect 25412 46922 25464 46928
rect 24860 39636 24912 39642
rect 24860 39578 24912 39584
rect 24952 37936 25004 37942
rect 24952 37878 25004 37884
rect 24860 35488 24912 35494
rect 24860 35430 24912 35436
rect 24872 35086 24900 35430
rect 24860 35080 24912 35086
rect 24860 35022 24912 35028
rect 24860 30184 24912 30190
rect 24860 30126 24912 30132
rect 24872 29594 24900 30126
rect 24780 29578 24900 29594
rect 24768 29572 24900 29578
rect 24820 29566 24900 29572
rect 24768 29514 24820 29520
rect 24964 26234 24992 37878
rect 25320 28076 25372 28082
rect 25320 28018 25372 28024
rect 24872 26206 24992 26234
rect 24768 24744 24820 24750
rect 24768 24686 24820 24692
rect 24780 24410 24808 24686
rect 24768 24404 24820 24410
rect 24768 24346 24820 24352
rect 24872 24206 24900 26206
rect 25332 25498 25360 28018
rect 25320 25492 25372 25498
rect 25320 25434 25372 25440
rect 25044 25220 25096 25226
rect 25044 25162 25096 25168
rect 25056 24886 25084 25162
rect 25044 24880 25096 24886
rect 25044 24822 25096 24828
rect 25332 24818 25360 25434
rect 25320 24812 25372 24818
rect 25320 24754 25372 24760
rect 25228 24676 25280 24682
rect 25228 24618 25280 24624
rect 24860 24200 24912 24206
rect 24860 24142 24912 24148
rect 24872 23866 24900 24142
rect 25240 24070 25268 24618
rect 25228 24064 25280 24070
rect 25228 24006 25280 24012
rect 24860 23860 24912 23866
rect 24860 23802 24912 23808
rect 24872 23322 24900 23802
rect 24860 23316 24912 23322
rect 24860 23258 24912 23264
rect 24676 22568 24728 22574
rect 24676 22510 24728 22516
rect 24768 22432 24820 22438
rect 24768 22374 24820 22380
rect 24780 21894 24808 22374
rect 24768 21888 24820 21894
rect 24768 21830 24820 21836
rect 24584 18148 24636 18154
rect 24584 18090 24636 18096
rect 24320 6886 24532 6914
rect 23756 5568 23808 5574
rect 23756 5510 23808 5516
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 23204 3392 23256 3398
rect 23204 3334 23256 3340
rect 23664 3392 23716 3398
rect 23664 3334 23716 3340
rect 23216 2990 23244 3334
rect 23204 2984 23256 2990
rect 23204 2926 23256 2932
rect 22284 2508 22336 2514
rect 22284 2450 22336 2456
rect 21928 2378 22048 2394
rect 21916 2372 22048 2378
rect 21968 2366 22048 2372
rect 21916 2314 21968 2320
rect 21928 800 21956 2314
rect 22560 1760 22612 1766
rect 22560 1702 22612 1708
rect 22572 800 22600 1702
rect 23216 800 23244 2926
rect 23676 2378 23704 3334
rect 23768 2650 23796 5510
rect 23756 2644 23808 2650
rect 23756 2586 23808 2592
rect 23848 2576 23900 2582
rect 23848 2518 23900 2524
rect 23664 2372 23716 2378
rect 23664 2314 23716 2320
rect 23676 1766 23704 2314
rect 23664 1760 23716 1766
rect 23664 1702 23716 1708
rect 23860 800 23888 2518
rect 24320 2038 24348 6886
rect 24400 5568 24452 5574
rect 24400 5510 24452 5516
rect 24412 5234 24440 5510
rect 24400 5228 24452 5234
rect 24400 5170 24452 5176
rect 24676 4140 24728 4146
rect 24676 4082 24728 4088
rect 24688 3670 24716 4082
rect 24676 3664 24728 3670
rect 24676 3606 24728 3612
rect 24492 3392 24544 3398
rect 24492 3334 24544 3340
rect 24400 3052 24452 3058
rect 24400 2994 24452 3000
rect 24412 2650 24440 2994
rect 24400 2644 24452 2650
rect 24400 2586 24452 2592
rect 24308 2032 24360 2038
rect 24308 1974 24360 1980
rect 24504 800 24532 3334
rect 24688 2990 24716 3606
rect 24780 3602 24808 21830
rect 24952 6452 25004 6458
rect 24952 6394 25004 6400
rect 24964 5778 24992 6394
rect 24952 5772 25004 5778
rect 24952 5714 25004 5720
rect 25240 4010 25268 24006
rect 25424 5914 25452 46922
rect 26068 46714 26096 46990
rect 26056 46708 26108 46714
rect 26056 46650 26108 46656
rect 26160 43450 26188 47126
rect 26976 47048 27028 47054
rect 26976 46990 27028 46996
rect 27344 47048 27396 47054
rect 27344 46990 27396 46996
rect 27896 47048 27948 47054
rect 27896 46990 27948 46996
rect 26148 43444 26200 43450
rect 26148 43386 26200 43392
rect 26424 43308 26476 43314
rect 26424 43250 26476 43256
rect 26436 42906 26464 43250
rect 26424 42900 26476 42906
rect 26424 42842 26476 42848
rect 26608 42560 26660 42566
rect 26608 42502 26660 42508
rect 26148 42016 26200 42022
rect 26148 41958 26200 41964
rect 26160 41414 26188 41958
rect 25976 41386 26188 41414
rect 25976 28694 26004 41386
rect 26148 33856 26200 33862
rect 26148 33798 26200 33804
rect 26056 30048 26108 30054
rect 26056 29990 26108 29996
rect 26068 29510 26096 29990
rect 26056 29504 26108 29510
rect 26056 29446 26108 29452
rect 25964 28688 26016 28694
rect 25964 28630 26016 28636
rect 25976 28014 26004 28630
rect 26068 28082 26096 29446
rect 26056 28076 26108 28082
rect 26056 28018 26108 28024
rect 25964 28008 26016 28014
rect 26160 27962 26188 33798
rect 25964 27950 26016 27956
rect 26068 27934 26188 27962
rect 26068 18630 26096 27934
rect 26148 27872 26200 27878
rect 26148 27814 26200 27820
rect 26056 18624 26108 18630
rect 26056 18566 26108 18572
rect 26160 16590 26188 27814
rect 26424 26512 26476 26518
rect 26424 26454 26476 26460
rect 26436 26042 26464 26454
rect 26424 26036 26476 26042
rect 26424 25978 26476 25984
rect 26240 25152 26292 25158
rect 26240 25094 26292 25100
rect 26252 23254 26280 25094
rect 26240 23248 26292 23254
rect 26240 23190 26292 23196
rect 26516 18080 26568 18086
rect 26516 18022 26568 18028
rect 26528 17678 26556 18022
rect 26516 17672 26568 17678
rect 26516 17614 26568 17620
rect 26148 16584 26200 16590
rect 26148 16526 26200 16532
rect 26160 16250 26188 16526
rect 26332 16448 26384 16454
rect 26332 16390 26384 16396
rect 26148 16244 26200 16250
rect 26148 16186 26200 16192
rect 25412 5908 25464 5914
rect 25412 5850 25464 5856
rect 25424 5642 25452 5850
rect 25412 5636 25464 5642
rect 25412 5578 25464 5584
rect 25596 5024 25648 5030
rect 25596 4966 25648 4972
rect 25228 4004 25280 4010
rect 25228 3946 25280 3952
rect 24768 3596 24820 3602
rect 24768 3538 24820 3544
rect 24676 2984 24728 2990
rect 24676 2926 24728 2932
rect 25608 2446 25636 4966
rect 25964 3460 26016 3466
rect 25964 3402 26016 3408
rect 25976 3194 26004 3402
rect 25964 3188 26016 3194
rect 25964 3130 26016 3136
rect 26160 2514 26188 16186
rect 26344 15366 26372 16390
rect 26332 15360 26384 15366
rect 26332 15302 26384 15308
rect 26424 14272 26476 14278
rect 26424 14214 26476 14220
rect 26436 14006 26464 14214
rect 26424 14000 26476 14006
rect 26424 13942 26476 13948
rect 26240 13796 26292 13802
rect 26240 13738 26292 13744
rect 26252 4146 26280 13738
rect 26332 5772 26384 5778
rect 26332 5714 26384 5720
rect 26344 5370 26372 5714
rect 26332 5364 26384 5370
rect 26332 5306 26384 5312
rect 26240 4140 26292 4146
rect 26240 4082 26292 4088
rect 26620 3738 26648 42502
rect 26988 41818 27016 46990
rect 27160 46436 27212 46442
rect 27160 46378 27212 46384
rect 27068 43104 27120 43110
rect 27068 43046 27120 43052
rect 27080 42702 27108 43046
rect 27068 42696 27120 42702
rect 27068 42638 27120 42644
rect 27172 42378 27200 46378
rect 27080 42350 27200 42378
rect 27356 42362 27384 46990
rect 27436 46980 27488 46986
rect 27436 46922 27488 46928
rect 27344 42356 27396 42362
rect 26976 41812 27028 41818
rect 26976 41754 27028 41760
rect 26884 35012 26936 35018
rect 26884 34954 26936 34960
rect 26792 23248 26844 23254
rect 26792 23190 26844 23196
rect 26804 22094 26832 23190
rect 26712 22066 26832 22094
rect 26712 14618 26740 22066
rect 26896 17218 26924 34954
rect 27080 32570 27108 42350
rect 27344 42298 27396 42304
rect 27160 42220 27212 42226
rect 27160 42162 27212 42168
rect 27172 41274 27200 42162
rect 27160 41268 27212 41274
rect 27160 41210 27212 41216
rect 27344 41132 27396 41138
rect 27344 41074 27396 41080
rect 27356 35290 27384 41074
rect 27344 35284 27396 35290
rect 27344 35226 27396 35232
rect 27448 34746 27476 46922
rect 27908 46374 27936 46990
rect 28644 46578 28672 49286
rect 28998 49200 29054 50000
rect 29642 49314 29698 50000
rect 29642 49286 29960 49314
rect 29642 49200 29698 49286
rect 29012 47054 29040 49200
rect 29000 47048 29052 47054
rect 29000 46990 29052 46996
rect 29644 47048 29696 47054
rect 29644 46990 29696 46996
rect 29552 46912 29604 46918
rect 29552 46854 29604 46860
rect 28632 46572 28684 46578
rect 28632 46514 28684 46520
rect 29564 46510 29592 46854
rect 29552 46504 29604 46510
rect 29552 46446 29604 46452
rect 27896 46368 27948 46374
rect 27896 46310 27948 46316
rect 28448 46368 28500 46374
rect 28448 46310 28500 46316
rect 27620 38752 27672 38758
rect 27620 38694 27672 38700
rect 27436 34740 27488 34746
rect 27436 34682 27488 34688
rect 27344 34604 27396 34610
rect 27344 34546 27396 34552
rect 27356 34202 27384 34546
rect 27344 34196 27396 34202
rect 27344 34138 27396 34144
rect 27632 33114 27660 38694
rect 27620 33108 27672 33114
rect 27620 33050 27672 33056
rect 27068 32564 27120 32570
rect 27068 32506 27120 32512
rect 27908 32230 27936 46310
rect 27988 43648 28040 43654
rect 27988 43590 28040 43596
rect 28000 43246 28028 43590
rect 27988 43240 28040 43246
rect 27988 43182 28040 43188
rect 28000 42770 28028 43182
rect 27988 42764 28040 42770
rect 27988 42706 28040 42712
rect 28000 42022 28028 42706
rect 27988 42016 28040 42022
rect 27988 41958 28040 41964
rect 28460 35834 28488 46310
rect 29656 46170 29684 46990
rect 29932 46578 29960 49286
rect 30286 49200 30342 50000
rect 30930 49200 30986 50000
rect 31574 49314 31630 50000
rect 31574 49286 31708 49314
rect 31574 49200 31630 49286
rect 30300 47274 30328 49200
rect 30300 47258 30420 47274
rect 30944 47258 30972 49200
rect 31680 47274 31708 49286
rect 32218 49200 32274 50000
rect 32862 49314 32918 50000
rect 33506 49314 33562 50000
rect 34150 49314 34206 50000
rect 32862 49286 32996 49314
rect 32862 49200 32918 49286
rect 31680 47258 31800 47274
rect 30300 47252 30432 47258
rect 30300 47246 30380 47252
rect 30380 47194 30432 47200
rect 30932 47252 30984 47258
rect 31680 47252 31812 47258
rect 31680 47246 31760 47252
rect 30932 47194 30984 47200
rect 31760 47194 31812 47200
rect 30932 47048 30984 47054
rect 30932 46990 30984 46996
rect 31484 47048 31536 47054
rect 31484 46990 31536 46996
rect 29920 46572 29972 46578
rect 29920 46514 29972 46520
rect 30944 46374 30972 46990
rect 31496 46374 31524 46990
rect 32232 46646 32260 49200
rect 32968 47122 32996 49286
rect 33506 49286 33824 49314
rect 33506 49200 33562 49286
rect 32956 47116 33008 47122
rect 32956 47058 33008 47064
rect 32220 46640 32272 46646
rect 32220 46582 32272 46588
rect 31576 46436 31628 46442
rect 31576 46378 31628 46384
rect 30932 46368 30984 46374
rect 30932 46310 30984 46316
rect 31484 46368 31536 46374
rect 31484 46310 31536 46316
rect 29644 46164 29696 46170
rect 29644 46106 29696 46112
rect 30380 45008 30432 45014
rect 30380 44950 30432 44956
rect 30392 43314 30420 44950
rect 30380 43308 30432 43314
rect 30380 43250 30432 43256
rect 28448 35828 28500 35834
rect 28448 35770 28500 35776
rect 29368 32904 29420 32910
rect 29368 32846 29420 32852
rect 29380 32570 29408 32846
rect 29368 32564 29420 32570
rect 29368 32506 29420 32512
rect 28724 32360 28776 32366
rect 28724 32302 28776 32308
rect 29828 32360 29880 32366
rect 29828 32302 29880 32308
rect 27896 32224 27948 32230
rect 27896 32166 27948 32172
rect 28736 31822 28764 32302
rect 28724 31816 28776 31822
rect 28724 31758 28776 31764
rect 27528 30252 27580 30258
rect 27528 30194 27580 30200
rect 26976 30048 27028 30054
rect 26976 29990 27028 29996
rect 26988 29714 27016 29990
rect 27540 29850 27568 30194
rect 27528 29844 27580 29850
rect 27528 29786 27580 29792
rect 26976 29708 27028 29714
rect 26976 29650 27028 29656
rect 27068 29504 27120 29510
rect 27068 29446 27120 29452
rect 27988 29504 28040 29510
rect 27988 29446 28040 29452
rect 27080 29306 27108 29446
rect 27068 29300 27120 29306
rect 27068 29242 27120 29248
rect 26976 29096 27028 29102
rect 26976 29038 27028 29044
rect 26804 17190 26924 17218
rect 26700 14612 26752 14618
rect 26700 14554 26752 14560
rect 26712 13802 26740 14554
rect 26700 13796 26752 13802
rect 26700 13738 26752 13744
rect 26804 11830 26832 17190
rect 26988 17134 27016 29038
rect 27712 26376 27764 26382
rect 27712 26318 27764 26324
rect 27724 26042 27752 26318
rect 27712 26036 27764 26042
rect 27712 25978 27764 25984
rect 27068 25832 27120 25838
rect 27068 25774 27120 25780
rect 27080 25158 27108 25774
rect 27068 25152 27120 25158
rect 27068 25094 27120 25100
rect 27896 24608 27948 24614
rect 27896 24550 27948 24556
rect 27908 24274 27936 24550
rect 27896 24268 27948 24274
rect 27896 24210 27948 24216
rect 27908 23662 27936 24210
rect 27896 23656 27948 23662
rect 27896 23598 27948 23604
rect 27908 23322 27936 23598
rect 27896 23316 27948 23322
rect 27896 23258 27948 23264
rect 26976 17128 27028 17134
rect 26976 17070 27028 17076
rect 26988 15450 27016 17070
rect 27068 16448 27120 16454
rect 27068 16390 27120 16396
rect 27080 16046 27108 16390
rect 27068 16040 27120 16046
rect 27068 15982 27120 15988
rect 26988 15422 27108 15450
rect 26976 15360 27028 15366
rect 26976 15302 27028 15308
rect 26884 13728 26936 13734
rect 26884 13670 26936 13676
rect 26896 13326 26924 13670
rect 26884 13320 26936 13326
rect 26884 13262 26936 13268
rect 26792 11824 26844 11830
rect 26792 11766 26844 11772
rect 26700 5704 26752 5710
rect 26700 5646 26752 5652
rect 26608 3732 26660 3738
rect 26608 3674 26660 3680
rect 26424 3392 26476 3398
rect 26424 3334 26476 3340
rect 26436 3058 26464 3334
rect 26424 3052 26476 3058
rect 26424 2994 26476 3000
rect 26148 2508 26200 2514
rect 26148 2450 26200 2456
rect 25596 2440 25648 2446
rect 25596 2382 25648 2388
rect 25780 2372 25832 2378
rect 25780 2314 25832 2320
rect 24860 2304 24912 2310
rect 24860 2246 24912 2252
rect 24872 1970 24900 2246
rect 24860 1964 24912 1970
rect 24860 1906 24912 1912
rect 25136 1896 25188 1902
rect 25136 1838 25188 1844
rect 25148 800 25176 1838
rect 25792 800 25820 2314
rect 26436 800 26464 2994
rect 26712 2650 26740 5646
rect 26988 3194 27016 15302
rect 27080 15162 27108 15422
rect 27068 15156 27120 15162
rect 27068 15098 27120 15104
rect 27896 14816 27948 14822
rect 27896 14758 27948 14764
rect 27908 14482 27936 14758
rect 27896 14476 27948 14482
rect 27896 14418 27948 14424
rect 27620 14408 27672 14414
rect 27620 14350 27672 14356
rect 27436 13864 27488 13870
rect 27436 13806 27488 13812
rect 27068 5568 27120 5574
rect 27068 5510 27120 5516
rect 27080 5234 27108 5510
rect 27068 5228 27120 5234
rect 27068 5170 27120 5176
rect 27160 3392 27212 3398
rect 27160 3334 27212 3340
rect 26976 3188 27028 3194
rect 26976 3130 27028 3136
rect 27068 2984 27120 2990
rect 27068 2926 27120 2932
rect 26700 2644 26752 2650
rect 26700 2586 26752 2592
rect 27080 800 27108 2926
rect 27172 2446 27200 3334
rect 27448 3194 27476 13806
rect 27632 5846 27660 14350
rect 27620 5840 27672 5846
rect 27620 5782 27672 5788
rect 27620 5704 27672 5710
rect 27620 5646 27672 5652
rect 27528 3392 27580 3398
rect 27528 3334 27580 3340
rect 27436 3188 27488 3194
rect 27436 3130 27488 3136
rect 27540 2990 27568 3334
rect 27528 2984 27580 2990
rect 27528 2926 27580 2932
rect 27632 2650 27660 5646
rect 27712 3528 27764 3534
rect 27712 3470 27764 3476
rect 27620 2644 27672 2650
rect 27620 2586 27672 2592
rect 27160 2440 27212 2446
rect 27160 2382 27212 2388
rect 27172 1902 27200 2382
rect 27724 2378 27752 3470
rect 27804 2848 27856 2854
rect 27804 2790 27856 2796
rect 27816 2650 27844 2790
rect 27804 2644 27856 2650
rect 27804 2586 27856 2592
rect 28000 2514 28028 29446
rect 29460 24200 29512 24206
rect 29460 24142 29512 24148
rect 28540 24064 28592 24070
rect 28540 24006 28592 24012
rect 28552 23118 28580 24006
rect 29472 23866 29500 24142
rect 29460 23860 29512 23866
rect 29460 23802 29512 23808
rect 28540 23112 28592 23118
rect 28540 23054 28592 23060
rect 28356 14952 28408 14958
rect 28356 14894 28408 14900
rect 28368 3194 28396 14894
rect 29736 11892 29788 11898
rect 29736 11834 29788 11840
rect 28908 5024 28960 5030
rect 28908 4966 28960 4972
rect 28920 3398 28948 4966
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 28356 3188 28408 3194
rect 28356 3130 28408 3136
rect 28540 3052 28592 3058
rect 28540 2994 28592 3000
rect 28552 2774 28580 2994
rect 29644 2848 29696 2854
rect 29644 2790 29696 2796
rect 28368 2746 28580 2774
rect 27988 2508 28040 2514
rect 27988 2450 28040 2456
rect 27712 2372 27764 2378
rect 27712 2314 27764 2320
rect 27160 1896 27212 1902
rect 27160 1838 27212 1844
rect 27724 800 27752 2314
rect 28368 800 28396 2746
rect 28448 2644 28500 2650
rect 28448 2586 28500 2592
rect 28460 2310 28488 2586
rect 29656 2446 29684 2790
rect 29748 2582 29776 11834
rect 29840 11626 29868 32302
rect 30380 30252 30432 30258
rect 30380 30194 30432 30200
rect 30392 26314 30420 30194
rect 30944 30054 30972 46310
rect 31496 37126 31524 46310
rect 31588 43450 31616 46378
rect 32232 46170 32260 46582
rect 32588 46368 32640 46374
rect 32588 46310 32640 46316
rect 32220 46164 32272 46170
rect 32220 46106 32272 46112
rect 31576 43444 31628 43450
rect 31576 43386 31628 43392
rect 31484 37120 31536 37126
rect 31484 37062 31536 37068
rect 30932 30048 30984 30054
rect 30932 29990 30984 29996
rect 30380 26308 30432 26314
rect 30380 26250 30432 26256
rect 29920 23520 29972 23526
rect 29920 23462 29972 23468
rect 29828 11620 29880 11626
rect 29828 11562 29880 11568
rect 29736 2576 29788 2582
rect 29736 2518 29788 2524
rect 29644 2440 29696 2446
rect 29644 2382 29696 2388
rect 28448 2304 28500 2310
rect 28448 2246 28500 2252
rect 29656 800 29684 2382
rect 29932 2038 29960 23462
rect 30840 22976 30892 22982
rect 30840 22918 30892 22924
rect 30472 6656 30524 6662
rect 30472 6598 30524 6604
rect 30484 3738 30512 6598
rect 30852 4146 30880 22918
rect 32600 20330 32628 46310
rect 32968 46170 32996 47058
rect 33796 46578 33824 49286
rect 34150 49286 34468 49314
rect 34150 49200 34206 49286
rect 34440 46578 34468 49286
rect 34794 49200 34850 50000
rect 35438 49314 35494 50000
rect 35360 49286 35494 49314
rect 34808 47190 34836 49200
rect 34934 47356 35242 47365
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47291 35242 47300
rect 34796 47184 34848 47190
rect 34716 47144 34796 47172
rect 34520 47048 34572 47054
rect 34520 46990 34572 46996
rect 33784 46572 33836 46578
rect 33784 46514 33836 46520
rect 34428 46572 34480 46578
rect 34428 46514 34480 46520
rect 33600 46368 33652 46374
rect 33600 46310 33652 46316
rect 32956 46164 33008 46170
rect 32956 46106 33008 46112
rect 33612 46102 33640 46310
rect 33796 46170 33824 46514
rect 34440 46170 34468 46514
rect 33784 46164 33836 46170
rect 33784 46106 33836 46112
rect 34428 46164 34480 46170
rect 34428 46106 34480 46112
rect 33600 46096 33652 46102
rect 33600 46038 33652 46044
rect 33600 44940 33652 44946
rect 33600 44882 33652 44888
rect 33612 44198 33640 44882
rect 33600 44192 33652 44198
rect 33600 44134 33652 44140
rect 33612 29102 33640 44134
rect 34244 29640 34296 29646
rect 34244 29582 34296 29588
rect 34256 29306 34284 29582
rect 34244 29300 34296 29306
rect 34244 29242 34296 29248
rect 33600 29096 33652 29102
rect 33600 29038 33652 29044
rect 32956 29028 33008 29034
rect 32956 28970 33008 28976
rect 32968 24177 32996 28970
rect 33612 28762 33640 29038
rect 33416 28756 33468 28762
rect 33416 28698 33468 28704
rect 33600 28756 33652 28762
rect 33600 28698 33652 28704
rect 33428 24750 33456 28698
rect 33416 24744 33468 24750
rect 33416 24686 33468 24692
rect 32954 24168 33010 24177
rect 32954 24103 33010 24112
rect 33428 20602 33456 24686
rect 33416 20596 33468 20602
rect 33416 20538 33468 20544
rect 32588 20324 32640 20330
rect 32588 20266 32640 20272
rect 33428 19922 33456 20538
rect 33784 20392 33836 20398
rect 33784 20334 33836 20340
rect 33140 19916 33192 19922
rect 33140 19858 33192 19864
rect 33416 19916 33468 19922
rect 33416 19858 33468 19864
rect 33152 19310 33180 19858
rect 33796 19514 33824 20334
rect 34244 19712 34296 19718
rect 34244 19654 34296 19660
rect 33784 19508 33836 19514
rect 33784 19450 33836 19456
rect 34256 19378 34284 19654
rect 34244 19372 34296 19378
rect 34244 19314 34296 19320
rect 33140 19304 33192 19310
rect 33140 19246 33192 19252
rect 33324 19304 33376 19310
rect 33324 19246 33376 19252
rect 33152 18970 33180 19246
rect 33140 18964 33192 18970
rect 33140 18906 33192 18912
rect 33336 18630 33364 19246
rect 33324 18624 33376 18630
rect 33324 18566 33376 18572
rect 30932 9376 30984 9382
rect 30932 9318 30984 9324
rect 30944 6914 30972 9318
rect 31024 7880 31076 7886
rect 31024 7822 31076 7828
rect 31036 7274 31064 7822
rect 31024 7268 31076 7274
rect 31024 7210 31076 7216
rect 30944 6886 31064 6914
rect 30840 4140 30892 4146
rect 30840 4082 30892 4088
rect 30472 3732 30524 3738
rect 30472 3674 30524 3680
rect 30484 2990 30512 3674
rect 30472 2984 30524 2990
rect 30472 2926 30524 2932
rect 30852 2446 30880 4082
rect 31036 3738 31064 6886
rect 31024 3732 31076 3738
rect 31024 3674 31076 3680
rect 33336 3670 33364 18566
rect 33784 18148 33836 18154
rect 33784 18090 33836 18096
rect 33796 9042 33824 18090
rect 33876 17536 33928 17542
rect 33876 17478 33928 17484
rect 33784 9036 33836 9042
rect 33784 8978 33836 8984
rect 33888 3738 33916 17478
rect 34428 14272 34480 14278
rect 34428 14214 34480 14220
rect 34440 13870 34468 14214
rect 34532 14074 34560 46990
rect 34612 45892 34664 45898
rect 34612 45834 34664 45840
rect 34624 29850 34652 45834
rect 34716 45558 34744 47144
rect 34796 47126 34848 47132
rect 34796 46572 34848 46578
rect 34796 46514 34848 46520
rect 34704 45552 34756 45558
rect 34704 45494 34756 45500
rect 34808 45286 34836 46514
rect 34934 46268 35242 46277
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46203 35242 46212
rect 35256 46028 35308 46034
rect 35256 45970 35308 45976
rect 35268 45490 35296 45970
rect 35360 45966 35388 49286
rect 35438 49200 35494 49286
rect 36082 49314 36138 50000
rect 36726 49314 36782 50000
rect 36082 49286 36400 49314
rect 36082 49200 36138 49286
rect 35438 49056 35494 49065
rect 35438 48991 35494 49000
rect 35452 46714 35480 48991
rect 35806 48376 35862 48385
rect 35806 48311 35862 48320
rect 35714 47696 35770 47705
rect 35714 47631 35770 47640
rect 35624 47116 35676 47122
rect 35624 47058 35676 47064
rect 35440 46708 35492 46714
rect 35440 46650 35492 46656
rect 35532 46504 35584 46510
rect 35532 46446 35584 46452
rect 35440 46436 35492 46442
rect 35440 46378 35492 46384
rect 35348 45960 35400 45966
rect 35348 45902 35400 45908
rect 35360 45626 35388 45902
rect 35348 45620 35400 45626
rect 35348 45562 35400 45568
rect 35256 45484 35308 45490
rect 35256 45426 35308 45432
rect 34796 45280 34848 45286
rect 34796 45222 34848 45228
rect 34704 44736 34756 44742
rect 34704 44678 34756 44684
rect 34716 43790 34744 44678
rect 34704 43784 34756 43790
rect 34704 43726 34756 43732
rect 34612 29844 34664 29850
rect 34612 29786 34664 29792
rect 34612 15020 34664 15026
rect 34612 14962 34664 14968
rect 34520 14068 34572 14074
rect 34520 14010 34572 14016
rect 34428 13864 34480 13870
rect 34428 13806 34480 13812
rect 33968 13728 34020 13734
rect 33968 13670 34020 13676
rect 33980 13326 34008 13670
rect 34440 13394 34468 13806
rect 34624 13530 34652 14962
rect 34612 13524 34664 13530
rect 34612 13466 34664 13472
rect 34428 13388 34480 13394
rect 34428 13330 34480 13336
rect 33968 13320 34020 13326
rect 33968 13262 34020 13268
rect 34440 12646 34468 13330
rect 34612 13184 34664 13190
rect 34612 13126 34664 13132
rect 34428 12640 34480 12646
rect 34428 12582 34480 12588
rect 34440 12442 34468 12582
rect 34428 12436 34480 12442
rect 34428 12378 34480 12384
rect 33876 3732 33928 3738
rect 33876 3674 33928 3680
rect 33324 3664 33376 3670
rect 33324 3606 33376 3612
rect 30932 3528 30984 3534
rect 30932 3470 30984 3476
rect 30012 2440 30064 2446
rect 30012 2382 30064 2388
rect 30840 2440 30892 2446
rect 30840 2382 30892 2388
rect 30024 2106 30052 2382
rect 30288 2304 30340 2310
rect 30288 2246 30340 2252
rect 30012 2100 30064 2106
rect 30012 2042 30064 2048
rect 29920 2032 29972 2038
rect 29920 1974 29972 1980
rect 30300 800 30328 2246
rect 30944 800 30972 3470
rect 32036 3392 32088 3398
rect 32036 3334 32088 3340
rect 32220 3392 32272 3398
rect 32220 3334 32272 3340
rect 32772 3392 32824 3398
rect 32772 3334 32824 3340
rect 32864 3392 32916 3398
rect 32864 3334 32916 3340
rect 31668 3188 31720 3194
rect 31496 3148 31668 3176
rect 31496 1970 31524 3148
rect 31668 3130 31720 3136
rect 32048 3126 32076 3334
rect 32036 3120 32088 3126
rect 32036 3062 32088 3068
rect 32232 2446 32260 3334
rect 32784 3058 32812 3334
rect 32312 3052 32364 3058
rect 32312 2994 32364 3000
rect 32772 3052 32824 3058
rect 32772 2994 32824 3000
rect 31760 2440 31812 2446
rect 31588 2400 31760 2428
rect 31484 1964 31536 1970
rect 31484 1906 31536 1912
rect 31588 800 31616 2400
rect 31760 2382 31812 2388
rect 32220 2440 32272 2446
rect 32220 2382 32272 2388
rect 32324 2258 32352 2994
rect 32876 2990 32904 3334
rect 32864 2984 32916 2990
rect 32864 2926 32916 2932
rect 32232 2230 32352 2258
rect 32232 800 32260 2230
rect 32876 800 32904 2926
rect 33888 2446 33916 3674
rect 34152 3392 34204 3398
rect 34152 3334 34204 3340
rect 34164 3058 34192 3334
rect 34624 3194 34652 13126
rect 34808 4486 34836 45222
rect 34934 45180 35242 45189
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45115 35242 45124
rect 34934 44092 35242 44101
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44027 35242 44036
rect 35348 43648 35400 43654
rect 35348 43590 35400 43596
rect 34934 43004 35242 43013
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42939 35242 42948
rect 34934 41916 35242 41925
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41851 35242 41860
rect 34934 40828 35242 40837
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40763 35242 40772
rect 34934 39740 35242 39749
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39675 35242 39684
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 35360 37874 35388 43590
rect 35348 37868 35400 37874
rect 35348 37810 35400 37816
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35452 25294 35480 46378
rect 35544 46034 35572 46446
rect 35532 46028 35584 46034
rect 35532 45970 35584 45976
rect 35636 45948 35664 47058
rect 35728 46102 35756 47631
rect 35820 46170 35848 48311
rect 36084 47048 36136 47054
rect 36084 46990 36136 46996
rect 35900 46572 35952 46578
rect 35900 46514 35952 46520
rect 35912 46345 35940 46514
rect 35898 46336 35954 46345
rect 35898 46271 35954 46280
rect 35808 46164 35860 46170
rect 35808 46106 35860 46112
rect 35716 46096 35768 46102
rect 35716 46038 35768 46044
rect 35636 45920 35756 45948
rect 35624 45824 35676 45830
rect 35624 45766 35676 45772
rect 35532 44192 35584 44198
rect 35532 44134 35584 44140
rect 35544 43382 35572 44134
rect 35532 43376 35584 43382
rect 35532 43318 35584 43324
rect 35636 42634 35664 45766
rect 35624 42628 35676 42634
rect 35624 42570 35676 42576
rect 35728 41274 35756 45920
rect 35912 45082 35940 46271
rect 35992 45960 36044 45966
rect 35992 45902 36044 45908
rect 36004 45354 36032 45902
rect 35992 45348 36044 45354
rect 35992 45290 36044 45296
rect 35900 45076 35952 45082
rect 35900 45018 35952 45024
rect 36096 44198 36124 46990
rect 36372 46918 36400 49286
rect 36648 49286 36782 49314
rect 36648 47258 36676 49286
rect 36726 49200 36782 49286
rect 37370 49200 37426 50000
rect 38014 49314 38070 50000
rect 38658 49314 38714 50000
rect 37476 49286 38070 49314
rect 36636 47252 36688 47258
rect 36636 47194 36688 47200
rect 36360 46912 36412 46918
rect 36360 46854 36412 46860
rect 37280 46912 37332 46918
rect 37280 46854 37332 46860
rect 36268 46572 36320 46578
rect 36268 46514 36320 46520
rect 36280 44198 36308 46514
rect 37186 45656 37242 45665
rect 37186 45591 37242 45600
rect 36820 45484 36872 45490
rect 36820 45426 36872 45432
rect 36832 45370 36860 45426
rect 36740 45342 36860 45370
rect 36544 45280 36596 45286
rect 36544 45222 36596 45228
rect 36556 44878 36584 45222
rect 36544 44872 36596 44878
rect 36544 44814 36596 44820
rect 36084 44192 36136 44198
rect 36084 44134 36136 44140
rect 36268 44192 36320 44198
rect 36268 44134 36320 44140
rect 35716 41268 35768 41274
rect 35716 41210 35768 41216
rect 35992 36168 36044 36174
rect 35992 36110 36044 36116
rect 36004 33114 36032 36110
rect 35992 33108 36044 33114
rect 35992 33050 36044 33056
rect 35440 25288 35492 25294
rect 35440 25230 35492 25236
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 36280 20466 36308 44134
rect 36740 43654 36768 45342
rect 37200 44878 37228 45591
rect 37188 44872 37240 44878
rect 37188 44814 37240 44820
rect 37292 44282 37320 46854
rect 37384 46714 37412 49200
rect 37476 46714 37504 49286
rect 38014 49200 38070 49286
rect 38120 49286 38714 49314
rect 38120 47138 38148 49286
rect 38658 49200 38714 49286
rect 39302 49200 39358 50000
rect 37568 47110 38148 47138
rect 37372 46708 37424 46714
rect 37372 46650 37424 46656
rect 37464 46708 37516 46714
rect 37464 46650 37516 46656
rect 37568 46594 37596 47110
rect 38106 47016 38162 47025
rect 38106 46951 38162 46960
rect 37648 46912 37700 46918
rect 37648 46854 37700 46860
rect 37384 46566 37596 46594
rect 37384 45558 37412 46566
rect 37464 46504 37516 46510
rect 37464 46446 37516 46452
rect 37372 45552 37424 45558
rect 37372 45494 37424 45500
rect 37292 44254 37412 44282
rect 37280 44192 37332 44198
rect 37280 44134 37332 44140
rect 37292 43790 37320 44134
rect 37384 43994 37412 44254
rect 37372 43988 37424 43994
rect 37372 43930 37424 43936
rect 37280 43784 37332 43790
rect 37280 43726 37332 43732
rect 36728 43648 36780 43654
rect 37292 43625 37320 43726
rect 36728 43590 36780 43596
rect 37278 43616 37334 43625
rect 36544 32768 36596 32774
rect 36544 32710 36596 32716
rect 36556 24410 36584 32710
rect 36740 29714 36768 43590
rect 37278 43551 37334 43560
rect 37372 42696 37424 42702
rect 37372 42638 37424 42644
rect 37384 41818 37412 42638
rect 37372 41812 37424 41818
rect 37372 41754 37424 41760
rect 36912 34740 36964 34746
rect 36912 34682 36964 34688
rect 36924 33930 36952 34682
rect 36912 33924 36964 33930
rect 36912 33866 36964 33872
rect 37372 31204 37424 31210
rect 37372 31146 37424 31152
rect 36728 29708 36780 29714
rect 36728 29650 36780 29656
rect 36636 29028 36688 29034
rect 36636 28970 36688 28976
rect 36648 25770 36676 28970
rect 37280 27328 37332 27334
rect 37280 27270 37332 27276
rect 37292 26790 37320 27270
rect 37280 26784 37332 26790
rect 37280 26726 37332 26732
rect 36636 25764 36688 25770
rect 36636 25706 36688 25712
rect 36544 24404 36596 24410
rect 36544 24346 36596 24352
rect 37384 23866 37412 31146
rect 37476 31142 37504 46446
rect 37660 46034 37688 46854
rect 37648 46028 37700 46034
rect 37648 45970 37700 45976
rect 37556 45960 37608 45966
rect 37556 45902 37608 45908
rect 37464 31136 37516 31142
rect 37464 31078 37516 31084
rect 37568 29102 37596 45902
rect 37660 44810 37688 45970
rect 38016 45280 38068 45286
rect 38016 45222 38068 45228
rect 38028 44985 38056 45222
rect 38014 44976 38070 44985
rect 38120 44946 38148 46951
rect 39316 46918 39344 49200
rect 39304 46912 39356 46918
rect 39304 46854 39356 46860
rect 38014 44911 38070 44920
rect 38108 44940 38160 44946
rect 38108 44882 38160 44888
rect 37648 44804 37700 44810
rect 37648 44746 37700 44752
rect 38200 44736 38252 44742
rect 38200 44678 38252 44684
rect 38014 44296 38070 44305
rect 38014 44231 38016 44240
rect 38068 44231 38070 44240
rect 38016 44202 38068 44208
rect 38016 43308 38068 43314
rect 38016 43250 38068 43256
rect 37648 43172 37700 43178
rect 37648 43114 37700 43120
rect 37556 29096 37608 29102
rect 37556 29038 37608 29044
rect 37556 27872 37608 27878
rect 37556 27814 37608 27820
rect 37372 23860 37424 23866
rect 37372 23802 37424 23808
rect 37372 22228 37424 22234
rect 37372 22170 37424 22176
rect 37280 21412 37332 21418
rect 37280 21354 37332 21360
rect 37292 21010 37320 21354
rect 37280 21004 37332 21010
rect 37280 20946 37332 20952
rect 36268 20460 36320 20466
rect 36268 20402 36320 20408
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35440 19848 35492 19854
rect 35440 19790 35492 19796
rect 35348 19168 35400 19174
rect 35348 19110 35400 19116
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35360 18766 35388 19110
rect 35348 18760 35400 18766
rect 35348 18702 35400 18708
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35452 16454 35480 19790
rect 37280 17536 37332 17542
rect 37280 17478 37332 17484
rect 35808 17332 35860 17338
rect 35808 17274 35860 17280
rect 35440 16448 35492 16454
rect 35440 16390 35492 16396
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 35072 13320 35124 13326
rect 35348 13320 35400 13326
rect 35124 13268 35348 13274
rect 35072 13262 35400 13268
rect 34980 13252 35032 13258
rect 35084 13246 35388 13262
rect 34980 13194 35032 13200
rect 34992 13138 35020 13194
rect 35348 13184 35400 13190
rect 34992 13132 35348 13138
rect 34992 13126 35400 13132
rect 34992 13110 35388 13126
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34796 4480 34848 4486
rect 34796 4422 34848 4428
rect 35716 4480 35768 4486
rect 35716 4422 35768 4428
rect 35440 3936 35492 3942
rect 35440 3878 35492 3884
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34612 3188 34664 3194
rect 34612 3130 34664 3136
rect 35452 3058 35480 3878
rect 34152 3052 34204 3058
rect 34152 2994 34204 3000
rect 35440 3052 35492 3058
rect 35440 2994 35492 3000
rect 33876 2440 33928 2446
rect 33876 2382 33928 2388
rect 33508 2304 33560 2310
rect 33508 2246 33560 2252
rect 33520 800 33548 2246
rect 34164 800 34192 2994
rect 34796 2916 34848 2922
rect 34796 2858 34848 2864
rect 34520 2848 34572 2854
rect 34520 2790 34572 2796
rect 34532 2650 34560 2790
rect 34520 2644 34572 2650
rect 34520 2586 34572 2592
rect 34808 2446 34836 2858
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 34796 2304 34848 2310
rect 34796 2246 34848 2252
rect 35164 2304 35216 2310
rect 35164 2246 35216 2252
rect 34808 800 34836 2246
rect 35176 2038 35204 2246
rect 35164 2032 35216 2038
rect 35164 1974 35216 1980
rect 35452 800 35480 2994
rect 35728 2514 35756 4422
rect 35820 2650 35848 17274
rect 37292 17134 37320 17478
rect 37280 17128 37332 17134
rect 37280 17070 37332 17076
rect 37188 16584 37240 16590
rect 37188 16526 37240 16532
rect 37200 16425 37228 16526
rect 37186 16416 37242 16425
rect 37186 16351 37242 16360
rect 37384 16250 37412 22170
rect 37372 16244 37424 16250
rect 37372 16186 37424 16192
rect 36820 13932 36872 13938
rect 36820 13874 36872 13880
rect 36832 13326 36860 13874
rect 36820 13320 36872 13326
rect 36820 13262 36872 13268
rect 37280 12096 37332 12102
rect 37280 12038 37332 12044
rect 37096 11824 37148 11830
rect 37096 11766 37148 11772
rect 36176 7812 36228 7818
rect 36176 7754 36228 7760
rect 36188 4826 36216 7754
rect 36636 5024 36688 5030
rect 36636 4966 36688 4972
rect 36176 4820 36228 4826
rect 36176 4762 36228 4768
rect 36084 3936 36136 3942
rect 36084 3878 36136 3884
rect 36096 3534 36124 3878
rect 36084 3528 36136 3534
rect 36084 3470 36136 3476
rect 35900 2848 35952 2854
rect 35900 2790 35952 2796
rect 35808 2644 35860 2650
rect 35808 2586 35860 2592
rect 35716 2508 35768 2514
rect 35716 2450 35768 2456
rect 35912 1465 35940 2790
rect 35898 1456 35954 1465
rect 35898 1391 35954 1400
rect 36096 800 36124 3470
rect 36188 3126 36216 4762
rect 36452 3936 36504 3942
rect 36452 3878 36504 3884
rect 36176 3120 36228 3126
rect 36176 3062 36228 3068
rect 36464 2378 36492 3878
rect 36544 3596 36596 3602
rect 36544 3538 36596 3544
rect 36556 3194 36584 3538
rect 36544 3188 36596 3194
rect 36544 3130 36596 3136
rect 36648 2446 36676 4966
rect 36728 4480 36780 4486
rect 36728 4422 36780 4428
rect 36740 2990 36768 4422
rect 37108 4146 37136 11766
rect 37292 11694 37320 12038
rect 37280 11688 37332 11694
rect 37278 11656 37280 11665
rect 37332 11656 37334 11665
rect 37278 11591 37334 11600
rect 37280 10600 37332 10606
rect 37280 10542 37332 10548
rect 37292 6458 37320 10542
rect 37568 10266 37596 27814
rect 37660 24274 37688 43114
rect 38028 42945 38056 43250
rect 38014 42936 38070 42945
rect 38014 42871 38070 42880
rect 38108 42696 38160 42702
rect 38108 42638 38160 42644
rect 37832 42560 37884 42566
rect 37832 42502 37884 42508
rect 37740 38208 37792 38214
rect 37740 38150 37792 38156
rect 37648 24268 37700 24274
rect 37648 24210 37700 24216
rect 37648 17536 37700 17542
rect 37648 17478 37700 17484
rect 37660 17338 37688 17478
rect 37752 17338 37780 38150
rect 37844 33998 37872 42502
rect 38120 42265 38148 42638
rect 38106 42256 38162 42265
rect 38106 42191 38162 42200
rect 38108 41608 38160 41614
rect 38106 41576 38108 41585
rect 38160 41576 38162 41585
rect 38106 41511 38162 41520
rect 38108 41132 38160 41138
rect 38108 41074 38160 41080
rect 38120 40905 38148 41074
rect 38106 40896 38162 40905
rect 38106 40831 38162 40840
rect 38108 40520 38160 40526
rect 38108 40462 38160 40468
rect 38120 40225 38148 40462
rect 38106 40216 38162 40225
rect 38106 40151 38162 40160
rect 38016 39840 38068 39846
rect 38016 39782 38068 39788
rect 38028 39545 38056 39782
rect 38014 39536 38070 39545
rect 38014 39471 38070 39480
rect 38014 38856 38070 38865
rect 38014 38791 38016 38800
rect 38068 38791 38070 38800
rect 38016 38762 38068 38768
rect 38108 38344 38160 38350
rect 38108 38286 38160 38292
rect 38120 38185 38148 38286
rect 38106 38176 38162 38185
rect 38106 38111 38162 38120
rect 38016 37664 38068 37670
rect 38016 37606 38068 37612
rect 38028 37505 38056 37606
rect 38014 37496 38070 37505
rect 38014 37431 38070 37440
rect 38108 37256 38160 37262
rect 38108 37198 38160 37204
rect 38120 36854 38148 37198
rect 38108 36848 38160 36854
rect 38106 36816 38108 36825
rect 38160 36816 38162 36825
rect 38106 36751 38162 36760
rect 38014 36136 38070 36145
rect 38014 36071 38070 36080
rect 38028 36038 38056 36071
rect 38016 36032 38068 36038
rect 38016 35974 38068 35980
rect 38108 35692 38160 35698
rect 38108 35634 38160 35640
rect 37924 35488 37976 35494
rect 38120 35465 38148 35634
rect 37924 35430 37976 35436
rect 38106 35456 38162 35465
rect 37832 33992 37884 33998
rect 37832 33934 37884 33940
rect 37936 30122 37964 35430
rect 38106 35391 38162 35400
rect 38108 34604 38160 34610
rect 38108 34546 38160 34552
rect 38120 34105 38148 34546
rect 38106 34096 38162 34105
rect 38106 34031 38162 34040
rect 38108 33516 38160 33522
rect 38108 33458 38160 33464
rect 38120 33425 38148 33458
rect 38106 33416 38162 33425
rect 38106 33351 38162 33360
rect 38108 32904 38160 32910
rect 38108 32846 38160 32852
rect 38120 32745 38148 32846
rect 38106 32736 38162 32745
rect 38106 32671 38162 32680
rect 38108 32428 38160 32434
rect 38108 32370 38160 32376
rect 38120 32065 38148 32370
rect 38106 32056 38162 32065
rect 38106 31991 38162 32000
rect 38016 31816 38068 31822
rect 38016 31758 38068 31764
rect 38028 31385 38056 31758
rect 38014 31376 38070 31385
rect 38014 31311 38070 31320
rect 37924 30116 37976 30122
rect 37924 30058 37976 30064
rect 38016 30048 38068 30054
rect 38014 30016 38016 30025
rect 38068 30016 38070 30025
rect 38014 29951 38070 29960
rect 38108 29640 38160 29646
rect 38108 29582 38160 29588
rect 37924 29504 37976 29510
rect 37924 29446 37976 29452
rect 37936 29238 37964 29446
rect 38120 29345 38148 29582
rect 38106 29336 38162 29345
rect 38106 29271 38162 29280
rect 37924 29232 37976 29238
rect 37924 29174 37976 29180
rect 38108 29164 38160 29170
rect 38108 29106 38160 29112
rect 38120 28665 38148 29106
rect 38106 28656 38162 28665
rect 38106 28591 38162 28600
rect 38014 27976 38070 27985
rect 38014 27911 38016 27920
rect 38068 27911 38070 27920
rect 38016 27882 38068 27888
rect 38016 27328 38068 27334
rect 38014 27296 38016 27305
rect 38068 27296 38070 27305
rect 38014 27231 38070 27240
rect 38108 26988 38160 26994
rect 38108 26930 38160 26936
rect 37924 26784 37976 26790
rect 37924 26726 37976 26732
rect 37936 26450 37964 26726
rect 38120 26625 38148 26930
rect 38106 26616 38162 26625
rect 38106 26551 38162 26560
rect 38016 26512 38068 26518
rect 38016 26454 38068 26460
rect 37924 26444 37976 26450
rect 37924 26386 37976 26392
rect 38028 25945 38056 26454
rect 38014 25936 38070 25945
rect 38014 25871 38070 25880
rect 37924 25832 37976 25838
rect 37924 25774 37976 25780
rect 37936 25498 37964 25774
rect 37924 25492 37976 25498
rect 37924 25434 37976 25440
rect 38108 25288 38160 25294
rect 38106 25256 38108 25265
rect 38160 25256 38162 25265
rect 38106 25191 38162 25200
rect 37832 25152 37884 25158
rect 37832 25094 37884 25100
rect 37844 21146 37872 25094
rect 38108 24812 38160 24818
rect 38108 24754 38160 24760
rect 38120 24585 38148 24754
rect 38106 24576 38162 24585
rect 38106 24511 38162 24520
rect 38016 24064 38068 24070
rect 38016 24006 38068 24012
rect 38028 23905 38056 24006
rect 38014 23896 38070 23905
rect 38014 23831 38070 23840
rect 38016 23520 38068 23526
rect 38016 23462 38068 23468
rect 38028 23225 38056 23462
rect 38014 23216 38070 23225
rect 38014 23151 38070 23160
rect 38108 22976 38160 22982
rect 38108 22918 38160 22924
rect 38120 22574 38148 22918
rect 38108 22568 38160 22574
rect 38106 22536 38108 22545
rect 38160 22536 38162 22545
rect 38106 22471 38162 22480
rect 38108 22024 38160 22030
rect 38108 21966 38160 21972
rect 38120 21865 38148 21966
rect 38106 21856 38162 21865
rect 38106 21791 38162 21800
rect 37924 21548 37976 21554
rect 37924 21490 37976 21496
rect 37832 21140 37884 21146
rect 37832 21082 37884 21088
rect 37832 21004 37884 21010
rect 37832 20946 37884 20952
rect 37648 17332 37700 17338
rect 37648 17274 37700 17280
rect 37740 17332 37792 17338
rect 37740 17274 37792 17280
rect 37648 17196 37700 17202
rect 37648 17138 37700 17144
rect 37660 12850 37688 17138
rect 37740 16448 37792 16454
rect 37740 16390 37792 16396
rect 37648 12844 37700 12850
rect 37648 12786 37700 12792
rect 37648 11756 37700 11762
rect 37648 11698 37700 11704
rect 37556 10260 37608 10266
rect 37556 10202 37608 10208
rect 37280 6452 37332 6458
rect 37280 6394 37332 6400
rect 37372 5568 37424 5574
rect 37372 5510 37424 5516
rect 37384 4214 37412 5510
rect 37660 4758 37688 11698
rect 37752 5234 37780 16390
rect 37844 14482 37872 20946
rect 37936 15450 37964 21490
rect 38016 21344 38068 21350
rect 38016 21286 38068 21292
rect 38028 21185 38056 21286
rect 38014 21176 38070 21185
rect 38014 21111 38070 21120
rect 38108 20936 38160 20942
rect 38108 20878 38160 20884
rect 38120 20505 38148 20878
rect 38106 20496 38162 20505
rect 38106 20431 38162 20440
rect 38014 19816 38070 19825
rect 38014 19751 38070 19760
rect 38028 19718 38056 19751
rect 38016 19712 38068 19718
rect 38016 19654 38068 19660
rect 38016 18624 38068 18630
rect 38016 18566 38068 18572
rect 38028 18465 38056 18566
rect 38014 18456 38070 18465
rect 38014 18391 38070 18400
rect 38108 18284 38160 18290
rect 38108 18226 38160 18232
rect 38120 17785 38148 18226
rect 38106 17776 38162 17785
rect 38106 17711 38162 17720
rect 38108 17672 38160 17678
rect 38108 17614 38160 17620
rect 38120 17105 38148 17614
rect 38106 17096 38162 17105
rect 38106 17031 38162 17040
rect 38016 16992 38068 16998
rect 38016 16934 38068 16940
rect 38028 16590 38056 16934
rect 38016 16584 38068 16590
rect 38016 16526 38068 16532
rect 38016 15904 38068 15910
rect 38016 15846 38068 15852
rect 38028 15745 38056 15846
rect 38014 15736 38070 15745
rect 38014 15671 38070 15680
rect 38108 15496 38160 15502
rect 37936 15422 38056 15450
rect 38108 15438 38160 15444
rect 37924 15360 37976 15366
rect 37924 15302 37976 15308
rect 37936 15094 37964 15302
rect 38028 15162 38056 15422
rect 38016 15156 38068 15162
rect 38016 15098 38068 15104
rect 37924 15088 37976 15094
rect 38120 15065 38148 15438
rect 37924 15030 37976 15036
rect 38106 15056 38162 15065
rect 38106 14991 38162 15000
rect 38108 14816 38160 14822
rect 38108 14758 38160 14764
rect 37832 14476 37884 14482
rect 37832 14418 37884 14424
rect 38120 14414 38148 14758
rect 38108 14408 38160 14414
rect 38106 14376 38108 14385
rect 38160 14376 38162 14385
rect 38106 14311 38162 14320
rect 38016 13728 38068 13734
rect 38014 13696 38016 13705
rect 38068 13696 38070 13705
rect 38014 13631 38070 13640
rect 37924 13252 37976 13258
rect 37924 13194 37976 13200
rect 37832 13184 37884 13190
rect 37832 13126 37884 13132
rect 37844 5710 37872 13126
rect 37936 11354 37964 13194
rect 38016 13184 38068 13190
rect 38016 13126 38068 13132
rect 38028 13025 38056 13126
rect 38014 13016 38070 13025
rect 38014 12951 38070 12960
rect 38108 12776 38160 12782
rect 38108 12718 38160 12724
rect 38120 12374 38148 12718
rect 38108 12368 38160 12374
rect 38106 12336 38108 12345
rect 38160 12336 38162 12345
rect 38106 12271 38162 12280
rect 37924 11348 37976 11354
rect 37924 11290 37976 11296
rect 38108 11144 38160 11150
rect 38108 11086 38160 11092
rect 38120 10985 38148 11086
rect 38106 10976 38162 10985
rect 38106 10911 38162 10920
rect 38108 10668 38160 10674
rect 38108 10610 38160 10616
rect 38120 10305 38148 10610
rect 38106 10296 38162 10305
rect 38106 10231 38162 10240
rect 38108 10056 38160 10062
rect 38108 9998 38160 10004
rect 38120 9625 38148 9998
rect 38106 9616 38162 9625
rect 38106 9551 38162 9560
rect 38108 9376 38160 9382
rect 38108 9318 38160 9324
rect 38120 8974 38148 9318
rect 38108 8968 38160 8974
rect 38106 8936 38108 8945
rect 38160 8936 38162 8945
rect 38106 8871 38162 8880
rect 38016 8356 38068 8362
rect 38016 8298 38068 8304
rect 38028 8265 38056 8298
rect 38014 8256 38070 8265
rect 38014 8191 38070 8200
rect 38016 7744 38068 7750
rect 38016 7686 38068 7692
rect 38028 7585 38056 7686
rect 38014 7576 38070 7585
rect 38014 7511 38070 7520
rect 38016 7404 38068 7410
rect 38016 7346 38068 7352
rect 38028 6905 38056 7346
rect 38014 6896 38070 6905
rect 38014 6831 38070 6840
rect 38014 6216 38070 6225
rect 38014 6151 38016 6160
rect 38068 6151 38070 6160
rect 38016 6122 38068 6128
rect 37832 5704 37884 5710
rect 37832 5646 37884 5652
rect 38212 5642 38240 44678
rect 38292 40044 38344 40050
rect 38292 39986 38344 39992
rect 38304 14006 38332 39986
rect 38384 31884 38436 31890
rect 38384 31826 38436 31832
rect 38292 14000 38344 14006
rect 38292 13942 38344 13948
rect 38396 6254 38424 31826
rect 38568 26376 38620 26382
rect 38568 26318 38620 26324
rect 38476 16040 38528 16046
rect 38476 15982 38528 15988
rect 38384 6248 38436 6254
rect 38384 6190 38436 6196
rect 38200 5636 38252 5642
rect 38200 5578 38252 5584
rect 38016 5568 38068 5574
rect 38014 5536 38016 5545
rect 38068 5536 38070 5545
rect 38014 5471 38070 5480
rect 38488 5370 38516 15982
rect 38580 14890 38608 26318
rect 38568 14884 38620 14890
rect 38568 14826 38620 14832
rect 37832 5364 37884 5370
rect 37832 5306 37884 5312
rect 38476 5364 38528 5370
rect 38476 5306 38528 5312
rect 37740 5228 37792 5234
rect 37740 5170 37792 5176
rect 37648 4752 37700 4758
rect 37648 4694 37700 4700
rect 37372 4208 37424 4214
rect 37372 4150 37424 4156
rect 37096 4140 37148 4146
rect 37096 4082 37148 4088
rect 37108 3534 37136 4082
rect 37844 3534 37872 5306
rect 38016 5024 38068 5030
rect 38016 4966 38068 4972
rect 38028 4865 38056 4966
rect 38014 4856 38070 4865
rect 38014 4791 38070 4800
rect 38016 4548 38068 4554
rect 38016 4490 38068 4496
rect 38028 4185 38056 4490
rect 39304 4208 39356 4214
rect 38014 4176 38070 4185
rect 39304 4150 39356 4156
rect 38014 4111 38070 4120
rect 38660 3664 38712 3670
rect 38660 3606 38712 3612
rect 37096 3528 37148 3534
rect 37096 3470 37148 3476
rect 37832 3528 37884 3534
rect 37832 3470 37884 3476
rect 36820 3392 36872 3398
rect 36820 3334 36872 3340
rect 38016 3392 38068 3398
rect 38016 3334 38068 3340
rect 36728 2984 36780 2990
rect 36728 2926 36780 2932
rect 36636 2440 36688 2446
rect 36688 2388 36768 2394
rect 36636 2382 36768 2388
rect 36452 2372 36504 2378
rect 36648 2366 36768 2382
rect 36452 2314 36504 2320
rect 2962 776 3018 785
rect 2962 711 3018 720
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36464 785 36492 2314
rect 36740 800 36768 2366
rect 36832 2145 36860 3334
rect 37924 2984 37976 2990
rect 37924 2926 37976 2932
rect 37372 2848 37424 2854
rect 37372 2790 37424 2796
rect 36818 2136 36874 2145
rect 36818 2071 36874 2080
rect 37384 800 37412 2790
rect 37936 2666 37964 2926
rect 38028 2825 38056 3334
rect 38014 2816 38070 2825
rect 38014 2751 38070 2760
rect 37936 2638 38056 2666
rect 37648 2508 37700 2514
rect 37648 2450 37700 2456
rect 36450 776 36506 785
rect 36450 711 36506 720
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 37660 105 37688 2450
rect 38028 800 38056 2638
rect 38672 800 38700 3606
rect 39316 800 39344 4150
rect 37646 96 37702 105
rect 37646 31 37702 40
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39302 0 39358 800
<< via2 >>
rect 2870 49680 2926 49736
rect 1490 45600 1546 45656
rect 1398 44240 1454 44296
rect 1398 43560 1454 43616
rect 1398 42880 1454 42936
rect 1398 42200 1454 42256
rect 1398 39516 1400 39536
rect 1400 39516 1452 39536
rect 1452 39516 1454 39536
rect 1398 39480 1454 39516
rect 1490 38820 1546 38856
rect 1490 38800 1492 38820
rect 1492 38800 1544 38820
rect 1544 38800 1546 38820
rect 1490 36760 1546 36816
rect 1490 36080 1546 36136
rect 1490 35436 1492 35456
rect 1492 35436 1544 35456
rect 1544 35436 1546 35456
rect 1490 35400 1546 35436
rect 1490 34720 1546 34776
rect 1398 33360 1454 33416
rect 1398 32680 1454 32736
rect 1490 32000 1546 32056
rect 1398 31320 1454 31376
rect 1858 41556 1860 41576
rect 1860 41556 1912 41576
rect 1912 41556 1914 41576
rect 1858 41520 1914 41556
rect 1858 40160 1914 40216
rect 2226 40840 2282 40896
rect 1490 29996 1492 30016
rect 1492 29996 1544 30016
rect 1544 29996 1546 30016
rect 1490 29960 1546 29996
rect 1490 29280 1546 29336
rect 1398 28600 1454 28656
rect 1398 27920 1454 27976
rect 1398 27240 1454 27296
rect 1490 26560 1546 26616
rect 1490 25880 1546 25936
rect 1398 24520 1454 24576
rect 1490 23160 1546 23216
rect 1398 22480 1454 22536
rect 1398 21800 1454 21856
rect 1398 20476 1400 20496
rect 1400 20476 1452 20496
rect 1452 20476 1454 20496
rect 1398 20440 1454 20476
rect 1490 19116 1492 19136
rect 1492 19116 1544 19136
rect 1544 19116 1546 19136
rect 1490 19080 1546 19116
rect 1490 18400 1546 18456
rect 1490 17720 1546 17776
rect 1398 17040 1454 17096
rect 1398 15700 1454 15736
rect 1398 15680 1400 15700
rect 1400 15680 1452 15700
rect 1452 15680 1454 15700
rect 1490 14320 1546 14376
rect 1398 12960 1454 13016
rect 1490 12280 1546 12336
rect 1490 11600 1546 11656
rect 2226 38120 2282 38176
rect 2226 37440 2282 37496
rect 2226 34040 2282 34096
rect 1858 25236 1860 25256
rect 1860 25236 1912 25256
rect 1912 25236 1914 25256
rect 1858 25200 1914 25236
rect 2042 24132 2098 24168
rect 2042 24112 2044 24132
rect 2044 24112 2096 24132
rect 2096 24112 2098 24132
rect 1858 23840 1914 23896
rect 2042 21140 2098 21176
rect 2042 21120 2044 21140
rect 2044 21120 2096 21140
rect 2096 21120 2098 21140
rect 1398 10920 1454 10976
rect 1398 10240 1454 10296
rect 1398 9560 1454 9616
rect 1490 8880 1546 8936
rect 1398 6876 1400 6896
rect 1400 6876 1452 6896
rect 1452 6876 1454 6896
rect 1398 6840 1454 6876
rect 2226 19796 2228 19816
rect 2228 19796 2280 19816
rect 2280 19796 2282 19816
rect 2226 19760 2282 19796
rect 1490 6180 1546 6216
rect 1490 6160 1492 6180
rect 1492 6160 1544 6180
rect 1544 6160 1546 6180
rect 1490 5516 1492 5536
rect 1492 5516 1544 5536
rect 1544 5516 1546 5536
rect 1490 5480 1546 5516
rect 1398 4800 1454 4856
rect 1490 4120 1546 4176
rect 2042 16360 2098 16416
rect 2042 13640 2098 13696
rect 2226 8200 2282 8256
rect 2042 7540 2098 7576
rect 2042 7520 2044 7540
rect 2044 7520 2096 7540
rect 2096 7520 2098 7540
rect 2778 47640 2834 47696
rect 2870 46960 2926 47016
rect 2778 44920 2834 44976
rect 3054 49000 3110 49056
rect 3146 48320 3202 48376
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 2226 3440 2282 3496
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 3330 2760 3386 2816
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 2870 2080 2926 2136
rect 2778 1400 2834 1456
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 32954 24112 33010 24168
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 35438 49000 35494 49056
rect 35806 48320 35862 48376
rect 35714 47640 35770 47696
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 35898 46280 35954 46336
rect 37186 45600 37242 45656
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 38106 46960 38162 47016
rect 37278 43560 37334 43616
rect 38014 44920 38070 44976
rect 38014 44260 38070 44296
rect 38014 44240 38016 44260
rect 38016 44240 38068 44260
rect 38068 44240 38070 44260
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 37186 16360 37242 16416
rect 35898 1400 35954 1456
rect 37278 11636 37280 11656
rect 37280 11636 37332 11656
rect 37332 11636 37334 11656
rect 37278 11600 37334 11636
rect 38014 42880 38070 42936
rect 38106 42200 38162 42256
rect 38106 41556 38108 41576
rect 38108 41556 38160 41576
rect 38160 41556 38162 41576
rect 38106 41520 38162 41556
rect 38106 40840 38162 40896
rect 38106 40160 38162 40216
rect 38014 39480 38070 39536
rect 38014 38820 38070 38856
rect 38014 38800 38016 38820
rect 38016 38800 38068 38820
rect 38068 38800 38070 38820
rect 38106 38120 38162 38176
rect 38014 37440 38070 37496
rect 38106 36796 38108 36816
rect 38108 36796 38160 36816
rect 38160 36796 38162 36816
rect 38106 36760 38162 36796
rect 38014 36080 38070 36136
rect 38106 35400 38162 35456
rect 38106 34040 38162 34096
rect 38106 33360 38162 33416
rect 38106 32680 38162 32736
rect 38106 32000 38162 32056
rect 38014 31320 38070 31376
rect 38014 29996 38016 30016
rect 38016 29996 38068 30016
rect 38068 29996 38070 30016
rect 38014 29960 38070 29996
rect 38106 29280 38162 29336
rect 38106 28600 38162 28656
rect 38014 27940 38070 27976
rect 38014 27920 38016 27940
rect 38016 27920 38068 27940
rect 38068 27920 38070 27940
rect 38014 27276 38016 27296
rect 38016 27276 38068 27296
rect 38068 27276 38070 27296
rect 38014 27240 38070 27276
rect 38106 26560 38162 26616
rect 38014 25880 38070 25936
rect 38106 25236 38108 25256
rect 38108 25236 38160 25256
rect 38160 25236 38162 25256
rect 38106 25200 38162 25236
rect 38106 24520 38162 24576
rect 38014 23840 38070 23896
rect 38014 23160 38070 23216
rect 38106 22516 38108 22536
rect 38108 22516 38160 22536
rect 38160 22516 38162 22536
rect 38106 22480 38162 22516
rect 38106 21800 38162 21856
rect 38014 21120 38070 21176
rect 38106 20440 38162 20496
rect 38014 19760 38070 19816
rect 38014 18400 38070 18456
rect 38106 17720 38162 17776
rect 38106 17040 38162 17096
rect 38014 15680 38070 15736
rect 38106 15000 38162 15056
rect 38106 14356 38108 14376
rect 38108 14356 38160 14376
rect 38160 14356 38162 14376
rect 38106 14320 38162 14356
rect 38014 13676 38016 13696
rect 38016 13676 38068 13696
rect 38068 13676 38070 13696
rect 38014 13640 38070 13676
rect 38014 12960 38070 13016
rect 38106 12316 38108 12336
rect 38108 12316 38160 12336
rect 38160 12316 38162 12336
rect 38106 12280 38162 12316
rect 38106 10920 38162 10976
rect 38106 10240 38162 10296
rect 38106 9560 38162 9616
rect 38106 8916 38108 8936
rect 38108 8916 38160 8936
rect 38160 8916 38162 8936
rect 38106 8880 38162 8916
rect 38014 8200 38070 8256
rect 38014 7520 38070 7576
rect 38014 6840 38070 6896
rect 38014 6180 38070 6216
rect 38014 6160 38016 6180
rect 38016 6160 38068 6180
rect 38068 6160 38070 6180
rect 38014 5516 38016 5536
rect 38016 5516 38068 5536
rect 38068 5516 38070 5536
rect 38014 5480 38070 5516
rect 38014 4800 38070 4856
rect 38014 4120 38070 4176
rect 2962 720 3018 776
rect 36818 2080 36874 2136
rect 38014 2760 38070 2816
rect 36450 720 36506 776
rect 37646 40 37702 96
<< metal3 >>
rect 0 49738 800 49768
rect 2865 49738 2931 49741
rect 0 49736 2931 49738
rect 0 49680 2870 49736
rect 2926 49680 2931 49736
rect 0 49678 2931 49680
rect 0 49648 800 49678
rect 2865 49675 2931 49678
rect 0 49058 800 49088
rect 3049 49058 3115 49061
rect 0 49056 3115 49058
rect 0 49000 3054 49056
rect 3110 49000 3115 49056
rect 0 48998 3115 49000
rect 0 48968 800 48998
rect 3049 48995 3115 48998
rect 35433 49058 35499 49061
rect 39200 49058 40000 49088
rect 35433 49056 40000 49058
rect 35433 49000 35438 49056
rect 35494 49000 40000 49056
rect 35433 48998 40000 49000
rect 35433 48995 35499 48998
rect 39200 48968 40000 48998
rect 0 48378 800 48408
rect 3141 48378 3207 48381
rect 0 48376 3207 48378
rect 0 48320 3146 48376
rect 3202 48320 3207 48376
rect 0 48318 3207 48320
rect 0 48288 800 48318
rect 3141 48315 3207 48318
rect 35801 48378 35867 48381
rect 39200 48378 40000 48408
rect 35801 48376 40000 48378
rect 35801 48320 35806 48376
rect 35862 48320 40000 48376
rect 35801 48318 40000 48320
rect 35801 48315 35867 48318
rect 39200 48288 40000 48318
rect 0 47698 800 47728
rect 2773 47698 2839 47701
rect 0 47696 2839 47698
rect 0 47640 2778 47696
rect 2834 47640 2839 47696
rect 0 47638 2839 47640
rect 0 47608 800 47638
rect 2773 47635 2839 47638
rect 35709 47698 35775 47701
rect 39200 47698 40000 47728
rect 35709 47696 40000 47698
rect 35709 47640 35714 47696
rect 35770 47640 40000 47696
rect 35709 47638 40000 47640
rect 35709 47635 35775 47638
rect 39200 47608 40000 47638
rect 4210 47360 4526 47361
rect 4210 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4526 47360
rect 4210 47295 4526 47296
rect 34930 47360 35246 47361
rect 34930 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35246 47360
rect 34930 47295 35246 47296
rect 0 47018 800 47048
rect 2865 47018 2931 47021
rect 0 47016 2931 47018
rect 0 46960 2870 47016
rect 2926 46960 2931 47016
rect 0 46958 2931 46960
rect 0 46928 800 46958
rect 2865 46955 2931 46958
rect 38101 47018 38167 47021
rect 39200 47018 40000 47048
rect 38101 47016 40000 47018
rect 38101 46960 38106 47016
rect 38162 46960 40000 47016
rect 38101 46958 40000 46960
rect 38101 46955 38167 46958
rect 39200 46928 40000 46958
rect 19570 46816 19886 46817
rect 19570 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19886 46816
rect 19570 46751 19886 46752
rect 35893 46338 35959 46341
rect 39200 46338 40000 46368
rect 35893 46336 40000 46338
rect 35893 46280 35898 46336
rect 35954 46280 40000 46336
rect 35893 46278 40000 46280
rect 35893 46275 35959 46278
rect 4210 46272 4526 46273
rect 4210 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4526 46272
rect 4210 46207 4526 46208
rect 34930 46272 35246 46273
rect 34930 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35246 46272
rect 39200 46248 40000 46278
rect 34930 46207 35246 46208
rect 19570 45728 19886 45729
rect 0 45658 800 45688
rect 19570 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19886 45728
rect 19570 45663 19886 45664
rect 1485 45658 1551 45661
rect 0 45656 1551 45658
rect 0 45600 1490 45656
rect 1546 45600 1551 45656
rect 0 45598 1551 45600
rect 0 45568 800 45598
rect 1485 45595 1551 45598
rect 37181 45658 37247 45661
rect 39200 45658 40000 45688
rect 37181 45656 40000 45658
rect 37181 45600 37186 45656
rect 37242 45600 40000 45656
rect 37181 45598 40000 45600
rect 37181 45595 37247 45598
rect 39200 45568 40000 45598
rect 4210 45184 4526 45185
rect 4210 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4526 45184
rect 4210 45119 4526 45120
rect 34930 45184 35246 45185
rect 34930 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35246 45184
rect 34930 45119 35246 45120
rect 0 44978 800 45008
rect 2773 44978 2839 44981
rect 0 44976 2839 44978
rect 0 44920 2778 44976
rect 2834 44920 2839 44976
rect 0 44918 2839 44920
rect 0 44888 800 44918
rect 2773 44915 2839 44918
rect 38009 44978 38075 44981
rect 39200 44978 40000 45008
rect 38009 44976 40000 44978
rect 38009 44920 38014 44976
rect 38070 44920 40000 44976
rect 38009 44918 40000 44920
rect 38009 44915 38075 44918
rect 39200 44888 40000 44918
rect 19570 44640 19886 44641
rect 19570 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19886 44640
rect 19570 44575 19886 44576
rect 0 44298 800 44328
rect 1393 44298 1459 44301
rect 0 44296 1459 44298
rect 0 44240 1398 44296
rect 1454 44240 1459 44296
rect 0 44238 1459 44240
rect 0 44208 800 44238
rect 1393 44235 1459 44238
rect 38009 44298 38075 44301
rect 39200 44298 40000 44328
rect 38009 44296 40000 44298
rect 38009 44240 38014 44296
rect 38070 44240 40000 44296
rect 38009 44238 40000 44240
rect 38009 44235 38075 44238
rect 39200 44208 40000 44238
rect 4210 44096 4526 44097
rect 4210 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4526 44096
rect 4210 44031 4526 44032
rect 34930 44096 35246 44097
rect 34930 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35246 44096
rect 34930 44031 35246 44032
rect 0 43618 800 43648
rect 1393 43618 1459 43621
rect 0 43616 1459 43618
rect 0 43560 1398 43616
rect 1454 43560 1459 43616
rect 0 43558 1459 43560
rect 0 43528 800 43558
rect 1393 43555 1459 43558
rect 37273 43618 37339 43621
rect 39200 43618 40000 43648
rect 37273 43616 40000 43618
rect 37273 43560 37278 43616
rect 37334 43560 40000 43616
rect 37273 43558 40000 43560
rect 37273 43555 37339 43558
rect 19570 43552 19886 43553
rect 19570 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19886 43552
rect 39200 43528 40000 43558
rect 19570 43487 19886 43488
rect 4210 43008 4526 43009
rect 0 42938 800 42968
rect 4210 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4526 43008
rect 4210 42943 4526 42944
rect 34930 43008 35246 43009
rect 34930 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35246 43008
rect 34930 42943 35246 42944
rect 1393 42938 1459 42941
rect 0 42936 1459 42938
rect 0 42880 1398 42936
rect 1454 42880 1459 42936
rect 0 42878 1459 42880
rect 0 42848 800 42878
rect 1393 42875 1459 42878
rect 38009 42938 38075 42941
rect 39200 42938 40000 42968
rect 38009 42936 40000 42938
rect 38009 42880 38014 42936
rect 38070 42880 40000 42936
rect 38009 42878 40000 42880
rect 38009 42875 38075 42878
rect 39200 42848 40000 42878
rect 19570 42464 19886 42465
rect 19570 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19886 42464
rect 19570 42399 19886 42400
rect 0 42258 800 42288
rect 1393 42258 1459 42261
rect 0 42256 1459 42258
rect 0 42200 1398 42256
rect 1454 42200 1459 42256
rect 0 42198 1459 42200
rect 0 42168 800 42198
rect 1393 42195 1459 42198
rect 38101 42258 38167 42261
rect 39200 42258 40000 42288
rect 38101 42256 40000 42258
rect 38101 42200 38106 42256
rect 38162 42200 40000 42256
rect 38101 42198 40000 42200
rect 38101 42195 38167 42198
rect 39200 42168 40000 42198
rect 4210 41920 4526 41921
rect 4210 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4526 41920
rect 4210 41855 4526 41856
rect 34930 41920 35246 41921
rect 34930 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35246 41920
rect 34930 41855 35246 41856
rect 0 41578 800 41608
rect 1853 41578 1919 41581
rect 0 41576 1919 41578
rect 0 41520 1858 41576
rect 1914 41520 1919 41576
rect 0 41518 1919 41520
rect 0 41488 800 41518
rect 1853 41515 1919 41518
rect 38101 41578 38167 41581
rect 39200 41578 40000 41608
rect 38101 41576 40000 41578
rect 38101 41520 38106 41576
rect 38162 41520 40000 41576
rect 38101 41518 40000 41520
rect 38101 41515 38167 41518
rect 39200 41488 40000 41518
rect 19570 41376 19886 41377
rect 19570 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19886 41376
rect 19570 41311 19886 41312
rect 0 40898 800 40928
rect 2221 40898 2287 40901
rect 0 40896 2287 40898
rect 0 40840 2226 40896
rect 2282 40840 2287 40896
rect 0 40838 2287 40840
rect 0 40808 800 40838
rect 2221 40835 2287 40838
rect 38101 40898 38167 40901
rect 39200 40898 40000 40928
rect 38101 40896 40000 40898
rect 38101 40840 38106 40896
rect 38162 40840 40000 40896
rect 38101 40838 40000 40840
rect 38101 40835 38167 40838
rect 4210 40832 4526 40833
rect 4210 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4526 40832
rect 4210 40767 4526 40768
rect 34930 40832 35246 40833
rect 34930 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35246 40832
rect 39200 40808 40000 40838
rect 34930 40767 35246 40768
rect 19570 40288 19886 40289
rect 0 40218 800 40248
rect 19570 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19886 40288
rect 19570 40223 19886 40224
rect 1853 40218 1919 40221
rect 0 40216 1919 40218
rect 0 40160 1858 40216
rect 1914 40160 1919 40216
rect 0 40158 1919 40160
rect 0 40128 800 40158
rect 1853 40155 1919 40158
rect 38101 40218 38167 40221
rect 39200 40218 40000 40248
rect 38101 40216 40000 40218
rect 38101 40160 38106 40216
rect 38162 40160 40000 40216
rect 38101 40158 40000 40160
rect 38101 40155 38167 40158
rect 39200 40128 40000 40158
rect 4210 39744 4526 39745
rect 4210 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4526 39744
rect 4210 39679 4526 39680
rect 34930 39744 35246 39745
rect 34930 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35246 39744
rect 34930 39679 35246 39680
rect 0 39538 800 39568
rect 1393 39538 1459 39541
rect 0 39536 1459 39538
rect 0 39480 1398 39536
rect 1454 39480 1459 39536
rect 0 39478 1459 39480
rect 0 39448 800 39478
rect 1393 39475 1459 39478
rect 38009 39538 38075 39541
rect 39200 39538 40000 39568
rect 38009 39536 40000 39538
rect 38009 39480 38014 39536
rect 38070 39480 40000 39536
rect 38009 39478 40000 39480
rect 38009 39475 38075 39478
rect 39200 39448 40000 39478
rect 19570 39200 19886 39201
rect 19570 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19886 39200
rect 19570 39135 19886 39136
rect 0 38858 800 38888
rect 1485 38858 1551 38861
rect 0 38856 1551 38858
rect 0 38800 1490 38856
rect 1546 38800 1551 38856
rect 0 38798 1551 38800
rect 0 38768 800 38798
rect 1485 38795 1551 38798
rect 38009 38858 38075 38861
rect 39200 38858 40000 38888
rect 38009 38856 40000 38858
rect 38009 38800 38014 38856
rect 38070 38800 40000 38856
rect 38009 38798 40000 38800
rect 38009 38795 38075 38798
rect 39200 38768 40000 38798
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 0 38178 800 38208
rect 2221 38178 2287 38181
rect 0 38176 2287 38178
rect 0 38120 2226 38176
rect 2282 38120 2287 38176
rect 0 38118 2287 38120
rect 0 38088 800 38118
rect 2221 38115 2287 38118
rect 38101 38178 38167 38181
rect 39200 38178 40000 38208
rect 38101 38176 40000 38178
rect 38101 38120 38106 38176
rect 38162 38120 40000 38176
rect 38101 38118 40000 38120
rect 38101 38115 38167 38118
rect 19570 38112 19886 38113
rect 19570 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19886 38112
rect 39200 38088 40000 38118
rect 19570 38047 19886 38048
rect 4210 37568 4526 37569
rect 0 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 2221 37498 2287 37501
rect 0 37496 2287 37498
rect 0 37440 2226 37496
rect 2282 37440 2287 37496
rect 0 37438 2287 37440
rect 0 37408 800 37438
rect 2221 37435 2287 37438
rect 38009 37498 38075 37501
rect 39200 37498 40000 37528
rect 38009 37496 40000 37498
rect 38009 37440 38014 37496
rect 38070 37440 40000 37496
rect 38009 37438 40000 37440
rect 38009 37435 38075 37438
rect 39200 37408 40000 37438
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 0 36818 800 36848
rect 1485 36818 1551 36821
rect 0 36816 1551 36818
rect 0 36760 1490 36816
rect 1546 36760 1551 36816
rect 0 36758 1551 36760
rect 0 36728 800 36758
rect 1485 36755 1551 36758
rect 38101 36818 38167 36821
rect 39200 36818 40000 36848
rect 38101 36816 40000 36818
rect 38101 36760 38106 36816
rect 38162 36760 40000 36816
rect 38101 36758 40000 36760
rect 38101 36755 38167 36758
rect 39200 36728 40000 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 0 36138 800 36168
rect 1485 36138 1551 36141
rect 0 36136 1551 36138
rect 0 36080 1490 36136
rect 1546 36080 1551 36136
rect 0 36078 1551 36080
rect 0 36048 800 36078
rect 1485 36075 1551 36078
rect 38009 36138 38075 36141
rect 39200 36138 40000 36168
rect 38009 36136 40000 36138
rect 38009 36080 38014 36136
rect 38070 36080 40000 36136
rect 38009 36078 40000 36080
rect 38009 36075 38075 36078
rect 39200 36048 40000 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 0 35458 800 35488
rect 1485 35458 1551 35461
rect 0 35456 1551 35458
rect 0 35400 1490 35456
rect 1546 35400 1551 35456
rect 0 35398 1551 35400
rect 0 35368 800 35398
rect 1485 35395 1551 35398
rect 38101 35458 38167 35461
rect 39200 35458 40000 35488
rect 38101 35456 40000 35458
rect 38101 35400 38106 35456
rect 38162 35400 40000 35456
rect 38101 35398 40000 35400
rect 38101 35395 38167 35398
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 39200 35368 40000 35398
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 0 34778 800 34808
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 1485 34778 1551 34781
rect 0 34776 1551 34778
rect 0 34720 1490 34776
rect 1546 34720 1551 34776
rect 0 34718 1551 34720
rect 0 34688 800 34718
rect 1485 34715 1551 34718
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 0 34098 800 34128
rect 2221 34098 2287 34101
rect 0 34096 2287 34098
rect 0 34040 2226 34096
rect 2282 34040 2287 34096
rect 0 34038 2287 34040
rect 0 34008 800 34038
rect 2221 34035 2287 34038
rect 38101 34098 38167 34101
rect 39200 34098 40000 34128
rect 38101 34096 40000 34098
rect 38101 34040 38106 34096
rect 38162 34040 40000 34096
rect 38101 34038 40000 34040
rect 38101 34035 38167 34038
rect 39200 34008 40000 34038
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 0 33418 800 33448
rect 1393 33418 1459 33421
rect 0 33416 1459 33418
rect 0 33360 1398 33416
rect 1454 33360 1459 33416
rect 0 33358 1459 33360
rect 0 33328 800 33358
rect 1393 33355 1459 33358
rect 38101 33418 38167 33421
rect 39200 33418 40000 33448
rect 38101 33416 40000 33418
rect 38101 33360 38106 33416
rect 38162 33360 40000 33416
rect 38101 33358 40000 33360
rect 38101 33355 38167 33358
rect 39200 33328 40000 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 0 32738 800 32768
rect 1393 32738 1459 32741
rect 0 32736 1459 32738
rect 0 32680 1398 32736
rect 1454 32680 1459 32736
rect 0 32678 1459 32680
rect 0 32648 800 32678
rect 1393 32675 1459 32678
rect 38101 32738 38167 32741
rect 39200 32738 40000 32768
rect 38101 32736 40000 32738
rect 38101 32680 38106 32736
rect 38162 32680 40000 32736
rect 38101 32678 40000 32680
rect 38101 32675 38167 32678
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 39200 32648 40000 32678
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 0 32058 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 1485 32058 1551 32061
rect 0 32056 1551 32058
rect 0 32000 1490 32056
rect 1546 32000 1551 32056
rect 0 31998 1551 32000
rect 0 31968 800 31998
rect 1485 31995 1551 31998
rect 38101 32058 38167 32061
rect 39200 32058 40000 32088
rect 38101 32056 40000 32058
rect 38101 32000 38106 32056
rect 38162 32000 40000 32056
rect 38101 31998 40000 32000
rect 38101 31995 38167 31998
rect 39200 31968 40000 31998
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 0 31378 800 31408
rect 1393 31378 1459 31381
rect 0 31376 1459 31378
rect 0 31320 1398 31376
rect 1454 31320 1459 31376
rect 0 31318 1459 31320
rect 0 31288 800 31318
rect 1393 31315 1459 31318
rect 38009 31378 38075 31381
rect 39200 31378 40000 31408
rect 38009 31376 40000 31378
rect 38009 31320 38014 31376
rect 38070 31320 40000 31376
rect 38009 31318 40000 31320
rect 38009 31315 38075 31318
rect 39200 31288 40000 31318
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 39200 30608 40000 30728
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 0 30018 800 30048
rect 1485 30018 1551 30021
rect 0 30016 1551 30018
rect 0 29960 1490 30016
rect 1546 29960 1551 30016
rect 0 29958 1551 29960
rect 0 29928 800 29958
rect 1485 29955 1551 29958
rect 38009 30018 38075 30021
rect 39200 30018 40000 30048
rect 38009 30016 40000 30018
rect 38009 29960 38014 30016
rect 38070 29960 40000 30016
rect 38009 29958 40000 29960
rect 38009 29955 38075 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 39200 29928 40000 29958
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 0 29338 800 29368
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 1485 29338 1551 29341
rect 0 29336 1551 29338
rect 0 29280 1490 29336
rect 1546 29280 1551 29336
rect 0 29278 1551 29280
rect 0 29248 800 29278
rect 1485 29275 1551 29278
rect 38101 29338 38167 29341
rect 39200 29338 40000 29368
rect 38101 29336 40000 29338
rect 38101 29280 38106 29336
rect 38162 29280 40000 29336
rect 38101 29278 40000 29280
rect 38101 29275 38167 29278
rect 39200 29248 40000 29278
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 0 28658 800 28688
rect 1393 28658 1459 28661
rect 0 28656 1459 28658
rect 0 28600 1398 28656
rect 1454 28600 1459 28656
rect 0 28598 1459 28600
rect 0 28568 800 28598
rect 1393 28595 1459 28598
rect 38101 28658 38167 28661
rect 39200 28658 40000 28688
rect 38101 28656 40000 28658
rect 38101 28600 38106 28656
rect 38162 28600 40000 28656
rect 38101 28598 40000 28600
rect 38101 28595 38167 28598
rect 39200 28568 40000 28598
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 0 27978 800 28008
rect 1393 27978 1459 27981
rect 0 27976 1459 27978
rect 0 27920 1398 27976
rect 1454 27920 1459 27976
rect 0 27918 1459 27920
rect 0 27888 800 27918
rect 1393 27915 1459 27918
rect 38009 27978 38075 27981
rect 39200 27978 40000 28008
rect 38009 27976 40000 27978
rect 38009 27920 38014 27976
rect 38070 27920 40000 27976
rect 38009 27918 40000 27920
rect 38009 27915 38075 27918
rect 39200 27888 40000 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 0 27298 800 27328
rect 1393 27298 1459 27301
rect 0 27296 1459 27298
rect 0 27240 1398 27296
rect 1454 27240 1459 27296
rect 0 27238 1459 27240
rect 0 27208 800 27238
rect 1393 27235 1459 27238
rect 38009 27298 38075 27301
rect 39200 27298 40000 27328
rect 38009 27296 40000 27298
rect 38009 27240 38014 27296
rect 38070 27240 40000 27296
rect 38009 27238 40000 27240
rect 38009 27235 38075 27238
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 39200 27208 40000 27238
rect 19570 27167 19886 27168
rect 4210 26688 4526 26689
rect 0 26618 800 26648
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 1485 26618 1551 26621
rect 0 26616 1551 26618
rect 0 26560 1490 26616
rect 1546 26560 1551 26616
rect 0 26558 1551 26560
rect 0 26528 800 26558
rect 1485 26555 1551 26558
rect 38101 26618 38167 26621
rect 39200 26618 40000 26648
rect 38101 26616 40000 26618
rect 38101 26560 38106 26616
rect 38162 26560 40000 26616
rect 38101 26558 40000 26560
rect 38101 26555 38167 26558
rect 39200 26528 40000 26558
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 0 25938 800 25968
rect 1485 25938 1551 25941
rect 0 25936 1551 25938
rect 0 25880 1490 25936
rect 1546 25880 1551 25936
rect 0 25878 1551 25880
rect 0 25848 800 25878
rect 1485 25875 1551 25878
rect 38009 25938 38075 25941
rect 39200 25938 40000 25968
rect 38009 25936 40000 25938
rect 38009 25880 38014 25936
rect 38070 25880 40000 25936
rect 38009 25878 40000 25880
rect 38009 25875 38075 25878
rect 39200 25848 40000 25878
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 0 25258 800 25288
rect 1853 25258 1919 25261
rect 0 25256 1919 25258
rect 0 25200 1858 25256
rect 1914 25200 1919 25256
rect 0 25198 1919 25200
rect 0 25168 800 25198
rect 1853 25195 1919 25198
rect 38101 25258 38167 25261
rect 39200 25258 40000 25288
rect 38101 25256 40000 25258
rect 38101 25200 38106 25256
rect 38162 25200 40000 25256
rect 38101 25198 40000 25200
rect 38101 25195 38167 25198
rect 39200 25168 40000 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 0 24578 800 24608
rect 1393 24578 1459 24581
rect 0 24576 1459 24578
rect 0 24520 1398 24576
rect 1454 24520 1459 24576
rect 0 24518 1459 24520
rect 0 24488 800 24518
rect 1393 24515 1459 24518
rect 38101 24578 38167 24581
rect 39200 24578 40000 24608
rect 38101 24576 40000 24578
rect 38101 24520 38106 24576
rect 38162 24520 40000 24576
rect 38101 24518 40000 24520
rect 38101 24515 38167 24518
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 39200 24488 40000 24518
rect 34930 24447 35246 24448
rect 2037 24170 2103 24173
rect 32949 24170 33015 24173
rect 2037 24168 33015 24170
rect 2037 24112 2042 24168
rect 2098 24112 32954 24168
rect 33010 24112 33015 24168
rect 2037 24110 33015 24112
rect 2037 24107 2103 24110
rect 32949 24107 33015 24110
rect 19570 23968 19886 23969
rect 0 23898 800 23928
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 1853 23898 1919 23901
rect 0 23896 1919 23898
rect 0 23840 1858 23896
rect 1914 23840 1919 23896
rect 0 23838 1919 23840
rect 0 23808 800 23838
rect 1853 23835 1919 23838
rect 38009 23898 38075 23901
rect 39200 23898 40000 23928
rect 38009 23896 40000 23898
rect 38009 23840 38014 23896
rect 38070 23840 40000 23896
rect 38009 23838 40000 23840
rect 38009 23835 38075 23838
rect 39200 23808 40000 23838
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 0 23218 800 23248
rect 1485 23218 1551 23221
rect 0 23216 1551 23218
rect 0 23160 1490 23216
rect 1546 23160 1551 23216
rect 0 23158 1551 23160
rect 0 23128 800 23158
rect 1485 23155 1551 23158
rect 38009 23218 38075 23221
rect 39200 23218 40000 23248
rect 38009 23216 40000 23218
rect 38009 23160 38014 23216
rect 38070 23160 40000 23216
rect 38009 23158 40000 23160
rect 38009 23155 38075 23158
rect 39200 23128 40000 23158
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 0 22538 800 22568
rect 1393 22538 1459 22541
rect 0 22536 1459 22538
rect 0 22480 1398 22536
rect 1454 22480 1459 22536
rect 0 22478 1459 22480
rect 0 22448 800 22478
rect 1393 22475 1459 22478
rect 38101 22538 38167 22541
rect 39200 22538 40000 22568
rect 38101 22536 40000 22538
rect 38101 22480 38106 22536
rect 38162 22480 40000 22536
rect 38101 22478 40000 22480
rect 38101 22475 38167 22478
rect 39200 22448 40000 22478
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 0 21858 800 21888
rect 1393 21858 1459 21861
rect 0 21856 1459 21858
rect 0 21800 1398 21856
rect 1454 21800 1459 21856
rect 0 21798 1459 21800
rect 0 21768 800 21798
rect 1393 21795 1459 21798
rect 38101 21858 38167 21861
rect 39200 21858 40000 21888
rect 38101 21856 40000 21858
rect 38101 21800 38106 21856
rect 38162 21800 40000 21856
rect 38101 21798 40000 21800
rect 38101 21795 38167 21798
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 39200 21768 40000 21798
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 0 21178 800 21208
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 2037 21178 2103 21181
rect 0 21176 2103 21178
rect 0 21120 2042 21176
rect 2098 21120 2103 21176
rect 0 21118 2103 21120
rect 0 21088 800 21118
rect 2037 21115 2103 21118
rect 38009 21178 38075 21181
rect 39200 21178 40000 21208
rect 38009 21176 40000 21178
rect 38009 21120 38014 21176
rect 38070 21120 40000 21176
rect 38009 21118 40000 21120
rect 38009 21115 38075 21118
rect 39200 21088 40000 21118
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 0 20498 800 20528
rect 1393 20498 1459 20501
rect 0 20496 1459 20498
rect 0 20440 1398 20496
rect 1454 20440 1459 20496
rect 0 20438 1459 20440
rect 0 20408 800 20438
rect 1393 20435 1459 20438
rect 38101 20498 38167 20501
rect 39200 20498 40000 20528
rect 38101 20496 40000 20498
rect 38101 20440 38106 20496
rect 38162 20440 40000 20496
rect 38101 20438 40000 20440
rect 38101 20435 38167 20438
rect 39200 20408 40000 20438
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 0 19818 800 19848
rect 2221 19818 2287 19821
rect 0 19816 2287 19818
rect 0 19760 2226 19816
rect 2282 19760 2287 19816
rect 0 19758 2287 19760
rect 0 19728 800 19758
rect 2221 19755 2287 19758
rect 38009 19818 38075 19821
rect 39200 19818 40000 19848
rect 38009 19816 40000 19818
rect 38009 19760 38014 19816
rect 38070 19760 40000 19816
rect 38009 19758 40000 19760
rect 38009 19755 38075 19758
rect 39200 19728 40000 19758
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 0 19138 800 19168
rect 1485 19138 1551 19141
rect 0 19136 1551 19138
rect 0 19080 1490 19136
rect 1546 19080 1551 19136
rect 0 19078 1551 19080
rect 0 19048 800 19078
rect 1485 19075 1551 19078
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 0 18458 800 18488
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 1485 18458 1551 18461
rect 0 18456 1551 18458
rect 0 18400 1490 18456
rect 1546 18400 1551 18456
rect 0 18398 1551 18400
rect 0 18368 800 18398
rect 1485 18395 1551 18398
rect 38009 18458 38075 18461
rect 39200 18458 40000 18488
rect 38009 18456 40000 18458
rect 38009 18400 38014 18456
rect 38070 18400 40000 18456
rect 38009 18398 40000 18400
rect 38009 18395 38075 18398
rect 39200 18368 40000 18398
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 0 17778 800 17808
rect 1485 17778 1551 17781
rect 0 17776 1551 17778
rect 0 17720 1490 17776
rect 1546 17720 1551 17776
rect 0 17718 1551 17720
rect 0 17688 800 17718
rect 1485 17715 1551 17718
rect 38101 17778 38167 17781
rect 39200 17778 40000 17808
rect 38101 17776 40000 17778
rect 38101 17720 38106 17776
rect 38162 17720 40000 17776
rect 38101 17718 40000 17720
rect 38101 17715 38167 17718
rect 39200 17688 40000 17718
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 0 17098 800 17128
rect 1393 17098 1459 17101
rect 0 17096 1459 17098
rect 0 17040 1398 17096
rect 1454 17040 1459 17096
rect 0 17038 1459 17040
rect 0 17008 800 17038
rect 1393 17035 1459 17038
rect 38101 17098 38167 17101
rect 39200 17098 40000 17128
rect 38101 17096 40000 17098
rect 38101 17040 38106 17096
rect 38162 17040 40000 17096
rect 38101 17038 40000 17040
rect 38101 17035 38167 17038
rect 39200 17008 40000 17038
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 0 16418 800 16448
rect 2037 16418 2103 16421
rect 0 16416 2103 16418
rect 0 16360 2042 16416
rect 2098 16360 2103 16416
rect 0 16358 2103 16360
rect 0 16328 800 16358
rect 2037 16355 2103 16358
rect 37181 16418 37247 16421
rect 39200 16418 40000 16448
rect 37181 16416 40000 16418
rect 37181 16360 37186 16416
rect 37242 16360 40000 16416
rect 37181 16358 40000 16360
rect 37181 16355 37247 16358
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 39200 16328 40000 16358
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 1393 15738 1459 15741
rect 0 15736 1459 15738
rect 0 15680 1398 15736
rect 1454 15680 1459 15736
rect 0 15678 1459 15680
rect 0 15648 800 15678
rect 1393 15675 1459 15678
rect 38009 15738 38075 15741
rect 39200 15738 40000 15768
rect 38009 15736 40000 15738
rect 38009 15680 38014 15736
rect 38070 15680 40000 15736
rect 38009 15678 40000 15680
rect 38009 15675 38075 15678
rect 39200 15648 40000 15678
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 38101 15058 38167 15061
rect 39200 15058 40000 15088
rect 38101 15056 40000 15058
rect 38101 15000 38106 15056
rect 38162 15000 40000 15056
rect 38101 14998 40000 15000
rect 38101 14995 38167 14998
rect 39200 14968 40000 14998
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 0 14378 800 14408
rect 1485 14378 1551 14381
rect 0 14376 1551 14378
rect 0 14320 1490 14376
rect 1546 14320 1551 14376
rect 0 14318 1551 14320
rect 0 14288 800 14318
rect 1485 14315 1551 14318
rect 38101 14378 38167 14381
rect 39200 14378 40000 14408
rect 38101 14376 40000 14378
rect 38101 14320 38106 14376
rect 38162 14320 40000 14376
rect 38101 14318 40000 14320
rect 38101 14315 38167 14318
rect 39200 14288 40000 14318
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 0 13698 800 13728
rect 2037 13698 2103 13701
rect 0 13696 2103 13698
rect 0 13640 2042 13696
rect 2098 13640 2103 13696
rect 0 13638 2103 13640
rect 0 13608 800 13638
rect 2037 13635 2103 13638
rect 38009 13698 38075 13701
rect 39200 13698 40000 13728
rect 38009 13696 40000 13698
rect 38009 13640 38014 13696
rect 38070 13640 40000 13696
rect 38009 13638 40000 13640
rect 38009 13635 38075 13638
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 39200 13608 40000 13638
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 0 13018 800 13048
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 1393 13018 1459 13021
rect 0 13016 1459 13018
rect 0 12960 1398 13016
rect 1454 12960 1459 13016
rect 0 12958 1459 12960
rect 0 12928 800 12958
rect 1393 12955 1459 12958
rect 38009 13018 38075 13021
rect 39200 13018 40000 13048
rect 38009 13016 40000 13018
rect 38009 12960 38014 13016
rect 38070 12960 40000 13016
rect 38009 12958 40000 12960
rect 38009 12955 38075 12958
rect 39200 12928 40000 12958
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 0 12338 800 12368
rect 1485 12338 1551 12341
rect 0 12336 1551 12338
rect 0 12280 1490 12336
rect 1546 12280 1551 12336
rect 0 12278 1551 12280
rect 0 12248 800 12278
rect 1485 12275 1551 12278
rect 38101 12338 38167 12341
rect 39200 12338 40000 12368
rect 38101 12336 40000 12338
rect 38101 12280 38106 12336
rect 38162 12280 40000 12336
rect 38101 12278 40000 12280
rect 38101 12275 38167 12278
rect 39200 12248 40000 12278
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 0 11658 800 11688
rect 1485 11658 1551 11661
rect 0 11656 1551 11658
rect 0 11600 1490 11656
rect 1546 11600 1551 11656
rect 0 11598 1551 11600
rect 0 11568 800 11598
rect 1485 11595 1551 11598
rect 37273 11658 37339 11661
rect 39200 11658 40000 11688
rect 37273 11656 40000 11658
rect 37273 11600 37278 11656
rect 37334 11600 40000 11656
rect 37273 11598 40000 11600
rect 37273 11595 37339 11598
rect 39200 11568 40000 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 38101 10978 38167 10981
rect 39200 10978 40000 11008
rect 38101 10976 40000 10978
rect 38101 10920 38106 10976
rect 38162 10920 40000 10976
rect 38101 10918 40000 10920
rect 38101 10915 38167 10918
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 39200 10888 40000 10918
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 0 10298 800 10328
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 1393 10298 1459 10301
rect 0 10296 1459 10298
rect 0 10240 1398 10296
rect 1454 10240 1459 10296
rect 0 10238 1459 10240
rect 0 10208 800 10238
rect 1393 10235 1459 10238
rect 38101 10298 38167 10301
rect 39200 10298 40000 10328
rect 38101 10296 40000 10298
rect 38101 10240 38106 10296
rect 38162 10240 40000 10296
rect 38101 10238 40000 10240
rect 38101 10235 38167 10238
rect 39200 10208 40000 10238
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 0 9618 800 9648
rect 1393 9618 1459 9621
rect 0 9616 1459 9618
rect 0 9560 1398 9616
rect 1454 9560 1459 9616
rect 0 9558 1459 9560
rect 0 9528 800 9558
rect 1393 9555 1459 9558
rect 38101 9618 38167 9621
rect 39200 9618 40000 9648
rect 38101 9616 40000 9618
rect 38101 9560 38106 9616
rect 38162 9560 40000 9616
rect 38101 9558 40000 9560
rect 38101 9555 38167 9558
rect 39200 9528 40000 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 0 8938 800 8968
rect 1485 8938 1551 8941
rect 0 8936 1551 8938
rect 0 8880 1490 8936
rect 1546 8880 1551 8936
rect 0 8878 1551 8880
rect 0 8848 800 8878
rect 1485 8875 1551 8878
rect 38101 8938 38167 8941
rect 39200 8938 40000 8968
rect 38101 8936 40000 8938
rect 38101 8880 38106 8936
rect 38162 8880 40000 8936
rect 38101 8878 40000 8880
rect 38101 8875 38167 8878
rect 39200 8848 40000 8878
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 0 8258 800 8288
rect 2221 8258 2287 8261
rect 0 8256 2287 8258
rect 0 8200 2226 8256
rect 2282 8200 2287 8256
rect 0 8198 2287 8200
rect 0 8168 800 8198
rect 2221 8195 2287 8198
rect 38009 8258 38075 8261
rect 39200 8258 40000 8288
rect 38009 8256 40000 8258
rect 38009 8200 38014 8256
rect 38070 8200 40000 8256
rect 38009 8198 40000 8200
rect 38009 8195 38075 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 39200 8168 40000 8198
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 0 7578 800 7608
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 2037 7578 2103 7581
rect 0 7576 2103 7578
rect 0 7520 2042 7576
rect 2098 7520 2103 7576
rect 0 7518 2103 7520
rect 0 7488 800 7518
rect 2037 7515 2103 7518
rect 38009 7578 38075 7581
rect 39200 7578 40000 7608
rect 38009 7576 40000 7578
rect 38009 7520 38014 7576
rect 38070 7520 40000 7576
rect 38009 7518 40000 7520
rect 38009 7515 38075 7518
rect 39200 7488 40000 7518
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 0 6898 800 6928
rect 1393 6898 1459 6901
rect 0 6896 1459 6898
rect 0 6840 1398 6896
rect 1454 6840 1459 6896
rect 0 6838 1459 6840
rect 0 6808 800 6838
rect 1393 6835 1459 6838
rect 38009 6898 38075 6901
rect 39200 6898 40000 6928
rect 38009 6896 40000 6898
rect 38009 6840 38014 6896
rect 38070 6840 40000 6896
rect 38009 6838 40000 6840
rect 38009 6835 38075 6838
rect 39200 6808 40000 6838
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 0 6218 800 6248
rect 1485 6218 1551 6221
rect 0 6216 1551 6218
rect 0 6160 1490 6216
rect 1546 6160 1551 6216
rect 0 6158 1551 6160
rect 0 6128 800 6158
rect 1485 6155 1551 6158
rect 38009 6218 38075 6221
rect 39200 6218 40000 6248
rect 38009 6216 40000 6218
rect 38009 6160 38014 6216
rect 38070 6160 40000 6216
rect 38009 6158 40000 6160
rect 38009 6155 38075 6158
rect 39200 6128 40000 6158
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 0 5538 800 5568
rect 1485 5538 1551 5541
rect 0 5536 1551 5538
rect 0 5480 1490 5536
rect 1546 5480 1551 5536
rect 0 5478 1551 5480
rect 0 5448 800 5478
rect 1485 5475 1551 5478
rect 38009 5538 38075 5541
rect 39200 5538 40000 5568
rect 38009 5536 40000 5538
rect 38009 5480 38014 5536
rect 38070 5480 40000 5536
rect 38009 5478 40000 5480
rect 38009 5475 38075 5478
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 39200 5448 40000 5478
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 0 4858 800 4888
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 1393 4858 1459 4861
rect 0 4856 1459 4858
rect 0 4800 1398 4856
rect 1454 4800 1459 4856
rect 0 4798 1459 4800
rect 0 4768 800 4798
rect 1393 4795 1459 4798
rect 38009 4858 38075 4861
rect 39200 4858 40000 4888
rect 38009 4856 40000 4858
rect 38009 4800 38014 4856
rect 38070 4800 40000 4856
rect 38009 4798 40000 4800
rect 38009 4795 38075 4798
rect 39200 4768 40000 4798
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 0 4178 800 4208
rect 1485 4178 1551 4181
rect 0 4176 1551 4178
rect 0 4120 1490 4176
rect 1546 4120 1551 4176
rect 0 4118 1551 4120
rect 0 4088 800 4118
rect 1485 4115 1551 4118
rect 38009 4178 38075 4181
rect 39200 4178 40000 4208
rect 38009 4176 40000 4178
rect 38009 4120 38014 4176
rect 38070 4120 40000 4176
rect 38009 4118 40000 4120
rect 38009 4115 38075 4118
rect 39200 4088 40000 4118
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 0 3498 800 3528
rect 2221 3498 2287 3501
rect 0 3496 2287 3498
rect 0 3440 2226 3496
rect 2282 3440 2287 3496
rect 0 3438 2287 3440
rect 0 3408 800 3438
rect 2221 3435 2287 3438
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 0 2818 800 2848
rect 3325 2818 3391 2821
rect 0 2816 3391 2818
rect 0 2760 3330 2816
rect 3386 2760 3391 2816
rect 0 2758 3391 2760
rect 0 2728 800 2758
rect 3325 2755 3391 2758
rect 38009 2818 38075 2821
rect 39200 2818 40000 2848
rect 38009 2816 40000 2818
rect 38009 2760 38014 2816
rect 38070 2760 40000 2816
rect 38009 2758 40000 2760
rect 38009 2755 38075 2758
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 39200 2728 40000 2758
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 0 2138 800 2168
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
rect 2865 2138 2931 2141
rect 0 2136 2931 2138
rect 0 2080 2870 2136
rect 2926 2080 2931 2136
rect 0 2078 2931 2080
rect 0 2048 800 2078
rect 2865 2075 2931 2078
rect 36813 2138 36879 2141
rect 39200 2138 40000 2168
rect 36813 2136 40000 2138
rect 36813 2080 36818 2136
rect 36874 2080 40000 2136
rect 36813 2078 40000 2080
rect 36813 2075 36879 2078
rect 39200 2048 40000 2078
rect 0 1458 800 1488
rect 2773 1458 2839 1461
rect 0 1456 2839 1458
rect 0 1400 2778 1456
rect 2834 1400 2839 1456
rect 0 1398 2839 1400
rect 0 1368 800 1398
rect 2773 1395 2839 1398
rect 35893 1458 35959 1461
rect 39200 1458 40000 1488
rect 35893 1456 40000 1458
rect 35893 1400 35898 1456
rect 35954 1400 40000 1456
rect 35893 1398 40000 1400
rect 35893 1395 35959 1398
rect 39200 1368 40000 1398
rect 0 778 800 808
rect 2957 778 3023 781
rect 0 776 3023 778
rect 0 720 2962 776
rect 3018 720 3023 776
rect 0 718 3023 720
rect 0 688 800 718
rect 2957 715 3023 718
rect 36445 778 36511 781
rect 39200 778 40000 808
rect 36445 776 40000 778
rect 36445 720 36450 776
rect 36506 720 40000 776
rect 36445 718 40000 720
rect 36445 715 36511 718
rect 39200 688 40000 718
rect 37641 98 37707 101
rect 39200 98 40000 128
rect 37641 96 40000 98
rect 37641 40 37646 96
rect 37702 40 40000 96
rect 37641 38 40000 40
rect 37641 35 37707 38
rect 39200 8 40000 38
<< via3 >>
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 47360 4528 47376
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 46816 19888 47376
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 47360 35248 47376
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 26128 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__110__A
timestamp 1649977179
transform 1 0 18584 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A0
timestamp 1649977179
transform 1 0 9660 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A1
timestamp 1649977179
transform -1 0 11684 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__S
timestamp 1649977179
transform 1 0 11040 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A1
timestamp 1649977179
transform -1 0 24564 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__S
timestamp 1649977179
transform 1 0 23552 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A0
timestamp 1649977179
transform 1 0 21804 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A1
timestamp 1649977179
transform -1 0 21436 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__S
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A1
timestamp 1649977179
transform 1 0 22632 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__S
timestamp 1649977179
transform 1 0 21160 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__A0
timestamp 1649977179
transform -1 0 26220 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__119__S
timestamp 1649977179
transform 1 0 25484 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__121__S
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__A0
timestamp 1649977179
transform 1 0 12696 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__S
timestamp 1649977179
transform 1 0 12328 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__A0
timestamp 1649977179
transform -1 0 10396 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__S
timestamp 1649977179
transform 1 0 9844 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__A1
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__S
timestamp 1649977179
transform -1 0 26496 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A0
timestamp 1649977179
transform 1 0 25576 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__A1
timestamp 1649977179
transform -1 0 23920 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__129__S
timestamp 1649977179
transform 1 0 24196 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__A
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__A1
timestamp 1649977179
transform 1 0 14352 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__S
timestamp 1649977179
transform 1 0 15364 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__S
timestamp 1649977179
transform 1 0 2760 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__S
timestamp 1649977179
transform -1 0 12972 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__S
timestamp 1649977179
transform 1 0 16008 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A0
timestamp 1649977179
transform 1 0 8740 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__S
timestamp 1649977179
transform 1 0 9292 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__S
timestamp 1649977179
transform 1 0 16008 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__S
timestamp 1649977179
transform 1 0 27324 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A1
timestamp 1649977179
transform -1 0 6532 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__S
timestamp 1649977179
transform 1 0 5888 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__A0
timestamp 1649977179
transform -1 0 36800 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__148__S
timestamp 1649977179
transform 1 0 37168 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A0
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A1
timestamp 1649977179
transform 1 0 24380 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__S
timestamp 1649977179
transform 1 0 22448 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__152__A
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__A0
timestamp 1649977179
transform 1 0 28060 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__A1
timestamp 1649977179
transform 1 0 29808 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__S
timestamp 1649977179
transform 1 0 28428 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A0
timestamp 1649977179
transform -1 0 23276 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A1
timestamp 1649977179
transform 1 0 23644 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__S
timestamp 1649977179
transform 1 0 21712 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A0
timestamp 1649977179
transform 1 0 28704 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__S
timestamp 1649977179
transform 1 0 26956 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A0
timestamp 1649977179
transform 1 0 23644 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A1
timestamp 1649977179
transform 1 0 23460 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__S
timestamp 1649977179
transform 1 0 21896 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__A0
timestamp 1649977179
transform 1 0 20792 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__A1
timestamp 1649977179
transform 1 0 20608 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__S
timestamp 1649977179
transform 1 0 20608 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A0
timestamp 1649977179
transform -1 0 27600 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A1
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__S
timestamp 1649977179
transform 1 0 27784 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__165__A1
timestamp 1649977179
transform 1 0 25300 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__165__S
timestamp 1649977179
transform 1 0 24380 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__A0
timestamp 1649977179
transform 1 0 20240 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__A1
timestamp 1649977179
transform -1 0 19780 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__S
timestamp 1649977179
transform 1 0 20792 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__A0
timestamp 1649977179
transform 1 0 27508 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__A1
timestamp 1649977179
transform 1 0 29900 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__S
timestamp 1649977179
transform 1 0 27876 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__171__A0
timestamp 1649977179
transform 1 0 20240 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__171__A1
timestamp 1649977179
transform -1 0 18768 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__171__S
timestamp 1649977179
transform -1 0 19320 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__A
timestamp 1649977179
transform 1 0 19044 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A0
timestamp 1649977179
transform 1 0 23644 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__A1
timestamp 1649977179
transform 1 0 23276 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__S
timestamp 1649977179
transform 1 0 20608 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__A0
timestamp 1649977179
transform -1 0 18768 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__A1
timestamp 1649977179
transform -1 0 19136 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__S
timestamp 1649977179
transform 1 0 19504 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__A0
timestamp 1649977179
transform 1 0 18584 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__A1
timestamp 1649977179
transform 1 0 21160 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__178__S
timestamp 1649977179
transform 1 0 19688 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__A0
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__A1
timestamp 1649977179
transform -1 0 12604 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__180__S
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__A0
timestamp 1649977179
transform 1 0 23460 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__A1
timestamp 1649977179
transform -1 0 21988 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__182__S
timestamp 1649977179
transform 1 0 22356 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__A0
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__184__S
timestamp 1649977179
transform 1 0 25116 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A0
timestamp 1649977179
transform 1 0 14812 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__A1
timestamp 1649977179
transform 1 0 13064 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__186__S
timestamp 1649977179
transform 1 0 14444 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A0
timestamp 1649977179
transform 1 0 22908 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__A1
timestamp 1649977179
transform 1 0 23644 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__S
timestamp 1649977179
transform 1 0 23092 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A0
timestamp 1649977179
transform 1 0 19688 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__A1
timestamp 1649977179
transform -1 0 22908 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__190__S
timestamp 1649977179
transform 1 0 19596 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A0
timestamp 1649977179
transform 1 0 20240 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__A1
timestamp 1649977179
transform 1 0 20056 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__192__S
timestamp 1649977179
transform 1 0 20056 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__194__A
timestamp 1649977179
transform 1 0 17480 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__A0
timestamp 1649977179
transform 1 0 26312 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__195__S
timestamp 1649977179
transform 1 0 26772 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__A0
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__A1
timestamp 1649977179
transform 1 0 21620 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__197__S
timestamp 1649977179
transform 1 0 23368 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__A0
timestamp 1649977179
transform 1 0 24932 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__A1
timestamp 1649977179
transform -1 0 20056 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__S
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__A0
timestamp 1649977179
transform 1 0 23368 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__A1
timestamp 1649977179
transform -1 0 24104 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__201__S
timestamp 1649977179
transform 1 0 22816 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__A0
timestamp 1649977179
transform -1 0 28152 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__A1
timestamp 1649977179
transform -1 0 27140 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__S
timestamp 1649977179
transform -1 0 27140 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__A1
timestamp 1649977179
transform -1 0 13984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__205__S
timestamp 1649977179
transform 1 0 15548 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__A0
timestamp 1649977179
transform -1 0 23920 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__A1
timestamp 1649977179
transform -1 0 25300 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__207__S
timestamp 1649977179
transform -1 0 25852 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__A0
timestamp 1649977179
transform -1 0 26496 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__S
timestamp 1649977179
transform 1 0 26772 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__S
timestamp 1649977179
transform 1 0 18400 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__S
timestamp 1649977179
transform 1 0 24380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__A0
timestamp 1649977179
transform -1 0 14812 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__215__S
timestamp 1649977179
transform 1 0 14260 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__S
timestamp 1649977179
transform -1 0 26496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A0
timestamp 1649977179
transform -1 0 5520 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__S
timestamp 1649977179
transform 1 0 4968 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A0
timestamp 1649977179
transform 1 0 3772 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__S
timestamp 1649977179
transform 1 0 5152 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__224__S
timestamp 1649977179
transform 1 0 4968 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__A1
timestamp 1649977179
transform 1 0 25116 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__226__S
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__A0
timestamp 1649977179
transform 1 0 5428 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__228__S
timestamp 1649977179
transform 1 0 7176 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__230__S
timestamp 1649977179
transform 1 0 4968 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__232__S
timestamp 1649977179
transform -1 0 27968 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__234__S
timestamp 1649977179
transform -1 0 27048 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__A1
timestamp 1649977179
transform -1 0 5152 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__236__S
timestamp 1649977179
transform 1 0 4600 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__A1
timestamp 1649977179
transform -1 0 4232 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__238__S
timestamp 1649977179
transform -1 0 3956 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__A0
timestamp 1649977179
transform -1 0 7268 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__240__S
timestamp 1649977179
transform 1 0 6900 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__242__S
timestamp 1649977179
transform 1 0 2760 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__244__A
timestamp 1649977179
transform 1 0 25484 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A0
timestamp 1649977179
transform -1 0 32660 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__A1
timestamp 1649977179
transform 1 0 33856 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__S
timestamp 1649977179
transform 1 0 32844 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__A0
timestamp 1649977179
transform 1 0 32476 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__247__S
timestamp 1649977179
transform 1 0 32844 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__A0
timestamp 1649977179
transform -1 0 14352 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__249__S
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__A0
timestamp 1649977179
transform -1 0 30452 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__251__S
timestamp 1649977179
transform 1 0 30452 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__A1
timestamp 1649977179
transform 1 0 32936 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__253__S
timestamp 1649977179
transform 1 0 33304 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__A1
timestamp 1649977179
transform 1 0 32844 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__255__S
timestamp 1649977179
transform 1 0 33212 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__A0
timestamp 1649977179
transform 1 0 19780 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__257__S
timestamp 1649977179
transform 1 0 21160 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__A0
timestamp 1649977179
transform 1 0 17848 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__259__S
timestamp 1649977179
transform 1 0 17480 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__A0
timestamp 1649977179
transform -1 0 33396 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__A1
timestamp 1649977179
transform -1 0 35144 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__261__S
timestamp 1649977179
transform 1 0 33580 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__A0
timestamp 1649977179
transform -1 0 19412 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__A1
timestamp 1649977179
transform -1 0 19964 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__263__S
timestamp 1649977179
transform 1 0 20148 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A0
timestamp 1649977179
transform 1 0 21160 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__A1
timestamp 1649977179
transform 1 0 23092 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__265__S
timestamp 1649977179
transform -1 0 23644 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__A1
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__267__S
timestamp 1649977179
transform 1 0 14536 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__A1
timestamp 1649977179
transform -1 0 7820 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__269__S
timestamp 1649977179
transform 1 0 8188 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__A1
timestamp 1649977179
transform -1 0 17296 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__271__S
timestamp 1649977179
transform -1 0 17112 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__273__S
timestamp 1649977179
transform 1 0 34500 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__A0
timestamp 1649977179
transform -1 0 11040 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__275__S
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__A0
timestamp 1649977179
transform -1 0 20976 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__A1
timestamp 1649977179
transform 1 0 23092 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__277__S
timestamp 1649977179
transform 1 0 22540 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__A
timestamp 1649977179
transform -1 0 21896 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__B
timestamp 1649977179
transform 1 0 23276 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__279__C_N
timestamp 1649977179
transform 1 0 23092 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__A
timestamp 1649977179
transform -1 0 22540 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__B
timestamp 1649977179
transform -1 0 22540 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__C
timestamp 1649977179
transform 1 0 20884 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__280__D
timestamp 1649977179
transform 1 0 20884 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__A
timestamp 1649977179
transform -1 0 23092 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__B
timestamp 1649977179
transform 1 0 24012 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__C
timestamp 1649977179
transform 1 0 24564 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__281__D
timestamp 1649977179
transform -1 0 25300 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__A
timestamp 1649977179
transform -1 0 21436 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__B
timestamp 1649977179
transform -1 0 23460 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__C
timestamp 1649977179
transform -1 0 23276 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__283__D
timestamp 1649977179
transform 1 0 21804 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__A_N
timestamp 1649977179
transform -1 0 24012 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__B
timestamp 1649977179
transform -1 0 24564 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__284__C
timestamp 1649977179
transform -1 0 23460 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__A
timestamp 1649977179
transform -1 0 17664 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__B
timestamp 1649977179
transform -1 0 19412 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__C
timestamp 1649977179
transform -1 0 17112 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__286__D_N
timestamp 1649977179
transform 1 0 17848 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__A
timestamp 1649977179
transform 1 0 24932 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__C
timestamp 1649977179
transform 1 0 25852 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__287__D
timestamp 1649977179
transform -1 0 24564 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__291__B1
timestamp 1649977179
transform -1 0 24012 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__292__A
timestamp 1649977179
transform 1 0 22356 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__294__A_N
timestamp 1649977179
transform 1 0 22356 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__A1
timestamp 1649977179
transform 1 0 24380 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__296__S
timestamp 1649977179
transform -1 0 25484 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__298__A
timestamp 1649977179
transform 1 0 15640 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__299__A
timestamp 1649977179
transform 1 0 17296 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__300__A
timestamp 1649977179
transform -1 0 22632 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__301__A
timestamp 1649977179
transform 1 0 21252 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__306__CLK
timestamp 1649977179
transform -1 0 21988 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__307__CLK
timestamp 1649977179
transform 1 0 22540 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_i_clk_A
timestamp 1649977179
transform -1 0 14352 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 2852 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 9108 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 18308 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 35604 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 36800 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 2208 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 2208 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 6532 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 2208 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 21528 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 37444 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 35512 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 4324 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 2852 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 2852 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 26956 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 1564 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 1564 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 38180 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 11040 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 33856 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 5060 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 37536 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 13984 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 38180 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 11040 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 2852 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 37536 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 4876 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 37444 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 36800 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 37628 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 2852 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 37536 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 2208 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 2208 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 37536 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 37536 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 33580 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 2208 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 37536 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 37444 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 18768 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 35788 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 30544 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 37536 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 19412 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 5888 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 13064 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 29256 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 24104 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 36800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 37536 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 2208 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 6808 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 2208 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 35696 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 2852 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 5060 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 2208 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1649977179
transform -1 0 20056 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1649977179
transform -1 0 16836 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1649977179
transform -1 0 5612 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1649977179
transform -1 0 3312 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1649977179
transform -1 0 35144 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1649977179
transform -1 0 14996 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1649977179
transform -1 0 33028 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1649977179
transform -1 0 21344 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1649977179
transform -1 0 2116 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1649977179
transform -1 0 2208 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1649977179
transform -1 0 15732 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1649977179
transform -1 0 2208 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1649977179
transform -1 0 18124 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1649977179
transform -1 0 34868 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1649977179
transform -1 0 2668 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1649977179
transform -1 0 1748 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1649977179
transform -1 0 1564 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1649977179
transform -1 0 12604 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1649977179
transform -1 0 37536 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1649977179
transform -1 0 37444 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1649977179
transform -1 0 4508 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1649977179
transform -1 0 23276 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1649977179
transform -1 0 2208 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1649977179
transform -1 0 2208 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1649977179
transform -1 0 2852 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1649977179
transform -1 0 12880 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1649977179
transform -1 0 37444 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1649977179
transform -1 0 36156 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1649977179
transform -1 0 37536 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1649977179
transform -1 0 31832 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1649977179
transform -1 0 3312 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1649977179
transform -1 0 8740 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1649977179
transform -1 0 37536 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1649977179
transform -1 0 19596 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1649977179
transform -1 0 36800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1649977179
transform -1 0 1564 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1649977179
transform -1 0 32936 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input98_A
timestamp 1649977179
transform -1 0 2668 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input99_A
timestamp 1649977179
transform -1 0 7176 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input100_A
timestamp 1649977179
transform -1 0 37536 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input101_A
timestamp 1649977179
transform -1 0 2208 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input102_A
timestamp 1649977179
transform -1 0 34408 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input103_A
timestamp 1649977179
transform -1 0 36708 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input104_A
timestamp 1649977179
transform -1 0 1564 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input105_A
timestamp 1649977179
transform -1 0 3956 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input106_A
timestamp 1649977179
transform -1 0 29256 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input107_A
timestamp 1649977179
transform -1 0 37536 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input108_A
timestamp 1649977179
transform -1 0 38180 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input109_A
timestamp 1649977179
transform -1 0 29808 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input110_A
timestamp 1649977179
transform -1 0 36248 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input111_A
timestamp 1649977179
transform -1 0 2208 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input112_A
timestamp 1649977179
transform -1 0 11684 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input113_A
timestamp 1649977179
transform -1 0 2760 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input114_A
timestamp 1649977179
transform -1 0 36892 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input115_A
timestamp 1649977179
transform -1 0 38180 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input116_A
timestamp 1649977179
transform -1 0 24564 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input117_A
timestamp 1649977179
transform -1 0 37536 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input118_A
timestamp 1649977179
transform -1 0 3956 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input119_A
timestamp 1649977179
transform -1 0 5244 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input120_A
timestamp 1649977179
transform -1 0 1564 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input121_A
timestamp 1649977179
transform 1 0 1564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input122_A
timestamp 1649977179
transform -1 0 7452 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input123_A
timestamp 1649977179
transform -1 0 37536 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input124_A
timestamp 1649977179
transform -1 0 22724 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input125_A
timestamp 1649977179
transform -1 0 36340 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input126_A
timestamp 1649977179
transform -1 0 37444 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input127_A
timestamp 1649977179
transform -1 0 11684 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input128_A
timestamp 1649977179
transform -1 0 6348 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input129_A
timestamp 1649977179
transform -1 0 37536 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input130_A
timestamp 1649977179
transform -1 0 37444 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input131_A
timestamp 1649977179
transform -1 0 1748 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input132_A
timestamp 1649977179
transform -1 0 37536 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input133_A
timestamp 1649977179
transform -1 0 28060 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input134_A
timestamp 1649977179
transform -1 0 2760 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input135_A
timestamp 1649977179
transform -1 0 37536 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input136_A
timestamp 1649977179
transform -1 0 34224 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input137_A
timestamp 1649977179
transform -1 0 37444 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input138_A
timestamp 1649977179
transform -1 0 32476 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input139_A
timestamp 1649977179
transform -1 0 1564 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input140_A
timestamp 1649977179
transform -1 0 2208 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input141_A
timestamp 1649977179
transform -1 0 28612 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input142_A
timestamp 1649977179
transform -1 0 4324 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input143_A
timestamp 1649977179
transform -1 0 33488 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input144_A
timestamp 1649977179
transform -1 0 2208 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input145_A
timestamp 1649977179
transform -1 0 3312 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input146_A
timestamp 1649977179
transform -1 0 2760 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input147_A
timestamp 1649977179
transform -1 0 2208 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input148_A
timestamp 1649977179
transform -1 0 8096 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input149_A
timestamp 1649977179
transform -1 0 3772 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input150_A
timestamp 1649977179
transform -1 0 23276 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input151_A
timestamp 1649977179
transform -1 0 12328 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input152_A
timestamp 1649977179
transform -1 0 23828 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input153_A
timestamp 1649977179
transform -1 0 29716 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input154_A
timestamp 1649977179
transform -1 0 37536 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input155_A
timestamp 1649977179
transform -1 0 2208 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input156_A
timestamp 1649977179
transform -1 0 37536 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input157_A
timestamp 1649977179
transform -1 0 9384 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input158_A
timestamp 1649977179
transform -1 0 16836 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input159_A
timestamp 1649977179
transform -1 0 27508 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input160_A
timestamp 1649977179
transform -1 0 38180 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input161_A
timestamp 1649977179
transform -1 0 29072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input162_A
timestamp 1649977179
transform -1 0 25944 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input163_A
timestamp 1649977179
transform -1 0 25392 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input164_A
timestamp 1649977179
transform -1 0 2208 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input165_A
timestamp 1649977179
transform -1 0 3956 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input166_A
timestamp 1649977179
transform -1 0 32384 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input167_A
timestamp 1649977179
transform -1 0 2208 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input168_A
timestamp 1649977179
transform -1 0 2852 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input169_A
timestamp 1649977179
transform -1 0 37536 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output170_A
timestamp 1649977179
transform -1 0 1748 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output171_A
timestamp 1649977179
transform -1 0 37444 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output172_A
timestamp 1649977179
transform 1 0 5612 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output173_A
timestamp 1649977179
transform 1 0 2116 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output174_A
timestamp 1649977179
transform 1 0 9752 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output175_A
timestamp 1649977179
transform -1 0 37444 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output176_A
timestamp 1649977179
transform 1 0 16100 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output178_A
timestamp 1649977179
transform -1 0 37444 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output179_A
timestamp 1649977179
transform -1 0 34040 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output180_A
timestamp 1649977179
transform -1 0 2300 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output181_A
timestamp 1649977179
transform 1 0 3220 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output182_A
timestamp 1649977179
transform 1 0 8188 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output184_A
timestamp 1649977179
transform 1 0 27876 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output186_A
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output187_A
timestamp 1649977179
transform -1 0 37444 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output188_A
timestamp 1649977179
transform -1 0 10488 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output190_A
timestamp 1649977179
transform -1 0 2300 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output192_A
timestamp 1649977179
transform 1 0 30820 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output193_A
timestamp 1649977179
transform -1 0 2300 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output194_A
timestamp 1649977179
transform 1 0 2116 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output196_A
timestamp 1649977179
transform 1 0 2116 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output197_A
timestamp 1649977179
transform -1 0 2300 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output198_A
timestamp 1649977179
transform -1 0 17756 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output201_A
timestamp 1649977179
transform 1 0 2116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output205_A
timestamp 1649977179
transform 1 0 36156 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output206_A
timestamp 1649977179
transform 1 0 10120 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output213_A
timestamp 1649977179
transform 1 0 30912 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output215_A
timestamp 1649977179
transform 1 0 37260 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output216_A
timestamp 1649977179
transform 1 0 2116 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output217_A
timestamp 1649977179
transform 1 0 31464 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output218_A
timestamp 1649977179
transform 1 0 35972 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output222_A
timestamp 1649977179
transform 1 0 36248 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output224_A
timestamp 1649977179
transform 1 0 2116 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output226_A
timestamp 1649977179
transform -1 0 37444 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output230_A
timestamp 1649977179
transform -1 0 37444 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output234_A
timestamp 1649977179
transform 1 0 20516 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output235_A
timestamp 1649977179
transform 1 0 4876 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output238_A
timestamp 1649977179
transform -1 0 2300 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output239_A
timestamp 1649977179
transform -1 0 2300 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output240_A
timestamp 1649977179
transform 1 0 14260 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output241_A
timestamp 1649977179
transform 1 0 36708 0 1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output243_A
timestamp 1649977179
transform 1 0 34776 0 -1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output245_A
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output248_A
timestamp 1649977179
transform 1 0 37260 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output253_A
timestamp 1649977179
transform 1 0 37260 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output254_A
timestamp 1649977179
transform 1 0 35696 0 -1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output255_A
timestamp 1649977179
transform 1 0 37260 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output256_A
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output258_A
timestamp 1649977179
transform -1 0 37444 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2300 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2852 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47
timestamp 1649977179
transform 1 0 5428 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1649977179
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63
timestamp 1649977179
transform 1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_77
timestamp 1649977179
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_83
timestamp 1649977179
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_89
timestamp 1649977179
transform 1 0 9292 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105
timestamp 1649977179
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111
timestamp 1649977179
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_133
timestamp 1649977179
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_139
timestamp 1649977179
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_145 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14444 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_157
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1649977179
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_175
timestamp 1649977179
transform 1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189
timestamp 1649977179
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1649977179
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_201
timestamp 1649977179
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217
timestamp 1649977179
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1649977179
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_237
timestamp 1649977179
transform 1 0 22908 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_245
timestamp 1649977179
transform 1 0 23644 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1649977179
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_262
timestamp 1649977179
transform 1 0 25208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_270
timestamp 1649977179
transform 1 0 25944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1649977179
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_284
timestamp 1649977179
transform 1 0 27232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_291
timestamp 1649977179
transform 1 0 27876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_298
timestamp 1649977179
transform 1 0 28520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1649977179
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_321
timestamp 1649977179
transform 1 0 30636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_329
timestamp 1649977179
transform 1 0 31372 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_335
timestamp 1649977179
transform 1 0 31924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_347
timestamp 1649977179
transform 1 0 33028 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_357
timestamp 1649977179
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_363
timestamp 1649977179
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_371
timestamp 1649977179
transform 1 0 35236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_375
timestamp 1649977179
transform 1 0 35604 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_380
timestamp 1649977179
transform 1 0 36064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_388
timestamp 1649977179
transform 1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1649977179
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_3
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_7
timestamp 1649977179
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_23
timestamp 1649977179
transform 1 0 3220 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_30
timestamp 1649977179
transform 1 0 3864 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_36
timestamp 1649977179
transform 1 0 4416 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_41
timestamp 1649977179
transform 1 0 4876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_49
timestamp 1649977179
transform 1 0 5612 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1649977179
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1649977179
transform 1 0 6808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_73
timestamp 1649977179
transform 1 0 7820 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_76
timestamp 1649977179
transform 1 0 8096 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_83
timestamp 1649977179
transform 1 0 8740 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_87
timestamp 1649977179
transform 1 0 9108 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_90
timestamp 1649977179
transform 1 0 9384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1649977179
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_102
timestamp 1649977179
transform 1 0 10488 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1649977179
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_116
timestamp 1649977179
transform 1 0 11776 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_122
timestamp 1649977179
transform 1 0 12328 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_132
timestamp 1649977179
transform 1 0 13248 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_138
timestamp 1649977179
transform 1 0 13800 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_155
timestamp 1649977179
transform 1 0 15364 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_162
timestamp 1649977179
transform 1 0 16008 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_171
timestamp 1649977179
transform 1 0 16836 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_177
timestamp 1649977179
transform 1 0 17388 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_187
timestamp 1649977179
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_191
timestamp 1649977179
transform 1 0 18676 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_195
timestamp 1649977179
transform 1 0 19044 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_201
timestamp 1649977179
transform 1 0 19596 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_209
timestamp 1649977179
transform 1 0 20332 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_213
timestamp 1649977179
transform 1 0 20700 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_220
timestamp 1649977179
transform 1 0 21344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_229
timestamp 1649977179
transform 1 0 22172 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_235
timestamp 1649977179
transform 1 0 22724 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_251
timestamp 1649977179
transform 1 0 24196 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_264
timestamp 1649977179
transform 1 0 25392 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_271
timestamp 1649977179
transform 1 0 26036 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1649977179
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_284
timestamp 1649977179
transform 1 0 27232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_291
timestamp 1649977179
transform 1 0 27876 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_300
timestamp 1649977179
transform 1 0 28704 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_306
timestamp 1649977179
transform 1 0 29256 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_312
timestamp 1649977179
transform 1 0 29808 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_316
timestamp 1649977179
transform 1 0 30176 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_319
timestamp 1649977179
transform 1 0 30452 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1649977179
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_340
timestamp 1649977179
transform 1 0 32384 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_347
timestamp 1649977179
transform 1 0 33028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_354
timestamp 1649977179
transform 1 0 33672 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_363
timestamp 1649977179
transform 1 0 34500 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_372
timestamp 1649977179
transform 1 0 35328 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_380
timestamp 1649977179
transform 1 0 36064 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1649977179
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_1_393
timestamp 1649977179
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_399
timestamp 1649977179
transform 1 0 37812 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_13
timestamp 1649977179
transform 1 0 2300 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_20
timestamp 1649977179
transform 1 0 2944 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_2_32
timestamp 1649977179
transform 1 0 4048 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_40
timestamp 1649977179
transform 1 0 4784 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_43
timestamp 1649977179
transform 1 0 5060 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_51
timestamp 1649977179
transform 1 0 5796 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_57 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_69
timestamp 1649977179
transform 1 0 7452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_81
timestamp 1649977179
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_115
timestamp 1649977179
transform 1 0 11684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_127
timestamp 1649977179
transform 1 0 12788 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_135
timestamp 1649977179
transform 1 0 13524 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_145
timestamp 1649977179
transform 1 0 14444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_151
timestamp 1649977179
transform 1 0 14996 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_171
timestamp 1649977179
transform 1 0 16836 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_184
timestamp 1649977179
transform 1 0 18032 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_190
timestamp 1649977179
transform 1 0 18584 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_217
timestamp 1649977179
transform 1 0 21068 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_2_222
timestamp 1649977179
transform 1 0 21528 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_234
timestamp 1649977179
transform 1 0 22632 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_238
timestamp 1649977179
transform 1 0 23000 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_241
timestamp 1649977179
transform 1 0 23276 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_247
timestamp 1649977179
transform 1 0 23828 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1649977179
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_259
timestamp 1649977179
transform 1 0 24932 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_271
timestamp 1649977179
transform 1 0 26036 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_281
timestamp 1649977179
transform 1 0 26956 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_287
timestamp 1649977179
transform 1 0 27508 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_293
timestamp 1649977179
transform 1 0 28060 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_299
timestamp 1649977179
transform 1 0 28612 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1649977179
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_317
timestamp 1649977179
transform 1 0 30268 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_321
timestamp 1649977179
transform 1 0 30636 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_328
timestamp 1649977179
transform 1 0 31280 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_334
timestamp 1649977179
transform 1 0 31832 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_340
timestamp 1649977179
transform 1 0 32384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_346
timestamp 1649977179
transform 1 0 32936 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_352
timestamp 1649977179
transform 1 0 33488 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_358
timestamp 1649977179
transform 1 0 34040 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_367
timestamp 1649977179
transform 1 0 34868 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_375
timestamp 1649977179
transform 1 0 35604 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_379
timestamp 1649977179
transform 1 0 35972 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_387
timestamp 1649977179
transform 1 0 36708 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_395
timestamp 1649977179
transform 1 0 37444 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_403
timestamp 1649977179
transform 1 0 38180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_6
timestamp 1649977179
transform 1 0 1656 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1649977179
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_19
timestamp 1649977179
transform 1 0 2852 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_29
timestamp 1649977179
transform 1 0 3772 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_35
timestamp 1649977179
transform 1 0 4324 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_41
timestamp 1649977179
transform 1 0 4876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_53
timestamp 1649977179
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_155
timestamp 1649977179
transform 1 0 15364 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1649977179
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1649977179
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1649977179
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_249
timestamp 1649977179
transform 1 0 24012 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_255
timestamp 1649977179
transform 1 0 24564 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_267
timestamp 1649977179
transform 1 0 25668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_317
timestamp 1649977179
transform 1 0 30268 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_325
timestamp 1649977179
transform 1 0 31004 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_333
timestamp 1649977179
transform 1 0 31740 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_361
timestamp 1649977179
transform 1 0 34316 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_369
timestamp 1649977179
transform 1 0 35052 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_374
timestamp 1649977179
transform 1 0 35512 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_378
timestamp 1649977179
transform 1 0 35880 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_381
timestamp 1649977179
transform 1 0 36156 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_387
timestamp 1649977179
transform 1 0 36708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1649977179
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_395
timestamp 1649977179
transform 1 0 37444 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_403
timestamp 1649977179
transform 1 0 38180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_7
timestamp 1649977179
transform 1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_13
timestamp 1649977179
transform 1 0 2300 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_19
timestamp 1649977179
transform 1 0 2852 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_31
timestamp 1649977179
transform 1 0 3956 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_43
timestamp 1649977179
transform 1 0 5060 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_55
timestamp 1649977179
transform 1 0 6164 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_67
timestamp 1649977179
transform 1 0 7268 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_79
timestamp 1649977179
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_159
timestamp 1649977179
transform 1 0 15732 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_171
timestamp 1649977179
transform 1 0 16836 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_4_183
timestamp 1649977179
transform 1 0 17940 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1649977179
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1649977179
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1649977179
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1649977179
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1649977179
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1649977179
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1649977179
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1649977179
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1649977179
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1649977179
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1649977179
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1649977179
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_373
timestamp 1649977179
transform 1 0 35420 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_383
timestamp 1649977179
transform 1 0 36340 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_389
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_395
timestamp 1649977179
transform 1 0 37444 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_403
timestamp 1649977179
transform 1 0 38180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_6
timestamp 1649977179
transform 1 0 1656 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_12
timestamp 1649977179
transform 1 0 2208 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_18
timestamp 1649977179
transform 1 0 2760 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_24
timestamp 1649977179
transform 1 0 3312 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_36
timestamp 1649977179
transform 1 0 4416 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_48
timestamp 1649977179
transform 1 0 5520 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_52
timestamp 1649977179
transform 1 0 5888 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_5_248
timestamp 1649977179
transform 1 0 23920 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_260
timestamp 1649977179
transform 1 0 25024 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_272
timestamp 1649977179
transform 1 0 26128 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_5_276
timestamp 1649977179
transform 1 0 26496 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_285
timestamp 1649977179
transform 1 0 27324 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_297
timestamp 1649977179
transform 1 0 28428 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_309
timestamp 1649977179
transform 1 0 29532 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_321
timestamp 1649977179
transform 1 0 30636 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_333
timestamp 1649977179
transform 1 0 31740 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1649977179
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_385
timestamp 1649977179
transform 1 0 36524 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_388
timestamp 1649977179
transform 1 0 36800 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_395
timestamp 1649977179
transform 1 0 37444 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_403
timestamp 1649977179
transform 1 0 38180 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_7
timestamp 1649977179
transform 1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_13
timestamp 1649977179
transform 1 0 2300 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_19
timestamp 1649977179
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_49
timestamp 1649977179
transform 1 0 5612 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_62
timestamp 1649977179
transform 1 0 6808 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_68
timestamp 1649977179
transform 1 0 7360 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_80
timestamp 1649977179
transform 1 0 8464 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_130
timestamp 1649977179
transform 1 0 13064 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_138
timestamp 1649977179
transform 1 0 13800 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_145
timestamp 1649977179
transform 1 0 14444 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_157
timestamp 1649977179
transform 1 0 15548 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_169
timestamp 1649977179
transform 1 0 16652 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_181
timestamp 1649977179
transform 1 0 17756 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_193
timestamp 1649977179
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_245
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_248
timestamp 1649977179
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_262
timestamp 1649977179
transform 1 0 25208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_268
timestamp 1649977179
transform 1 0 25760 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_6_285
timestamp 1649977179
transform 1 0 27324 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_291
timestamp 1649977179
transform 1 0 27876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_303
timestamp 1649977179
transform 1 0 28980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1649977179
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1649977179
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1649977179
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1649977179
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1649977179
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1649977179
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1649977179
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_389
timestamp 1649977179
transform 1 0 36892 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_395
timestamp 1649977179
transform 1 0 37444 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_403
timestamp 1649977179
transform 1 0 38180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_7
timestamp 1649977179
transform 1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_13
timestamp 1649977179
transform 1 0 2300 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_25
timestamp 1649977179
transform 1 0 3404 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_37
timestamp 1649977179
transform 1 0 4508 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_49
timestamp 1649977179
transform 1 0 5612 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_122
timestamp 1649977179
transform 1 0 12328 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_7_128
timestamp 1649977179
transform 1 0 12880 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_7_143
timestamp 1649977179
transform 1 0 14260 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_249
timestamp 1649977179
transform 1 0 24012 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_7_253
timestamp 1649977179
transform 1 0 24380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_265
timestamp 1649977179
transform 1 0 25484 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_277
timestamp 1649977179
transform 1 0 26588 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1649977179
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1649977179
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1649977179
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1649977179
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1649977179
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_395
timestamp 1649977179
transform 1 0 37444 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_403
timestamp 1649977179
transform 1 0 38180 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_5
timestamp 1649977179
transform 1 0 1564 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_17
timestamp 1649977179
transform 1 0 2668 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_25
timestamp 1649977179
transform 1 0 3404 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_8_107
timestamp 1649977179
transform 1 0 10948 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_119
timestamp 1649977179
transform 1 0 12052 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_8_124
timestamp 1649977179
transform 1 0 12512 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_136
timestamp 1649977179
transform 1 0 13616 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_227
timestamp 1649977179
transform 1 0 21988 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1649977179
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1649977179
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1649977179
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1649977179
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1649977179
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1649977179
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1649977179
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1649977179
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1649977179
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1649977179
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1649977179
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1649977179
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1649977179
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1649977179
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_6
timestamp 1649977179
transform 1 0 1656 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_12
timestamp 1649977179
transform 1 0 2208 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_24
timestamp 1649977179
transform 1 0 3312 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_36
timestamp 1649977179
transform 1 0 4416 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_48
timestamp 1649977179
transform 1 0 5520 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1649977179
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_236
timestamp 1649977179
transform 1 0 22816 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_248
timestamp 1649977179
transform 1 0 23920 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_260
timestamp 1649977179
transform 1 0 25024 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_272
timestamp 1649977179
transform 1 0 26128 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1649977179
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1649977179
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1649977179
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1649977179
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1649977179
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1649977179
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1649977179
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1649977179
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_395
timestamp 1649977179
transform 1 0 37444 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_403
timestamp 1649977179
transform 1 0 38180 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_13
timestamp 1649977179
transform 1 0 2300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1649977179
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_175
timestamp 1649977179
transform 1 0 17204 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_187
timestamp 1649977179
transform 1 0 18308 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1649977179
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1649977179
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1649977179
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1649977179
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1649977179
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1649977179
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1649977179
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1649977179
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1649977179
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1649977179
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1649977179
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1649977179
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1649977179
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_389
timestamp 1649977179
transform 1 0 36892 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_10_397
timestamp 1649977179
transform 1 0 37628 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_403
timestamp 1649977179
transform 1 0 38180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_13
timestamp 1649977179
transform 1 0 2300 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_19
timestamp 1649977179
transform 1 0 2852 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_31
timestamp 1649977179
transform 1 0 3956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_43
timestamp 1649977179
transform 1 0 5060 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_164
timestamp 1649977179
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_171
timestamp 1649977179
transform 1 0 16836 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_183
timestamp 1649977179
transform 1 0 17940 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_195
timestamp 1649977179
transform 1 0 19044 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_207
timestamp 1649977179
transform 1 0 20148 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_219
timestamp 1649977179
transform 1 0 21252 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1649977179
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1649977179
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1649977179
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1649977179
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1649977179
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1649977179
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1649977179
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1649977179
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1649977179
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1649977179
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1649977179
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_395
timestamp 1649977179
transform 1 0 37444 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_403
timestamp 1649977179
transform 1 0 38180 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_7
timestamp 1649977179
transform 1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_13
timestamp 1649977179
transform 1 0 2300 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_25
timestamp 1649977179
transform 1 0 3404 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1649977179
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1649977179
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1649977179
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1649977179
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1649977179
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1649977179
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1649977179
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1649977179
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1649977179
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1649977179
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1649977179
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1649977179
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1649977179
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_389
timestamp 1649977179
transform 1 0 36892 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_403
timestamp 1649977179
transform 1 0 38180 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_145
timestamp 1649977179
transform 1 0 14444 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_148
timestamp 1649977179
transform 1 0 14720 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_171
timestamp 1649977179
transform 1 0 16836 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_183
timestamp 1649977179
transform 1 0 17940 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_195
timestamp 1649977179
transform 1 0 19044 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_207
timestamp 1649977179
transform 1 0 20148 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_219
timestamp 1649977179
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1649977179
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1649977179
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1649977179
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1649977179
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1649977179
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1649977179
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1649977179
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1649977179
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1649977179
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1649977179
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1649977179
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1649977179
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_403
timestamp 1649977179
transform 1 0 38180 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_6
timestamp 1649977179
transform 1 0 1656 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_12
timestamp 1649977179
transform 1 0 2208 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1649977179
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_109
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_117
timestamp 1649977179
transform 1 0 11868 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_14_123
timestamp 1649977179
transform 1 0 12420 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_135
timestamp 1649977179
transform 1 0 13524 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_159
timestamp 1649977179
transform 1 0 15732 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_163
timestamp 1649977179
transform 1 0 16100 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_175
timestamp 1649977179
transform 1 0 17204 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_187
timestamp 1649977179
transform 1 0 18308 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1649977179
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1649977179
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1649977179
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1649977179
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1649977179
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1649977179
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1649977179
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1649977179
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1649977179
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1649977179
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_389
timestamp 1649977179
transform 1 0 36892 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_395
timestamp 1649977179
transform 1 0 37444 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_403
timestamp 1649977179
transform 1 0 38180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_6
timestamp 1649977179
transform 1 0 1656 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_12
timestamp 1649977179
transform 1 0 2208 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_24
timestamp 1649977179
transform 1 0 3312 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_36
timestamp 1649977179
transform 1 0 4416 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_48
timestamp 1649977179
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_73
timestamp 1649977179
transform 1 0 7820 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_79
timestamp 1649977179
transform 1 0 8372 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_92
timestamp 1649977179
transform 1 0 9568 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_104
timestamp 1649977179
transform 1 0 10672 0 -1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_140
timestamp 1649977179
transform 1 0 13984 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1649977179
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_159
timestamp 1649977179
transform 1 0 15732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1649977179
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1649977179
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1649977179
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1649977179
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1649977179
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1649977179
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1649977179
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1649977179
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1649977179
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1649977179
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1649977179
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1649977179
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1649977179
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_396
timestamp 1649977179
transform 1 0 37536 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_403
timestamp 1649977179
transform 1 0 38180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_6
timestamp 1649977179
transform 1 0 1656 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_12
timestamp 1649977179
transform 1 0 2208 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1649977179
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1649977179
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1649977179
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1649977179
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1649977179
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1649977179
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1649977179
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1649977179
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1649977179
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1649977179
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1649977179
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1649977179
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1649977179
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1649977179
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1649977179
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_389
timestamp 1649977179
transform 1 0 36892 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_393
timestamp 1649977179
transform 1 0 37260 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_396
timestamp 1649977179
transform 1 0 37536 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_403
timestamp 1649977179
transform 1 0 38180 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_12
timestamp 1649977179
transform 1 0 2208 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_24
timestamp 1649977179
transform 1 0 3312 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_28
timestamp 1649977179
transform 1 0 3680 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_38
timestamp 1649977179
transform 1 0 4600 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_44
timestamp 1649977179
transform 1 0 5152 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_105
timestamp 1649977179
transform 1 0 10764 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1649977179
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_115
timestamp 1649977179
transform 1 0 11684 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_127
timestamp 1649977179
transform 1 0 12788 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_139
timestamp 1649977179
transform 1 0 13892 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_145
timestamp 1649977179
transform 1 0 14444 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_156
timestamp 1649977179
transform 1 0 15456 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1649977179
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1649977179
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1649977179
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1649977179
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1649977179
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1649977179
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1649977179
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1649977179
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1649977179
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1649977179
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1649977179
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_403
timestamp 1649977179
transform 1 0 38180 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_5
timestamp 1649977179
transform 1 0 1564 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_17
timestamp 1649977179
transform 1 0 2668 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1649977179
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_106
timestamp 1649977179
transform 1 0 10856 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_119
timestamp 1649977179
transform 1 0 12052 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_131
timestamp 1649977179
transform 1 0 13156 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1649977179
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1649977179
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1649977179
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1649977179
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1649977179
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1649977179
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1649977179
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1649977179
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1649977179
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1649977179
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1649977179
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1649977179
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_389
timestamp 1649977179
transform 1 0 36892 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_397
timestamp 1649977179
transform 1 0 37628 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_403
timestamp 1649977179
transform 1 0 38180 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_7
timestamp 1649977179
transform 1 0 1748 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_19
timestamp 1649977179
transform 1 0 2852 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_31
timestamp 1649977179
transform 1 0 3956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_43
timestamp 1649977179
transform 1 0 5060 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1649977179
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1649977179
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1649977179
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1649977179
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1649977179
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1649977179
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1649977179
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1649977179
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1649977179
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1649977179
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_361
timestamp 1649977179
transform 1 0 34316 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_19_365
timestamp 1649977179
transform 1 0 34684 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_377
timestamp 1649977179
transform 1 0 35788 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_389
timestamp 1649977179
transform 1 0 36892 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_403
timestamp 1649977179
transform 1 0 38180 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_6
timestamp 1649977179
transform 1 0 1656 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_12
timestamp 1649977179
transform 1 0 2208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_18
timestamp 1649977179
transform 1 0 2760 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_26
timestamp 1649977179
transform 1 0 3496 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_38
timestamp 1649977179
transform 1 0 4600 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_44
timestamp 1649977179
transform 1 0 5152 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_56
timestamp 1649977179
transform 1 0 6256 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_68
timestamp 1649977179
transform 1 0 7360 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_80
timestamp 1649977179
transform 1 0 8464 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1649977179
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1649977179
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1649977179
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_277
timestamp 1649977179
transform 1 0 26588 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_283
timestamp 1649977179
transform 1 0 27140 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_295
timestamp 1649977179
transform 1 0 28244 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1649977179
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1649977179
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1649977179
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1649977179
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_360
timestamp 1649977179
transform 1 0 34224 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_374
timestamp 1649977179
transform 1 0 35512 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_386
timestamp 1649977179
transform 1 0 36616 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_392
timestamp 1649977179
transform 1 0 37168 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_395
timestamp 1649977179
transform 1 0 37444 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_403
timestamp 1649977179
transform 1 0 38180 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_13
timestamp 1649977179
transform 1 0 2300 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_25
timestamp 1649977179
transform 1 0 3404 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_37
timestamp 1649977179
transform 1 0 4508 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_42
timestamp 1649977179
transform 1 0 4968 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_54
timestamp 1649977179
transform 1 0 6072 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1649977179
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1649977179
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1649977179
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_273
timestamp 1649977179
transform 1 0 26220 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1649977179
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_290
timestamp 1649977179
transform 1 0 27784 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_302
timestamp 1649977179
transform 1 0 28888 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_314
timestamp 1649977179
transform 1 0 29992 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_326
timestamp 1649977179
transform 1 0 31096 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_334
timestamp 1649977179
transform 1 0 31832 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_351
timestamp 1649977179
transform 1 0 33396 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_364
timestamp 1649977179
transform 1 0 34592 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_370
timestamp 1649977179
transform 1 0 35144 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_382
timestamp 1649977179
transform 1 0 36248 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_390
timestamp 1649977179
transform 1 0 36984 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_403
timestamp 1649977179
transform 1 0 38180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_7
timestamp 1649977179
transform 1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_13
timestamp 1649977179
transform 1 0 2300 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_25
timestamp 1649977179
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1649977179
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_277
timestamp 1649977179
transform 1 0 26588 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_281
timestamp 1649977179
transform 1 0 26956 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_295
timestamp 1649977179
transform 1 0 28244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1649977179
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1649977179
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1649977179
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_345
timestamp 1649977179
transform 1 0 32844 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_355
timestamp 1649977179
transform 1 0 33764 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1649977179
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1649977179
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_389
timestamp 1649977179
transform 1 0 36892 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_403
timestamp 1649977179
transform 1 0 38180 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_43
timestamp 1649977179
transform 1 0 5060 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1649977179
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1649977179
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1649977179
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1649977179
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_287
timestamp 1649977179
transform 1 0 27508 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_300
timestamp 1649977179
transform 1 0 28704 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_312
timestamp 1649977179
transform 1 0 29808 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_324
timestamp 1649977179
transform 1 0 30912 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1649977179
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_23_361
timestamp 1649977179
transform 1 0 34316 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_23_367
timestamp 1649977179
transform 1 0 34868 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_379
timestamp 1649977179
transform 1 0 35972 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1649977179
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_393
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_403
timestamp 1649977179
transform 1 0 38180 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_5
timestamp 1649977179
transform 1 0 1564 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_17
timestamp 1649977179
transform 1 0 2668 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_25
timestamp 1649977179
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_24_166
timestamp 1649977179
transform 1 0 16376 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_178
timestamp 1649977179
transform 1 0 17480 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_190
timestamp 1649977179
transform 1 0 18584 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1649977179
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1649977179
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1649977179
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1649977179
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1649977179
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1649977179
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1649977179
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1649977179
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1649977179
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1649977179
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1649977179
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1649977179
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_389
timestamp 1649977179
transform 1 0 36892 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_393
timestamp 1649977179
transform 1 0 37260 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_396
timestamp 1649977179
transform 1 0 37536 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_403
timestamp 1649977179
transform 1 0 38180 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_6
timestamp 1649977179
transform 1 0 1656 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_12
timestamp 1649977179
transform 1 0 2208 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_24
timestamp 1649977179
transform 1 0 3312 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_36
timestamp 1649977179
transform 1 0 4416 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_48
timestamp 1649977179
transform 1 0 5520 0 -1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_141
timestamp 1649977179
transform 1 0 14076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_144
timestamp 1649977179
transform 1 0 14352 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_157
timestamp 1649977179
transform 1 0 15548 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_163
timestamp 1649977179
transform 1 0 16100 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1649977179
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1649977179
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1649977179
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_283
timestamp 1649977179
transform 1 0 27140 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_295
timestamp 1649977179
transform 1 0 28244 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_307
timestamp 1649977179
transform 1 0 29348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_319
timestamp 1649977179
transform 1 0 30452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_331
timestamp 1649977179
transform 1 0 31556 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1649977179
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1649977179
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1649977179
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1649977179
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1649977179
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1649977179
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_395
timestamp 1649977179
transform 1 0 37444 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_403
timestamp 1649977179
transform 1 0 38180 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_13
timestamp 1649977179
transform 1 0 2300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_25
timestamp 1649977179
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1649977179
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1649977179
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_263
timestamp 1649977179
transform 1 0 25300 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_276
timestamp 1649977179
transform 1 0 26496 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_283
timestamp 1649977179
transform 1 0 27140 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_295
timestamp 1649977179
transform 1 0 28244 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1649977179
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1649977179
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1649977179
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1649977179
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1649977179
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_377
timestamp 1649977179
transform 1 0 35788 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_385
timestamp 1649977179
transform 1 0 36524 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_388
timestamp 1649977179
transform 1 0 36800 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_395
timestamp 1649977179
transform 1 0 37444 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_402
timestamp 1649977179
transform 1 0 38088 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_406
timestamp 1649977179
transform 1 0 38456 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_6
timestamp 1649977179
transform 1 0 1656 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_12
timestamp 1649977179
transform 1 0 2208 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_24
timestamp 1649977179
transform 1 0 3312 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_36
timestamp 1649977179
transform 1 0 4416 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_27_40
timestamp 1649977179
transform 1 0 4784 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_52
timestamp 1649977179
transform 1 0 5888 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1649977179
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1649977179
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1649977179
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1649977179
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1649977179
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1649977179
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1649977179
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1649977179
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1649977179
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1649977179
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1649977179
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1649977179
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_385
timestamp 1649977179
transform 1 0 36524 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_388
timestamp 1649977179
transform 1 0 36800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_393
timestamp 1649977179
transform 1 0 37260 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_403
timestamp 1649977179
transform 1 0 38180 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_38
timestamp 1649977179
transform 1 0 4600 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_44
timestamp 1649977179
transform 1 0 5152 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_56
timestamp 1649977179
transform 1 0 6256 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_68
timestamp 1649977179
transform 1 0 7360 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1649977179
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_144
timestamp 1649977179
transform 1 0 14352 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_168
timestamp 1649977179
transform 1 0 16560 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_180
timestamp 1649977179
transform 1 0 17664 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1649977179
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1649977179
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1649977179
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_265
timestamp 1649977179
transform 1 0 25484 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_273
timestamp 1649977179
transform 1 0 26220 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_28_279
timestamp 1649977179
transform 1 0 26772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_291
timestamp 1649977179
transform 1 0 27876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_303
timestamp 1649977179
transform 1 0 28980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1649977179
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1649977179
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1649977179
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1649977179
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1649977179
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_377
timestamp 1649977179
transform 1 0 35788 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_385
timestamp 1649977179
transform 1 0 36524 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_388
timestamp 1649977179
transform 1 0 36800 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_394
timestamp 1649977179
transform 1 0 37352 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_403
timestamp 1649977179
transform 1 0 38180 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_7
timestamp 1649977179
transform 1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_13
timestamp 1649977179
transform 1 0 2300 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_25
timestamp 1649977179
transform 1 0 3404 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_37
timestamp 1649977179
transform 1 0 4508 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_49
timestamp 1649977179
transform 1 0 5612 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1649977179
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_263
timestamp 1649977179
transform 1 0 25300 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1649977179
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_283
timestamp 1649977179
transform 1 0 27140 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_295
timestamp 1649977179
transform 1 0 28244 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_307
timestamp 1649977179
transform 1 0 29348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_319
timestamp 1649977179
transform 1 0 30452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_331
timestamp 1649977179
transform 1 0 31556 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1649977179
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1649977179
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1649977179
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1649977179
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1649977179
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1649977179
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_396
timestamp 1649977179
transform 1 0 37536 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_403
timestamp 1649977179
transform 1 0 38180 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_7
timestamp 1649977179
transform 1 0 1748 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_19
timestamp 1649977179
transform 1 0 2852 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_217
timestamp 1649977179
transform 1 0 21068 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_30_230
timestamp 1649977179
transform 1 0 22264 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_242
timestamp 1649977179
transform 1 0 23368 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1649977179
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1649977179
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1649977179
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1649977179
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1649977179
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1649977179
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1649977179
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1649977179
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_347
timestamp 1649977179
transform 1 0 33028 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_355
timestamp 1649977179
transform 1 0 33764 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_358
timestamp 1649977179
transform 1 0 34040 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_389
timestamp 1649977179
transform 1 0 36892 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_397
timestamp 1649977179
transform 1 0 37628 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_403
timestamp 1649977179
transform 1 0 38180 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_7
timestamp 1649977179
transform 1 0 1748 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_19
timestamp 1649977179
transform 1 0 2852 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_23
timestamp 1649977179
transform 1 0 3220 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_121
timestamp 1649977179
transform 1 0 12236 0 -1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_31_127
timestamp 1649977179
transform 1 0 12788 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_139
timestamp 1649977179
transform 1 0 13892 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_151
timestamp 1649977179
transform 1 0 14996 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_163
timestamp 1649977179
transform 1 0 16100 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1649977179
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_235
timestamp 1649977179
transform 1 0 22724 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_241
timestamp 1649977179
transform 1 0 23276 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_247
timestamp 1649977179
transform 1 0 23828 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_259
timestamp 1649977179
transform 1 0 24932 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_271
timestamp 1649977179
transform 1 0 26036 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1649977179
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1649977179
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1649977179
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1649977179
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_343
timestamp 1649977179
transform 1 0 32660 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_356
timestamp 1649977179
transform 1 0 33856 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_363
timestamp 1649977179
transform 1 0 34500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_375
timestamp 1649977179
transform 1 0 35604 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_387
timestamp 1649977179
transform 1 0 36708 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1649977179
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1649977179
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_13
timestamp 1649977179
transform 1 0 2300 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_20
timestamp 1649977179
transform 1 0 2944 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_31
timestamp 1649977179
transform 1 0 3956 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_43
timestamp 1649977179
transform 1 0 5060 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_55
timestamp 1649977179
transform 1 0 6164 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_67
timestamp 1649977179
transform 1 0 7268 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_79
timestamp 1649977179
transform 1 0 8372 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_123
timestamp 1649977179
transform 1 0 12420 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1649977179
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_143
timestamp 1649977179
transform 1 0 14260 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_155
timestamp 1649977179
transform 1 0 15364 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_167
timestamp 1649977179
transform 1 0 16468 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_179
timestamp 1649977179
transform 1 0 17572 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_191
timestamp 1649977179
transform 1 0 18676 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_32_226
timestamp 1649977179
transform 1 0 21896 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_238
timestamp 1649977179
transform 1 0 23000 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_250
timestamp 1649977179
transform 1 0 24104 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1649977179
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1649977179
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1649977179
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1649977179
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1649977179
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_333
timestamp 1649977179
transform 1 0 31740 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_343
timestamp 1649977179
transform 1 0 32660 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_356
timestamp 1649977179
transform 1 0 33856 0 1 19584
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1649977179
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_389
timestamp 1649977179
transform 1 0 36892 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_395
timestamp 1649977179
transform 1 0 37444 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_403
timestamp 1649977179
transform 1 0 38180 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_5
timestamp 1649977179
transform 1 0 1564 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_11
timestamp 1649977179
transform 1 0 2116 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_28
timestamp 1649977179
transform 1 0 3680 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_34
timestamp 1649977179
transform 1 0 4232 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_46
timestamp 1649977179
transform 1 0 5336 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1649977179
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_33_67
timestamp 1649977179
transform 1 0 7268 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_79
timestamp 1649977179
transform 1 0 8372 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_91
timestamp 1649977179
transform 1 0 9476 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_103
timestamp 1649977179
transform 1 0 10580 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_121
timestamp 1649977179
transform 1 0 12236 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1649977179
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1649977179
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_225
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_237
timestamp 1649977179
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_249
timestamp 1649977179
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_261
timestamp 1649977179
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1649977179
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1649977179
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1649977179
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1649977179
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1649977179
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1649977179
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_347
timestamp 1649977179
transform 1 0 33028 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_363
timestamp 1649977179
transform 1 0 34500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_375
timestamp 1649977179
transform 1 0 35604 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_387
timestamp 1649977179
transform 1 0 36708 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1649977179
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1649977179
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_6
timestamp 1649977179
transform 1 0 1656 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_12
timestamp 1649977179
transform 1 0 2208 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_24
timestamp 1649977179
transform 1 0 3312 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_63
timestamp 1649977179
transform 1 0 6900 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_71
timestamp 1649977179
transform 1 0 7636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1649977179
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1649977179
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1649977179
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1649977179
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1649977179
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1649977179
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_221
timestamp 1649977179
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_233
timestamp 1649977179
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_245
timestamp 1649977179
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1649977179
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1649977179
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1649977179
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1649977179
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1649977179
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1649977179
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1649977179
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1649977179
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1649977179
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1649977179
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1649977179
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_389
timestamp 1649977179
transform 1 0 36892 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_393
timestamp 1649977179
transform 1 0 37260 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_396
timestamp 1649977179
transform 1 0 37536 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_403
timestamp 1649977179
transform 1 0 38180 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_13
timestamp 1649977179
transform 1 0 2300 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_25
timestamp 1649977179
transform 1 0 3404 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_37
timestamp 1649977179
transform 1 0 4508 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_49
timestamp 1649977179
transform 1 0 5612 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1649977179
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_65
timestamp 1649977179
transform 1 0 7084 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_77
timestamp 1649977179
transform 1 0 8188 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_89
timestamp 1649977179
transform 1 0 9292 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_101
timestamp 1649977179
transform 1 0 10396 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_109
timestamp 1649977179
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1649977179
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1649977179
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_205
timestamp 1649977179
transform 1 0 19964 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_209
timestamp 1649977179
transform 1 0 20332 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_213
timestamp 1649977179
transform 1 0 20700 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_217
timestamp 1649977179
transform 1 0 21068 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_220
timestamp 1649977179
transform 1 0 21344 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_237
timestamp 1649977179
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_249
timestamp 1649977179
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_261
timestamp 1649977179
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_273
timestamp 1649977179
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1649977179
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1649977179
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1649977179
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1649977179
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1649977179
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1649977179
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1649977179
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1649977179
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1649977179
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1649977179
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_403
timestamp 1649977179
transform 1 0 38180 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_6
timestamp 1649977179
transform 1 0 1656 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_12
timestamp 1649977179
transform 1 0 2208 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1649977179
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1649977179
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1649977179
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1649977179
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_97
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_105
timestamp 1649977179
transform 1 0 10764 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_36_110
timestamp 1649977179
transform 1 0 11224 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_122
timestamp 1649977179
transform 1 0 12328 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_134
timestamp 1649977179
transform 1 0 13432 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1649977179
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_177
timestamp 1649977179
transform 1 0 17388 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_180
timestamp 1649977179
transform 1 0 17664 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1649977179
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_205
timestamp 1649977179
transform 1 0 19964 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_218
timestamp 1649977179
transform 1 0 21160 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_224
timestamp 1649977179
transform 1 0 21712 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_227
timestamp 1649977179
transform 1 0 21988 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_233
timestamp 1649977179
transform 1 0 22540 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_239
timestamp 1649977179
transform 1 0 23092 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1649977179
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1649977179
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1649977179
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1649977179
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1649977179
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1649977179
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1649977179
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1649977179
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1649977179
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1649977179
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1649977179
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1649977179
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_389
timestamp 1649977179
transform 1 0 36892 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_393
timestamp 1649977179
transform 1 0 37260 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_396
timestamp 1649977179
transform 1 0 37536 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_403
timestamp 1649977179
transform 1 0 38180 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_6
timestamp 1649977179
transform 1 0 1656 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_12
timestamp 1649977179
transform 1 0 2208 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_24
timestamp 1649977179
transform 1 0 3312 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_36
timestamp 1649977179
transform 1 0 4416 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_48
timestamp 1649977179
transform 1 0 5520 0 -1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1649977179
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_95
timestamp 1649977179
transform 1 0 9844 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_108
timestamp 1649977179
transform 1 0 11040 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_115
timestamp 1649977179
transform 1 0 11684 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_127
timestamp 1649977179
transform 1 0 12788 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_139
timestamp 1649977179
transform 1 0 13892 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_151
timestamp 1649977179
transform 1 0 14996 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_163
timestamp 1649977179
transform 1 0 16100 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_178
timestamp 1649977179
transform 1 0 17480 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_184
timestamp 1649977179
transform 1 0 18032 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_37_192
timestamp 1649977179
transform 1 0 18768 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_198
timestamp 1649977179
transform 1 0 19320 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_204
timestamp 1649977179
transform 1 0 19872 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_210
timestamp 1649977179
transform 1 0 20424 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1649977179
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_227
timestamp 1649977179
transform 1 0 21988 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_231
timestamp 1649977179
transform 1 0 22356 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_238
timestamp 1649977179
transform 1 0 23000 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_245
timestamp 1649977179
transform 1 0 23644 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_251
timestamp 1649977179
transform 1 0 24196 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_257
timestamp 1649977179
transform 1 0 24748 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_263
timestamp 1649977179
transform 1 0 25300 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1649977179
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1649977179
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1649977179
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1649977179
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1649977179
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1649977179
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1649977179
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1649977179
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1649977179
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1649977179
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1649977179
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1649977179
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_403
timestamp 1649977179
transform 1 0 38180 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1649977179
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1649977179
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1649977179
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_107
timestamp 1649977179
transform 1 0 10948 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_119
timestamp 1649977179
transform 1 0 12052 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_131
timestamp 1649977179
transform 1 0 13156 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_147
timestamp 1649977179
transform 1 0 14628 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_169
timestamp 1649977179
transform 1 0 16652 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_181
timestamp 1649977179
transform 1 0 17756 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_189
timestamp 1649977179
transform 1 0 18492 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1649977179
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_206
timestamp 1649977179
transform 1 0 20056 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_219
timestamp 1649977179
transform 1 0 21252 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_225
timestamp 1649977179
transform 1 0 21804 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_238
timestamp 1649977179
transform 1 0 23000 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_244
timestamp 1649977179
transform 1 0 23552 0 1 22848
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_38_255
timestamp 1649977179
transform 1 0 24564 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_267
timestamp 1649977179
transform 1 0 25668 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_279
timestamp 1649977179
transform 1 0 26772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_293
timestamp 1649977179
transform 1 0 28060 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_297
timestamp 1649977179
transform 1 0 28428 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_301
timestamp 1649977179
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1649977179
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1649977179
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1649977179
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1649977179
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1649977179
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1649977179
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1649977179
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1649977179
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_403
timestamp 1649977179
transform 1 0 38180 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_7
timestamp 1649977179
transform 1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_13
timestamp 1649977179
transform 1 0 2300 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_25
timestamp 1649977179
transform 1 0 3404 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_37
timestamp 1649977179
transform 1 0 4508 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_49
timestamp 1649977179
transform 1 0 5612 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1649977179
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1649977179
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1649977179
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1649977179
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_129
timestamp 1649977179
transform 1 0 12972 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_132
timestamp 1649977179
transform 1 0 13248 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_145
timestamp 1649977179
transform 1 0 14444 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_151
timestamp 1649977179
transform 1 0 14996 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_163
timestamp 1649977179
transform 1 0 16100 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_177
timestamp 1649977179
transform 1 0 17388 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_180
timestamp 1649977179
transform 1 0 17664 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_195
timestamp 1649977179
transform 1 0 19044 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_209
timestamp 1649977179
transform 1 0 20332 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1649977179
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_234
timestamp 1649977179
transform 1 0 22632 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_238
timestamp 1649977179
transform 1 0 23000 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_249
timestamp 1649977179
transform 1 0 24012 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_255
timestamp 1649977179
transform 1 0 24564 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_261
timestamp 1649977179
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_273
timestamp 1649977179
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1649977179
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_289
timestamp 1649977179
transform 1 0 27692 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_302
timestamp 1649977179
transform 1 0 28888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_309
timestamp 1649977179
transform 1 0 29532 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_315
timestamp 1649977179
transform 1 0 30084 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_327
timestamp 1649977179
transform 1 0 31188 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1649977179
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1649977179
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1649977179
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1649977179
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1649977179
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1649977179
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_395
timestamp 1649977179
transform 1 0 37444 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_403
timestamp 1649977179
transform 1 0 38180 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_11
timestamp 1649977179
transform 1 0 2116 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_17
timestamp 1649977179
transform 1 0 2668 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_25
timestamp 1649977179
transform 1 0 3404 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1649977179
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1649977179
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1649977179
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1649977179
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1649977179
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1649977179
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1649977179
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1649977179
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1649977179
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_165
timestamp 1649977179
transform 1 0 16284 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_171
timestamp 1649977179
transform 1 0 16836 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_174
timestamp 1649977179
transform 1 0 17112 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_180
timestamp 1649977179
transform 1 0 17664 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_192
timestamp 1649977179
transform 1 0 18768 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_199
timestamp 1649977179
transform 1 0 19412 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_203
timestamp 1649977179
transform 1 0 19780 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_214
timestamp 1649977179
transform 1 0 20792 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_220
timestamp 1649977179
transform 1 0 21344 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_225
timestamp 1649977179
transform 1 0 21804 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_239
timestamp 1649977179
transform 1 0 23092 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1649977179
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_259
timestamp 1649977179
transform 1 0 24932 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_265
timestamp 1649977179
transform 1 0 25484 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_271
timestamp 1649977179
transform 1 0 26036 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_283
timestamp 1649977179
transform 1 0 27140 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_288
timestamp 1649977179
transform 1 0 27600 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_301
timestamp 1649977179
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1649977179
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_311
timestamp 1649977179
transform 1 0 29716 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_323
timestamp 1649977179
transform 1 0 30820 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_335
timestamp 1649977179
transform 1 0 31924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_347
timestamp 1649977179
transform 1 0 33028 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_359
timestamp 1649977179
transform 1 0 34132 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1649977179
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_389
timestamp 1649977179
transform 1 0 36892 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_397
timestamp 1649977179
transform 1 0 37628 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_403
timestamp 1649977179
transform 1 0 38180 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_6
timestamp 1649977179
transform 1 0 1656 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_12
timestamp 1649977179
transform 1 0 2208 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_24
timestamp 1649977179
transform 1 0 3312 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_36
timestamp 1649977179
transform 1 0 4416 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_48
timestamp 1649977179
transform 1 0 5520 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1649977179
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1649977179
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1649977179
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1649977179
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1649977179
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1649977179
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1649977179
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1649977179
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_184
timestamp 1649977179
transform 1 0 18032 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_198
timestamp 1649977179
transform 1 0 19320 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_206
timestamp 1649977179
transform 1 0 20056 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1649977179
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_228
timestamp 1649977179
transform 1 0 22080 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_241
timestamp 1649977179
transform 1 0 23276 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_254
timestamp 1649977179
transform 1 0 24472 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_41_271
timestamp 1649977179
transform 1 0 26036 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1649977179
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_289
timestamp 1649977179
transform 1 0 27692 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_292
timestamp 1649977179
transform 1 0 27968 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_304
timestamp 1649977179
transform 1 0 29072 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_316
timestamp 1649977179
transform 1 0 30176 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_328
timestamp 1649977179
transform 1 0 31280 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1649977179
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1649977179
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1649977179
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1649977179
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1649977179
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_396
timestamp 1649977179
transform 1 0 37536 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_403
timestamp 1649977179
transform 1 0 38180 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_11
timestamp 1649977179
transform 1 0 2116 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_23
timestamp 1649977179
transform 1 0 3220 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1649977179
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1649977179
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1649977179
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1649977179
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1649977179
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1649977179
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1649977179
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1649977179
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1649977179
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1649977179
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_177
timestamp 1649977179
transform 1 0 17388 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_190
timestamp 1649977179
transform 1 0 18584 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_42_206
timestamp 1649977179
transform 1 0 20056 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_214
timestamp 1649977179
transform 1 0 20792 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_227
timestamp 1649977179
transform 1 0 21988 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_241
timestamp 1649977179
transform 1 0 23276 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_247
timestamp 1649977179
transform 1 0 23828 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1649977179
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_255
timestamp 1649977179
transform 1 0 24564 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_261
timestamp 1649977179
transform 1 0 25116 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_267
timestamp 1649977179
transform 1 0 25668 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_281
timestamp 1649977179
transform 1 0 26956 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_293
timestamp 1649977179
transform 1 0 28060 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_42_305
timestamp 1649977179
transform 1 0 29164 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1649977179
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1649977179
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1649977179
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1649977179
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1649977179
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1649977179
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_389
timestamp 1649977179
transform 1 0 36892 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_393
timestamp 1649977179
transform 1 0 37260 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_396
timestamp 1649977179
transform 1 0 37536 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_403
timestamp 1649977179
transform 1 0 38180 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_7
timestamp 1649977179
transform 1 0 1748 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_19
timestamp 1649977179
transform 1 0 2852 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_31
timestamp 1649977179
transform 1 0 3956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_43
timestamp 1649977179
transform 1 0 5060 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1649977179
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1649977179
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1649977179
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1649977179
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1649977179
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1649977179
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1649977179
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1649977179
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1649977179
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1649977179
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1649977179
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_181
timestamp 1649977179
transform 1 0 17756 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_191
timestamp 1649977179
transform 1 0 18676 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_197
timestamp 1649977179
transform 1 0 19228 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_203
timestamp 1649977179
transform 1 0 19780 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_207
timestamp 1649977179
transform 1 0 20148 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_210
timestamp 1649977179
transform 1 0 20424 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_216
timestamp 1649977179
transform 1 0 20976 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_43_225
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_229
timestamp 1649977179
transform 1 0 22172 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_237
timestamp 1649977179
transform 1 0 22908 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_243
timestamp 1649977179
transform 1 0 23460 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1649977179
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1649977179
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_273
timestamp 1649977179
transform 1 0 26220 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1649977179
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_290
timestamp 1649977179
transform 1 0 27784 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_302
timestamp 1649977179
transform 1 0 28888 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_314
timestamp 1649977179
transform 1 0 29992 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_326
timestamp 1649977179
transform 1 0 31096 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_334
timestamp 1649977179
transform 1 0 31832 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1649977179
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1649977179
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1649977179
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1649977179
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1649977179
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1649977179
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_7
timestamp 1649977179
transform 1 0 1748 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_19
timestamp 1649977179
transform 1 0 2852 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1649977179
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1649977179
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1649977179
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1649977179
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1649977179
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1649977179
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1649977179
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1649977179
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1649977179
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1649977179
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1649977179
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1649977179
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1649977179
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_189
timestamp 1649977179
transform 1 0 18492 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1649977179
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_209
timestamp 1649977179
transform 1 0 20332 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_44_217
timestamp 1649977179
transform 1 0 21068 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_223
timestamp 1649977179
transform 1 0 21620 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_226
timestamp 1649977179
transform 1 0 21896 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_237
timestamp 1649977179
transform 1 0 22908 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_243
timestamp 1649977179
transform 1 0 23460 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1649977179
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1649977179
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_277
timestamp 1649977179
transform 1 0 26588 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_283
timestamp 1649977179
transform 1 0 27140 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_287
timestamp 1649977179
transform 1 0 27508 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_299
timestamp 1649977179
transform 1 0 28612 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1649977179
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1649977179
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1649977179
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1649977179
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1649977179
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1649977179
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1649977179
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_389
timestamp 1649977179
transform 1 0 36892 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_395
timestamp 1649977179
transform 1 0 37444 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_403
timestamp 1649977179
transform 1 0 38180 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_7
timestamp 1649977179
transform 1 0 1748 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_13
timestamp 1649977179
transform 1 0 2300 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_25
timestamp 1649977179
transform 1 0 3404 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_37
timestamp 1649977179
transform 1 0 4508 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_49
timestamp 1649977179
transform 1 0 5612 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1649977179
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1649977179
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1649977179
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1649977179
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1649977179
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1649977179
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1649977179
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1649977179
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1649977179
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1649977179
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1649977179
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1649977179
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_193
timestamp 1649977179
transform 1 0 18860 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_196
timestamp 1649977179
transform 1 0 19136 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_202
timestamp 1649977179
transform 1 0 19688 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_209
timestamp 1649977179
transform 1 0 20332 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_219
timestamp 1649977179
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1649977179
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_227
timestamp 1649977179
transform 1 0 21988 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_233
timestamp 1649977179
transform 1 0 22540 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_241
timestamp 1649977179
transform 1 0 23276 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_253
timestamp 1649977179
transform 1 0 24380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_265
timestamp 1649977179
transform 1 0 25484 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_277
timestamp 1649977179
transform 1 0 26588 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1649977179
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1649977179
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1649977179
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1649977179
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1649977179
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1649977179
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1649977179
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1649977179
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1649977179
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1649977179
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_396
timestamp 1649977179
transform 1 0 37536 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_403
timestamp 1649977179
transform 1 0 38180 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_6
timestamp 1649977179
transform 1 0 1656 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_12
timestamp 1649977179
transform 1 0 2208 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_24
timestamp 1649977179
transform 1 0 3312 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_41
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_48
timestamp 1649977179
transform 1 0 5520 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_60
timestamp 1649977179
transform 1 0 6624 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_72
timestamp 1649977179
transform 1 0 7728 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1649977179
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1649977179
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1649977179
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1649977179
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1649977179
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1649977179
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1649977179
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1649977179
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_189
timestamp 1649977179
transform 1 0 18492 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1649977179
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_201
timestamp 1649977179
transform 1 0 19596 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_211
timestamp 1649977179
transform 1 0 20516 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_217
timestamp 1649977179
transform 1 0 21068 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_227
timestamp 1649977179
transform 1 0 21988 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_233
timestamp 1649977179
transform 1 0 22540 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_239
timestamp 1649977179
transform 1 0 23092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1649977179
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1649977179
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1649977179
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1649977179
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1649977179
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1649977179
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1649977179
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1649977179
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1649977179
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1649977179
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1649977179
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1649977179
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_389
timestamp 1649977179
transform 1 0 36892 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_395
timestamp 1649977179
transform 1 0 37444 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_403
timestamp 1649977179
transform 1 0 38180 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_6
timestamp 1649977179
transform 1 0 1656 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_12
timestamp 1649977179
transform 1 0 2208 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_24
timestamp 1649977179
transform 1 0 3312 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_32
timestamp 1649977179
transform 1 0 4048 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_42
timestamp 1649977179
transform 1 0 4968 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_48
timestamp 1649977179
transform 1 0 5520 0 -1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1649977179
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1649977179
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1649977179
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1649977179
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1649977179
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1649977179
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1649977179
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1649977179
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1649977179
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1649977179
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1649977179
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_193
timestamp 1649977179
transform 1 0 18860 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_199
timestamp 1649977179
transform 1 0 19412 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_205
timestamp 1649977179
transform 1 0 19964 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_218
timestamp 1649977179
transform 1 0 21160 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_235
timestamp 1649977179
transform 1 0 22724 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_241
timestamp 1649977179
transform 1 0 23276 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_247
timestamp 1649977179
transform 1 0 23828 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_259
timestamp 1649977179
transform 1 0 24932 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_47_274
timestamp 1649977179
transform 1 0 26312 0 -1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_283
timestamp 1649977179
transform 1 0 27140 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_295
timestamp 1649977179
transform 1 0 28244 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_307
timestamp 1649977179
transform 1 0 29348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_319
timestamp 1649977179
transform 1 0 30452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_331
timestamp 1649977179
transform 1 0 31556 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1649977179
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1649977179
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1649977179
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1649977179
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1649977179
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1649977179
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1649977179
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_395
timestamp 1649977179
transform 1 0 37444 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_403
timestamp 1649977179
transform 1 0 38180 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1649977179
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_41
timestamp 1649977179
transform 1 0 4876 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_44
timestamp 1649977179
transform 1 0 5152 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_56
timestamp 1649977179
transform 1 0 6256 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_68
timestamp 1649977179
transform 1 0 7360 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 1649977179
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1649977179
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1649977179
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1649977179
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1649977179
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1649977179
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1649977179
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1649977179
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1649977179
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1649977179
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1649977179
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_203
timestamp 1649977179
transform 1 0 19780 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_209
timestamp 1649977179
transform 1 0 20332 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_213
timestamp 1649977179
transform 1 0 20700 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_223
timestamp 1649977179
transform 1 0 21620 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_231
timestamp 1649977179
transform 1 0 22356 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_237
timestamp 1649977179
transform 1 0 22908 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_249
timestamp 1649977179
transform 1 0 24012 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1649977179
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1649977179
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1649977179
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1649977179
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1649977179
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1649977179
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1649977179
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_345
timestamp 1649977179
transform 1 0 32844 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_349
timestamp 1649977179
transform 1 0 33212 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_352
timestamp 1649977179
transform 1 0 33488 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1649977179
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1649977179
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1649977179
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1649977179
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_6
timestamp 1649977179
transform 1 0 1656 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_12
timestamp 1649977179
transform 1 0 2208 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_24
timestamp 1649977179
transform 1 0 3312 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_36
timestamp 1649977179
transform 1 0 4416 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_48
timestamp 1649977179
transform 1 0 5520 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1649977179
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1649977179
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1649977179
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1649977179
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1649977179
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1649977179
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1649977179
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_149
timestamp 1649977179
transform 1 0 14812 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1649977179
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_171
timestamp 1649977179
transform 1 0 16836 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_183
timestamp 1649977179
transform 1 0 17940 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_195
timestamp 1649977179
transform 1 0 19044 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_201
timestamp 1649977179
transform 1 0 19596 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_204
timestamp 1649977179
transform 1 0 19872 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_218
timestamp 1649977179
transform 1 0 21160 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_238
timestamp 1649977179
transform 1 0 23000 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_244
timestamp 1649977179
transform 1 0 23552 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_250
timestamp 1649977179
transform 1 0 24104 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_262
timestamp 1649977179
transform 1 0 25208 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_274
timestamp 1649977179
transform 1 0 26312 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_283
timestamp 1649977179
transform 1 0 27140 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_295
timestamp 1649977179
transform 1 0 28244 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_307
timestamp 1649977179
transform 1 0 29348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_319
timestamp 1649977179
transform 1 0 30452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_331
timestamp 1649977179
transform 1 0 31556 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1649977179
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_337
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_345
timestamp 1649977179
transform 1 0 32844 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_348
timestamp 1649977179
transform 1 0 33120 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1649977179
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1649977179
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1649977179
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1649977179
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_393
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_396
timestamp 1649977179
transform 1 0 37536 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_403
timestamp 1649977179
transform 1 0 38180 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_7
timestamp 1649977179
transform 1 0 1748 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_19
timestamp 1649977179
transform 1 0 2852 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1649977179
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1649977179
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1649977179
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1649977179
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1649977179
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1649977179
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1649977179
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1649977179
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1649977179
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1649977179
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1649977179
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1649977179
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1649977179
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1649977179
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1649977179
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1649977179
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_209
timestamp 1649977179
transform 1 0 20332 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_213
timestamp 1649977179
transform 1 0 20700 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_221
timestamp 1649977179
transform 1 0 21436 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_232
timestamp 1649977179
transform 1 0 22448 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_238
timestamp 1649977179
transform 1 0 23000 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1649977179
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_253
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_268
timestamp 1649977179
transform 1 0 25760 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_274
timestamp 1649977179
transform 1 0 26312 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_278
timestamp 1649977179
transform 1 0 26680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_288
timestamp 1649977179
transform 1 0 27600 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_294
timestamp 1649977179
transform 1 0 28152 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_306
timestamp 1649977179
transform 1 0 29256 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1649977179
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1649977179
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1649977179
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1649977179
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1649977179
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1649977179
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_368
timestamp 1649977179
transform 1 0 34960 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_380
timestamp 1649977179
transform 1 0 36064 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_392
timestamp 1649977179
transform 1 0 37168 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_396
timestamp 1649977179
transform 1 0 37536 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_403
timestamp 1649977179
transform 1 0 38180 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_7
timestamp 1649977179
transform 1 0 1748 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_13
timestamp 1649977179
transform 1 0 2300 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_25
timestamp 1649977179
transform 1 0 3404 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_37
timestamp 1649977179
transform 1 0 4508 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_49
timestamp 1649977179
transform 1 0 5612 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1649977179
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1649977179
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1649977179
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1649977179
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1649977179
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1649977179
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1649977179
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1649977179
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1649977179
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1649977179
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1649977179
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1649977179
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1649977179
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1649977179
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1649977179
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1649977179
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_225
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_235
timestamp 1649977179
transform 1 0 22724 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_239
timestamp 1649977179
transform 1 0 23092 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_244
timestamp 1649977179
transform 1 0 23552 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_257
timestamp 1649977179
transform 1 0 24748 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_263
timestamp 1649977179
transform 1 0 25300 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_269
timestamp 1649977179
transform 1 0 25852 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_277
timestamp 1649977179
transform 1 0 26588 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_283
timestamp 1649977179
transform 1 0 27140 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_290
timestamp 1649977179
transform 1 0 27784 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_302
timestamp 1649977179
transform 1 0 28888 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_314
timestamp 1649977179
transform 1 0 29992 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_326
timestamp 1649977179
transform 1 0 31096 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_334
timestamp 1649977179
transform 1 0 31832 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1649977179
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1649977179
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1649977179
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1649977179
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1649977179
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_393
timestamp 1649977179
transform 1 0 37260 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_403
timestamp 1649977179
transform 1 0 38180 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_5
timestamp 1649977179
transform 1 0 1564 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_17
timestamp 1649977179
transform 1 0 2668 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_25
timestamp 1649977179
transform 1 0 3404 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1649977179
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1649977179
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1649977179
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1649977179
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1649977179
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1649977179
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1649977179
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1649977179
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1649977179
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1649977179
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_141
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_145
timestamp 1649977179
transform 1 0 14444 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_149
timestamp 1649977179
transform 1 0 14812 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_176
timestamp 1649977179
transform 1 0 17296 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_188
timestamp 1649977179
transform 1 0 18400 0 1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1649977179
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_221
timestamp 1649977179
transform 1 0 21436 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_229
timestamp 1649977179
transform 1 0 22172 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_234
timestamp 1649977179
transform 1 0 22632 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_247
timestamp 1649977179
transform 1 0 23828 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1649977179
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_255
timestamp 1649977179
transform 1 0 24564 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_267
timestamp 1649977179
transform 1 0 25668 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_279
timestamp 1649977179
transform 1 0 26772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_291
timestamp 1649977179
transform 1 0 27876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_303
timestamp 1649977179
transform 1 0 28980 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1649977179
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1649977179
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1649977179
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1649977179
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1649977179
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1649977179
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1649977179
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_389
timestamp 1649977179
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_401
timestamp 1649977179
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_14
timestamp 1649977179
transform 1 0 2392 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_20
timestamp 1649977179
transform 1 0 2944 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_32
timestamp 1649977179
transform 1 0 4048 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_40
timestamp 1649977179
transform 1 0 4784 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_45
timestamp 1649977179
transform 1 0 5244 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_53
timestamp 1649977179
transform 1 0 5980 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1649977179
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1649977179
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1649977179
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1649977179
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1649977179
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1649977179
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_137
timestamp 1649977179
transform 1 0 13708 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_141
timestamp 1649977179
transform 1 0 14076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_163
timestamp 1649977179
transform 1 0 16100 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1649977179
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_177
timestamp 1649977179
transform 1 0 17388 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_189
timestamp 1649977179
transform 1 0 18492 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_201
timestamp 1649977179
transform 1 0 19596 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_207
timestamp 1649977179
transform 1 0 20148 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_210
timestamp 1649977179
transform 1 0 20424 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1649977179
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_53_227
timestamp 1649977179
transform 1 0 21988 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_237
timestamp 1649977179
transform 1 0 22908 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_243
timestamp 1649977179
transform 1 0 23460 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_249
timestamp 1649977179
transform 1 0 24012 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_255
timestamp 1649977179
transform 1 0 24564 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_267
timestamp 1649977179
transform 1 0 25668 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1649977179
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1649977179
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1649977179
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1649977179
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1649977179
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1649977179
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1649977179
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1649977179
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1649977179
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1649977179
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1649977179
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1649977179
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_13
timestamp 1649977179
transform 1 0 2300 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_20
timestamp 1649977179
transform 1 0 2944 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1649977179
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1649977179
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1649977179
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1649977179
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1649977179
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1649977179
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1649977179
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1649977179
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1649977179
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_141
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_149
timestamp 1649977179
transform 1 0 14812 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_154
timestamp 1649977179
transform 1 0 15272 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_160
timestamp 1649977179
transform 1 0 15824 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_168
timestamp 1649977179
transform 1 0 16560 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_172
timestamp 1649977179
transform 1 0 16928 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_178
timestamp 1649977179
transform 1 0 17480 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_192
timestamp 1649977179
transform 1 0 18768 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_197
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_205
timestamp 1649977179
transform 1 0 19964 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_208
timestamp 1649977179
transform 1 0 20240 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_221
timestamp 1649977179
transform 1 0 21436 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_227
timestamp 1649977179
transform 1 0 21988 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_54_243
timestamp 1649977179
transform 1 0 23460 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1649977179
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_255
timestamp 1649977179
transform 1 0 24564 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_267
timestamp 1649977179
transform 1 0 25668 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_279
timestamp 1649977179
transform 1 0 26772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_291
timestamp 1649977179
transform 1 0 27876 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_54_299
timestamp 1649977179
transform 1 0 28612 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1649977179
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1649977179
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1649977179
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1649977179
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1649977179
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1649977179
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1649977179
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_389
timestamp 1649977179
transform 1 0 36892 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_395
timestamp 1649977179
transform 1 0 37444 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_403
timestamp 1649977179
transform 1 0 38180 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_7
timestamp 1649977179
transform 1 0 1748 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_19
timestamp 1649977179
transform 1 0 2852 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_31
timestamp 1649977179
transform 1 0 3956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_43
timestamp 1649977179
transform 1 0 5060 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1649977179
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1649977179
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1649977179
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1649977179
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1649977179
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1649977179
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1649977179
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1649977179
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1649977179
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1649977179
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1649977179
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1649977179
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1649977179
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_205
timestamp 1649977179
transform 1 0 19964 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_208
timestamp 1649977179
transform 1 0 20240 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_216
timestamp 1649977179
transform 1 0 20976 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1649977179
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_55_234
timestamp 1649977179
transform 1 0 22632 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_249
timestamp 1649977179
transform 1 0 24012 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_255
timestamp 1649977179
transform 1 0 24564 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_267
timestamp 1649977179
transform 1 0 25668 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1649977179
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_295
timestamp 1649977179
transform 1 0 28244 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_308
timestamp 1649977179
transform 1 0 29440 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_314
timestamp 1649977179
transform 1 0 29992 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_326
timestamp 1649977179
transform 1 0 31096 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_334
timestamp 1649977179
transform 1 0 31832 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1649977179
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1649977179
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1649977179
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1649977179
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1649977179
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_55_393
timestamp 1649977179
transform 1 0 37260 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_396
timestamp 1649977179
transform 1 0 37536 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_403
timestamp 1649977179
transform 1 0 38180 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_6
timestamp 1649977179
transform 1 0 1656 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_12
timestamp 1649977179
transform 1 0 2208 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_24
timestamp 1649977179
transform 1 0 3312 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_41
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_49
timestamp 1649977179
transform 1 0 5612 0 1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_56_54
timestamp 1649977179
transform 1 0 6072 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_66
timestamp 1649977179
transform 1 0 7176 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_78
timestamp 1649977179
transform 1 0 8280 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1649977179
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1649977179
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1649977179
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1649977179
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1649977179
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1649977179
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_165
timestamp 1649977179
transform 1 0 16284 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_173
timestamp 1649977179
transform 1 0 17020 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_176
timestamp 1649977179
transform 1 0 17296 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_188
timestamp 1649977179
transform 1 0 18400 0 1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_209
timestamp 1649977179
transform 1 0 20332 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_217
timestamp 1649977179
transform 1 0 21068 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_56_221
timestamp 1649977179
transform 1 0 21436 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_230
timestamp 1649977179
transform 1 0 22264 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_240
timestamp 1649977179
transform 1 0 23184 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_246
timestamp 1649977179
transform 1 0 23736 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1649977179
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1649977179
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1649977179
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1649977179
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1649977179
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_312
timestamp 1649977179
transform 1 0 29808 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_324
timestamp 1649977179
transform 1 0 30912 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_336
timestamp 1649977179
transform 1 0 32016 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_348
timestamp 1649977179
transform 1 0 33120 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_360
timestamp 1649977179
transform 1 0 34224 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1649977179
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_389
timestamp 1649977179
transform 1 0 36892 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_393
timestamp 1649977179
transform 1 0 37260 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_396
timestamp 1649977179
transform 1 0 37536 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_403
timestamp 1649977179
transform 1 0 38180 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_6
timestamp 1649977179
transform 1 0 1656 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_12
timestamp 1649977179
transform 1 0 2208 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_24
timestamp 1649977179
transform 1 0 3312 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_36
timestamp 1649977179
transform 1 0 4416 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_42
timestamp 1649977179
transform 1 0 4968 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_52
timestamp 1649977179
transform 1 0 5888 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_59
timestamp 1649977179
transform 1 0 6532 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_71
timestamp 1649977179
transform 1 0 7636 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_83
timestamp 1649977179
transform 1 0 8740 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_95
timestamp 1649977179
transform 1 0 9844 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_107
timestamp 1649977179
transform 1 0 10948 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1649977179
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1649977179
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1649977179
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1649977179
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1649977179
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_169
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_174
timestamp 1649977179
transform 1 0 17112 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_187
timestamp 1649977179
transform 1 0 18308 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_199
timestamp 1649977179
transform 1 0 19412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_211
timestamp 1649977179
transform 1 0 20516 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_217
timestamp 1649977179
transform 1 0 21068 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_220
timestamp 1649977179
transform 1 0 21344 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_225
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_229
timestamp 1649977179
transform 1 0 22172 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_239
timestamp 1649977179
transform 1 0 23092 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_245
timestamp 1649977179
transform 1 0 23644 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_257
timestamp 1649977179
transform 1 0 24748 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_269
timestamp 1649977179
transform 1 0 25852 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_277
timestamp 1649977179
transform 1 0 26588 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1649977179
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1649977179
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1649977179
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1649977179
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1649977179
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1649977179
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1649977179
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1649977179
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1649977179
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1649977179
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_57_393
timestamp 1649977179
transform 1 0 37260 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_396
timestamp 1649977179
transform 1 0 37536 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_403
timestamp 1649977179
transform 1 0 38180 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_58_3
timestamp 1649977179
transform 1 0 1380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_14
timestamp 1649977179
transform 1 0 2392 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_20
timestamp 1649977179
transform 1 0 2944 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1649977179
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1649977179
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1649977179
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1649977179
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1649977179
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1649977179
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1649977179
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1649977179
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1649977179
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1649977179
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1649977179
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1649977179
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1649977179
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1649977179
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_209
timestamp 1649977179
transform 1 0 20332 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_215
timestamp 1649977179
transform 1 0 20884 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_226
timestamp 1649977179
transform 1 0 21896 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_230
timestamp 1649977179
transform 1 0 22264 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_234
timestamp 1649977179
transform 1 0 22632 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_238
timestamp 1649977179
transform 1 0 23000 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_241
timestamp 1649977179
transform 1 0 23276 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_249
timestamp 1649977179
transform 1 0 24012 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_267
timestamp 1649977179
transform 1 0 25668 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_273
timestamp 1649977179
transform 1 0 26220 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_58_286
timestamp 1649977179
transform 1 0 27416 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_298
timestamp 1649977179
transform 1 0 28520 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_306
timestamp 1649977179
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1649977179
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1649977179
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1649977179
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1649977179
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1649977179
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1649977179
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1649977179
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1649977179
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1649977179
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_59_13
timestamp 1649977179
transform 1 0 2300 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_19
timestamp 1649977179
transform 1 0 2852 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_31
timestamp 1649977179
transform 1 0 3956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_43
timestamp 1649977179
transform 1 0 5060 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1649977179
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1649977179
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1649977179
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1649977179
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1649977179
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1649977179
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1649977179
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1649977179
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1649977179
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1649977179
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1649977179
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1649977179
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1649977179
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1649977179
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1649977179
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1649977179
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_225
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_233
timestamp 1649977179
transform 1 0 22540 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_241
timestamp 1649977179
transform 1 0 23276 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_253
timestamp 1649977179
transform 1 0 24380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_265
timestamp 1649977179
transform 1 0 25484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_277
timestamp 1649977179
transform 1 0 26588 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_281
timestamp 1649977179
transform 1 0 26956 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_59_288
timestamp 1649977179
transform 1 0 27600 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_300
timestamp 1649977179
transform 1 0 28704 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_312
timestamp 1649977179
transform 1 0 29808 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_324
timestamp 1649977179
transform 1 0 30912 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1649977179
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1649977179
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1649977179
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1649977179
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1649977179
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1649977179
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_59_393
timestamp 1649977179
transform 1 0 37260 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_396
timestamp 1649977179
transform 1 0 37536 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_403
timestamp 1649977179
transform 1 0 38180 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_7
timestamp 1649977179
transform 1 0 1748 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_14
timestamp 1649977179
transform 1 0 2392 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_26
timestamp 1649977179
transform 1 0 3496 0 1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1649977179
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1649977179
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1649977179
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1649977179
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1649977179
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1649977179
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1649977179
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1649977179
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1649977179
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1649977179
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1649977179
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1649977179
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1649977179
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1649977179
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1649977179
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_209
timestamp 1649977179
transform 1 0 20332 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_217
timestamp 1649977179
transform 1 0 21068 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_221
timestamp 1649977179
transform 1 0 21436 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_227
timestamp 1649977179
transform 1 0 21988 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_237
timestamp 1649977179
transform 1 0 22908 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_243
timestamp 1649977179
transform 1 0 23460 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1649977179
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_253
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_261
timestamp 1649977179
transform 1 0 25116 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_273
timestamp 1649977179
transform 1 0 26220 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_285
timestamp 1649977179
transform 1 0 27324 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_297
timestamp 1649977179
transform 1 0 28428 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_305
timestamp 1649977179
transform 1 0 29164 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1649977179
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1649977179
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1649977179
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1649977179
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1649977179
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1649977179
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1649977179
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1649977179
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_401
timestamp 1649977179
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_7
timestamp 1649977179
transform 1 0 1748 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_13
timestamp 1649977179
transform 1 0 2300 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_25
timestamp 1649977179
transform 1 0 3404 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_37
timestamp 1649977179
transform 1 0 4508 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_49
timestamp 1649977179
transform 1 0 5612 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1649977179
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_57
timestamp 1649977179
transform 1 0 6348 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_66
timestamp 1649977179
transform 1 0 7176 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_79
timestamp 1649977179
transform 1 0 8372 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_85
timestamp 1649977179
transform 1 0 8924 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_91
timestamp 1649977179
transform 1 0 9476 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_103
timestamp 1649977179
transform 1 0 10580 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_111
timestamp 1649977179
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1649977179
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1649977179
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1649977179
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1649977179
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1649977179
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1649977179
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1649977179
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1649977179
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1649977179
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1649977179
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_225
timestamp 1649977179
transform 1 0 21804 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_228
timestamp 1649977179
transform 1 0 22080 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_61_241
timestamp 1649977179
transform 1 0 23276 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_249
timestamp 1649977179
transform 1 0 24012 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_259
timestamp 1649977179
transform 1 0 24932 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_61_265
timestamp 1649977179
transform 1 0 25484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_277
timestamp 1649977179
transform 1 0 26588 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1649977179
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1649977179
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1649977179
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1649977179
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1649977179
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1649977179
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1649977179
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1649977179
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1649977179
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1649977179
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1649977179
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_61_393
timestamp 1649977179
transform 1 0 37260 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_396
timestamp 1649977179
transform 1 0 37536 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_403
timestamp 1649977179
transform 1 0 38180 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_7
timestamp 1649977179
transform 1 0 1748 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_19
timestamp 1649977179
transform 1 0 2852 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1649977179
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1649977179
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1649977179
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1649977179
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1649977179
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1649977179
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1649977179
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1649977179
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1649977179
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1649977179
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1649977179
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1649977179
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1649977179
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1649977179
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1649977179
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1649977179
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_209
timestamp 1649977179
transform 1 0 20332 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_213
timestamp 1649977179
transform 1 0 20700 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_216
timestamp 1649977179
transform 1 0 20976 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_229
timestamp 1649977179
transform 1 0 22172 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_235
timestamp 1649977179
transform 1 0 22724 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_241
timestamp 1649977179
transform 1 0 23276 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_247
timestamp 1649977179
transform 1 0 23828 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1649977179
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_255
timestamp 1649977179
transform 1 0 24564 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_267
timestamp 1649977179
transform 1 0 25668 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_279
timestamp 1649977179
transform 1 0 26772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_291
timestamp 1649977179
transform 1 0 27876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_303
timestamp 1649977179
transform 1 0 28980 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1649977179
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1649977179
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1649977179
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1649977179
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1649977179
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1649977179
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1649977179
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1649977179
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1649977179
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_389
timestamp 1649977179
transform 1 0 36892 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_397
timestamp 1649977179
transform 1 0 37628 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_403
timestamp 1649977179
transform 1 0 38180 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1649977179
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1649977179
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1649977179
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1649977179
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1649977179
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1649977179
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1649977179
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1649977179
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_93
timestamp 1649977179
transform 1 0 9660 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_63_97
timestamp 1649977179
transform 1 0 10028 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_63_109
timestamp 1649977179
transform 1 0 11132 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1649977179
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_137
timestamp 1649977179
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_149
timestamp 1649977179
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1649977179
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1649977179
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1649977179
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1649977179
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1649977179
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1649977179
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_217
timestamp 1649977179
transform 1 0 21068 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_220
timestamp 1649977179
transform 1 0 21344 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_234
timestamp 1649977179
transform 1 0 22632 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_242
timestamp 1649977179
transform 1 0 23368 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_245
timestamp 1649977179
transform 1 0 23644 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_257
timestamp 1649977179
transform 1 0 24748 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_269
timestamp 1649977179
transform 1 0 25852 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_277
timestamp 1649977179
transform 1 0 26588 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1649977179
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1649977179
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1649977179
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1649977179
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1649977179
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1649977179
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1649977179
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1649977179
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1649977179
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1649977179
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1649977179
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1649977179
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_393
timestamp 1649977179
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_403
timestamp 1649977179
transform 1 0 38180 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_7
timestamp 1649977179
transform 1 0 1748 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_13
timestamp 1649977179
transform 1 0 2300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_25
timestamp 1649977179
transform 1 0 3404 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1649977179
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_53
timestamp 1649977179
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_65
timestamp 1649977179
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_77
timestamp 1649977179
transform 1 0 8188 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_83
timestamp 1649977179
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_95
timestamp 1649977179
transform 1 0 9844 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_101
timestamp 1649977179
transform 1 0 10396 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_113
timestamp 1649977179
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_125
timestamp 1649977179
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 1649977179
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_141
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_153
timestamp 1649977179
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_165
timestamp 1649977179
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_177
timestamp 1649977179
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1649977179
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1649977179
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1649977179
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_221
timestamp 1649977179
transform 1 0 21436 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_230
timestamp 1649977179
transform 1 0 22264 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_236
timestamp 1649977179
transform 1 0 22816 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_248
timestamp 1649977179
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1649977179
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1649977179
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_277
timestamp 1649977179
transform 1 0 26588 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_289
timestamp 1649977179
transform 1 0 27692 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1649977179
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1649977179
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_309
timestamp 1649977179
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_321
timestamp 1649977179
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_333
timestamp 1649977179
transform 1 0 31740 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_345
timestamp 1649977179
transform 1 0 32844 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_357
timestamp 1649977179
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_363
timestamp 1649977179
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1649977179
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1649977179
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_389
timestamp 1649977179
transform 1 0 36892 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_403
timestamp 1649977179
transform 1 0 38180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_13
timestamp 1649977179
transform 1 0 2300 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_65_19
timestamp 1649977179
transform 1 0 2852 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_31
timestamp 1649977179
transform 1 0 3956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_43
timestamp 1649977179
transform 1 0 5060 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1649977179
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_57
timestamp 1649977179
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_69
timestamp 1649977179
transform 1 0 7452 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_65_77
timestamp 1649977179
transform 1 0 8188 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_65_82
timestamp 1649977179
transform 1 0 8648 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_94
timestamp 1649977179
transform 1 0 9752 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_106
timestamp 1649977179
transform 1 0 10856 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_65_113
timestamp 1649977179
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_125
timestamp 1649977179
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_137
timestamp 1649977179
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_149
timestamp 1649977179
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1649977179
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1649977179
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_169
timestamp 1649977179
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_181
timestamp 1649977179
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_193
timestamp 1649977179
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_205
timestamp 1649977179
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_217
timestamp 1649977179
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_223
timestamp 1649977179
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_225
timestamp 1649977179
transform 1 0 21804 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_237
timestamp 1649977179
transform 1 0 22908 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_249
timestamp 1649977179
transform 1 0 24012 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_261
timestamp 1649977179
transform 1 0 25116 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_273
timestamp 1649977179
transform 1 0 26220 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1649977179
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_281
timestamp 1649977179
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_293
timestamp 1649977179
transform 1 0 28060 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_305
timestamp 1649977179
transform 1 0 29164 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_317
timestamp 1649977179
transform 1 0 30268 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_329
timestamp 1649977179
transform 1 0 31372 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_335
timestamp 1649977179
transform 1 0 31924 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_65_337
timestamp 1649977179
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_349
timestamp 1649977179
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_361
timestamp 1649977179
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_65_373
timestamp 1649977179
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1649977179
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1649977179
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_393
timestamp 1649977179
transform 1 0 37260 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_65_403
timestamp 1649977179
transform 1 0 38180 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_13
timestamp 1649977179
transform 1 0 2300 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_19
timestamp 1649977179
transform 1 0 2852 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_66_27
timestamp 1649977179
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_29
timestamp 1649977179
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_41
timestamp 1649977179
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_53
timestamp 1649977179
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_65
timestamp 1649977179
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1649977179
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1649977179
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_85
timestamp 1649977179
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_97
timestamp 1649977179
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_109
timestamp 1649977179
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_121
timestamp 1649977179
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1649977179
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1649977179
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_141
timestamp 1649977179
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_153
timestamp 1649977179
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_165
timestamp 1649977179
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_177
timestamp 1649977179
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_189
timestamp 1649977179
transform 1 0 18492 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_195
timestamp 1649977179
transform 1 0 19044 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_197
timestamp 1649977179
transform 1 0 19228 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_209
timestamp 1649977179
transform 1 0 20332 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_215
timestamp 1649977179
transform 1 0 20884 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_221
timestamp 1649977179
transform 1 0 21436 0 1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_66_227
timestamp 1649977179
transform 1 0 21988 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_239
timestamp 1649977179
transform 1 0 23092 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1649977179
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_253
timestamp 1649977179
transform 1 0 24380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_265
timestamp 1649977179
transform 1 0 25484 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_277
timestamp 1649977179
transform 1 0 26588 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_289
timestamp 1649977179
transform 1 0 27692 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_301
timestamp 1649977179
transform 1 0 28796 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_307
timestamp 1649977179
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_309
timestamp 1649977179
transform 1 0 29532 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_321
timestamp 1649977179
transform 1 0 30636 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_333
timestamp 1649977179
transform 1 0 31740 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_345
timestamp 1649977179
transform 1 0 32844 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_357
timestamp 1649977179
transform 1 0 33948 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_363
timestamp 1649977179
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_66_365
timestamp 1649977179
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_66_377
timestamp 1649977179
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_66_389
timestamp 1649977179
transform 1 0 36892 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_66_393
timestamp 1649977179
transform 1 0 37260 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_396
timestamp 1649977179
transform 1 0 37536 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_403
timestamp 1649977179
transform 1 0 38180 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_7
timestamp 1649977179
transform 1 0 1748 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_13
timestamp 1649977179
transform 1 0 2300 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_25
timestamp 1649977179
transform 1 0 3404 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_37
timestamp 1649977179
transform 1 0 4508 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_49
timestamp 1649977179
transform 1 0 5612 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1649977179
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_57
timestamp 1649977179
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_69
timestamp 1649977179
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_81
timestamp 1649977179
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_93
timestamp 1649977179
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1649977179
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1649977179
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_113
timestamp 1649977179
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_125
timestamp 1649977179
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_137
timestamp 1649977179
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_149
timestamp 1649977179
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1649977179
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1649977179
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_169
timestamp 1649977179
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_181
timestamp 1649977179
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_193
timestamp 1649977179
transform 1 0 18860 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_197
timestamp 1649977179
transform 1 0 19228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_219
timestamp 1649977179
transform 1 0 21252 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1649977179
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_228
timestamp 1649977179
transform 1 0 22080 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_67_234
timestamp 1649977179
transform 1 0 22632 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_246
timestamp 1649977179
transform 1 0 23736 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_258
timestamp 1649977179
transform 1 0 24840 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_270
timestamp 1649977179
transform 1 0 25944 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_278
timestamp 1649977179
transform 1 0 26680 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_67_281
timestamp 1649977179
transform 1 0 26956 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_293
timestamp 1649977179
transform 1 0 28060 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_305
timestamp 1649977179
transform 1 0 29164 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_317
timestamp 1649977179
transform 1 0 30268 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_329
timestamp 1649977179
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_335
timestamp 1649977179
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_67_337
timestamp 1649977179
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_349
timestamp 1649977179
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_361
timestamp 1649977179
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_67_373
timestamp 1649977179
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1649977179
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1649977179
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_395
timestamp 1649977179
transform 1 0 37444 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_403
timestamp 1649977179
transform 1 0 38180 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_5
timestamp 1649977179
transform 1 0 1564 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_17
timestamp 1649977179
transform 1 0 2668 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_25
timestamp 1649977179
transform 1 0 3404 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_68_29
timestamp 1649977179
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_41
timestamp 1649977179
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_53
timestamp 1649977179
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_65
timestamp 1649977179
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1649977179
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1649977179
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_85
timestamp 1649977179
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_97
timestamp 1649977179
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_109
timestamp 1649977179
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_121
timestamp 1649977179
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1649977179
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1649977179
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_141
timestamp 1649977179
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_153
timestamp 1649977179
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_165
timestamp 1649977179
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_177
timestamp 1649977179
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_189
timestamp 1649977179
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_195
timestamp 1649977179
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_197
timestamp 1649977179
transform 1 0 19228 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_204
timestamp 1649977179
transform 1 0 19872 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_68_229
timestamp 1649977179
transform 1 0 22172 0 1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_68_235
timestamp 1649977179
transform 1 0 22724 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_247
timestamp 1649977179
transform 1 0 23828 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_68_251
timestamp 1649977179
transform 1 0 24196 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_253
timestamp 1649977179
transform 1 0 24380 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_265
timestamp 1649977179
transform 1 0 25484 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_277
timestamp 1649977179
transform 1 0 26588 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_289
timestamp 1649977179
transform 1 0 27692 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_301
timestamp 1649977179
transform 1 0 28796 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_307
timestamp 1649977179
transform 1 0 29348 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_309
timestamp 1649977179
transform 1 0 29532 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_321
timestamp 1649977179
transform 1 0 30636 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_333
timestamp 1649977179
transform 1 0 31740 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_345
timestamp 1649977179
transform 1 0 32844 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_357
timestamp 1649977179
transform 1 0 33948 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_363
timestamp 1649977179
transform 1 0 34500 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_68_365
timestamp 1649977179
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_377
timestamp 1649977179
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_68_389
timestamp 1649977179
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_401
timestamp 1649977179
transform 1 0 37996 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_69_13
timestamp 1649977179
transform 1 0 2300 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_25
timestamp 1649977179
transform 1 0 3404 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_37
timestamp 1649977179
transform 1 0 4508 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_49
timestamp 1649977179
transform 1 0 5612 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1649977179
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_57
timestamp 1649977179
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_69
timestamp 1649977179
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_81
timestamp 1649977179
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_93
timestamp 1649977179
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1649977179
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1649977179
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_113
timestamp 1649977179
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_125
timestamp 1649977179
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_137
timestamp 1649977179
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_149
timestamp 1649977179
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1649977179
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1649977179
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_169
timestamp 1649977179
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_181
timestamp 1649977179
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_193
timestamp 1649977179
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_205
timestamp 1649977179
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_217
timestamp 1649977179
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1649977179
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_225
timestamp 1649977179
transform 1 0 21804 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_237
timestamp 1649977179
transform 1 0 22908 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_249
timestamp 1649977179
transform 1 0 24012 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_261
timestamp 1649977179
transform 1 0 25116 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1649977179
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1649977179
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_281
timestamp 1649977179
transform 1 0 26956 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_293
timestamp 1649977179
transform 1 0 28060 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_305
timestamp 1649977179
transform 1 0 29164 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_317
timestamp 1649977179
transform 1 0 30268 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_329
timestamp 1649977179
transform 1 0 31372 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1649977179
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_69_337
timestamp 1649977179
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_349
timestamp 1649977179
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_361
timestamp 1649977179
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_69_373
timestamp 1649977179
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1649977179
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1649977179
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_395
timestamp 1649977179
transform 1 0 37444 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_403
timestamp 1649977179
transform 1 0 38180 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_3
timestamp 1649977179
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_11
timestamp 1649977179
transform 1 0 2116 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_70_17
timestamp 1649977179
transform 1 0 2668 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_70_25
timestamp 1649977179
transform 1 0 3404 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_70_29
timestamp 1649977179
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_41
timestamp 1649977179
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_53
timestamp 1649977179
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_65
timestamp 1649977179
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1649977179
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1649977179
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_85
timestamp 1649977179
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_97
timestamp 1649977179
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_109
timestamp 1649977179
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_121
timestamp 1649977179
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1649977179
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1649977179
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_141
timestamp 1649977179
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_153
timestamp 1649977179
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_165
timestamp 1649977179
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_177
timestamp 1649977179
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1649977179
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1649977179
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_197
timestamp 1649977179
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_209
timestamp 1649977179
transform 1 0 20332 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_221
timestamp 1649977179
transform 1 0 21436 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_233
timestamp 1649977179
transform 1 0 22540 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_245
timestamp 1649977179
transform 1 0 23644 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1649977179
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_253
timestamp 1649977179
transform 1 0 24380 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_265
timestamp 1649977179
transform 1 0 25484 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_277
timestamp 1649977179
transform 1 0 26588 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_289
timestamp 1649977179
transform 1 0 27692 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_301
timestamp 1649977179
transform 1 0 28796 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_307
timestamp 1649977179
transform 1 0 29348 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_309
timestamp 1649977179
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_321
timestamp 1649977179
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_333
timestamp 1649977179
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_345
timestamp 1649977179
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1649977179
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1649977179
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_70_365
timestamp 1649977179
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_70_377
timestamp 1649977179
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_389
timestamp 1649977179
transform 1 0 36892 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_70_393
timestamp 1649977179
transform 1 0 37260 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_396
timestamp 1649977179
transform 1 0 37536 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_70_403
timestamp 1649977179
transform 1 0 38180 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_13
timestamp 1649977179
transform 1 0 2300 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_19
timestamp 1649977179
transform 1 0 2852 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_31
timestamp 1649977179
transform 1 0 3956 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_43
timestamp 1649977179
transform 1 0 5060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_55
timestamp 1649977179
transform 1 0 6164 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_57
timestamp 1649977179
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_69
timestamp 1649977179
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_81
timestamp 1649977179
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_93
timestamp 1649977179
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1649977179
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1649977179
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_113
timestamp 1649977179
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_125
timestamp 1649977179
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_137
timestamp 1649977179
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_149
timestamp 1649977179
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1649977179
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1649977179
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_71_169
timestamp 1649977179
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_181
timestamp 1649977179
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_193
timestamp 1649977179
transform 1 0 18860 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_205
timestamp 1649977179
transform 1 0 19964 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_71_213
timestamp 1649977179
transform 1 0 20700 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_216
timestamp 1649977179
transform 1 0 20976 0 -1 41344
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_71_225
timestamp 1649977179
transform 1 0 21804 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_237
timestamp 1649977179
transform 1 0 22908 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_249
timestamp 1649977179
transform 1 0 24012 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_261
timestamp 1649977179
transform 1 0 25116 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_273
timestamp 1649977179
transform 1 0 26220 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_279
timestamp 1649977179
transform 1 0 26772 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_283
timestamp 1649977179
transform 1 0 27140 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_296
timestamp 1649977179
transform 1 0 28336 0 -1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_71_302
timestamp 1649977179
transform 1 0 28888 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_314
timestamp 1649977179
transform 1 0 29992 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_326
timestamp 1649977179
transform 1 0 31096 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_334
timestamp 1649977179
transform 1 0 31832 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_71_337
timestamp 1649977179
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_349
timestamp 1649977179
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_361
timestamp 1649977179
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_71_373
timestamp 1649977179
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1649977179
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1649977179
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_71_393
timestamp 1649977179
transform 1 0 37260 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_71_396
timestamp 1649977179
transform 1 0 37536 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_403
timestamp 1649977179
transform 1 0 38180 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_3
timestamp 1649977179
transform 1 0 1380 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_11
timestamp 1649977179
transform 1 0 2116 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_23
timestamp 1649977179
transform 1 0 3220 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_27
timestamp 1649977179
transform 1 0 3588 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_29
timestamp 1649977179
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_41
timestamp 1649977179
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_53
timestamp 1649977179
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_65
timestamp 1649977179
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1649977179
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1649977179
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_85
timestamp 1649977179
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_97
timestamp 1649977179
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_109
timestamp 1649977179
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_121
timestamp 1649977179
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1649977179
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1649977179
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_141
timestamp 1649977179
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_153
timestamp 1649977179
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_165
timestamp 1649977179
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_177
timestamp 1649977179
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1649977179
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1649977179
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_197
timestamp 1649977179
transform 1 0 19228 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_72_209
timestamp 1649977179
transform 1 0 20332 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_72_214
timestamp 1649977179
transform 1 0 20792 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_227
timestamp 1649977179
transform 1 0 21988 0 1 41344
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_72_234
timestamp 1649977179
transform 1 0 22632 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_246
timestamp 1649977179
transform 1 0 23736 0 1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_72_253
timestamp 1649977179
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_265
timestamp 1649977179
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_277
timestamp 1649977179
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_289
timestamp 1649977179
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1649977179
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1649977179
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_309
timestamp 1649977179
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_321
timestamp 1649977179
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_333
timestamp 1649977179
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_345
timestamp 1649977179
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1649977179
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1649977179
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_72_365
timestamp 1649977179
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_72_377
timestamp 1649977179
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_389
timestamp 1649977179
transform 1 0 36892 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_393
timestamp 1649977179
transform 1 0 37260 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_396
timestamp 1649977179
transform 1 0 37536 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_403
timestamp 1649977179
transform 1 0 38180 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_73_3
timestamp 1649977179
transform 1 0 1380 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_7
timestamp 1649977179
transform 1 0 1748 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_19
timestamp 1649977179
transform 1 0 2852 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_27
timestamp 1649977179
transform 1 0 3588 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_31
timestamp 1649977179
transform 1 0 3956 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_43
timestamp 1649977179
transform 1 0 5060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1649977179
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_57
timestamp 1649977179
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_69
timestamp 1649977179
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_81
timestamp 1649977179
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_93
timestamp 1649977179
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1649977179
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1649977179
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_113
timestamp 1649977179
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_125
timestamp 1649977179
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_137
timestamp 1649977179
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_149
timestamp 1649977179
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1649977179
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1649977179
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_169
timestamp 1649977179
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_181
timestamp 1649977179
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_193
timestamp 1649977179
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_205
timestamp 1649977179
transform 1 0 19964 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_211
timestamp 1649977179
transform 1 0 20516 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_214
timestamp 1649977179
transform 1 0 20792 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_73_222
timestamp 1649977179
transform 1 0 21528 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_73_225
timestamp 1649977179
transform 1 0 21804 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_237
timestamp 1649977179
transform 1 0 22908 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_249
timestamp 1649977179
transform 1 0 24012 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_261
timestamp 1649977179
transform 1 0 25116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_273
timestamp 1649977179
transform 1 0 26220 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1649977179
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_281
timestamp 1649977179
transform 1 0 26956 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_73_286
timestamp 1649977179
transform 1 0 27416 0 -1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_73_292
timestamp 1649977179
transform 1 0 27968 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_304
timestamp 1649977179
transform 1 0 29072 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_316
timestamp 1649977179
transform 1 0 30176 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_328
timestamp 1649977179
transform 1 0 31280 0 -1 42432
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_73_337
timestamp 1649977179
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_349
timestamp 1649977179
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_361
timestamp 1649977179
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_73_373
timestamp 1649977179
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1649977179
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1649977179
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_73_393
timestamp 1649977179
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_405
timestamp 1649977179
transform 1 0 38364 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_6
timestamp 1649977179
transform 1 0 1656 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_12
timestamp 1649977179
transform 1 0 2208 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_24
timestamp 1649977179
transform 1 0 3312 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_74_29
timestamp 1649977179
transform 1 0 3772 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_40
timestamp 1649977179
transform 1 0 4784 0 1 42432
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_74_46
timestamp 1649977179
transform 1 0 5336 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_58
timestamp 1649977179
transform 1 0 6440 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_70
timestamp 1649977179
transform 1 0 7544 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_82
timestamp 1649977179
transform 1 0 8648 0 1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_74_85
timestamp 1649977179
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_97
timestamp 1649977179
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_109
timestamp 1649977179
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_121
timestamp 1649977179
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1649977179
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1649977179
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_141
timestamp 1649977179
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_153
timestamp 1649977179
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_165
timestamp 1649977179
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_177
timestamp 1649977179
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1649977179
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1649977179
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_197
timestamp 1649977179
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_209
timestamp 1649977179
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_221
timestamp 1649977179
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_233
timestamp 1649977179
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1649977179
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1649977179
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_253
timestamp 1649977179
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_265
timestamp 1649977179
transform 1 0 25484 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_74_277
timestamp 1649977179
transform 1 0 26588 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_74_285
timestamp 1649977179
transform 1 0 27324 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_295
timestamp 1649977179
transform 1 0 28244 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1649977179
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_309
timestamp 1649977179
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_321
timestamp 1649977179
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_333
timestamp 1649977179
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_345
timestamp 1649977179
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1649977179
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1649977179
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_74_365
timestamp 1649977179
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_74_377
timestamp 1649977179
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_389
timestamp 1649977179
transform 1 0 36892 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_74_393
timestamp 1649977179
transform 1 0 37260 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_74_396
timestamp 1649977179
transform 1 0 37536 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_74_403
timestamp 1649977179
transform 1 0 38180 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_6
timestamp 1649977179
transform 1 0 1656 0 -1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_75_12
timestamp 1649977179
transform 1 0 2208 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_24
timestamp 1649977179
transform 1 0 3312 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_36
timestamp 1649977179
transform 1 0 4416 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_40
timestamp 1649977179
transform 1 0 4784 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1649977179
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1649977179
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_57
timestamp 1649977179
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_69
timestamp 1649977179
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_81
timestamp 1649977179
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_93
timestamp 1649977179
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1649977179
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1649977179
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_113
timestamp 1649977179
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_125
timestamp 1649977179
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_137
timestamp 1649977179
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_149
timestamp 1649977179
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1649977179
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1649977179
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_169
timestamp 1649977179
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_181
timestamp 1649977179
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_193
timestamp 1649977179
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_205
timestamp 1649977179
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1649977179
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1649977179
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_225
timestamp 1649977179
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_237
timestamp 1649977179
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_249
timestamp 1649977179
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_261
timestamp 1649977179
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_276
timestamp 1649977179
transform 1 0 26496 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_281
timestamp 1649977179
transform 1 0 26956 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_291
timestamp 1649977179
transform 1 0 27876 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_303
timestamp 1649977179
transform 1 0 28980 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_315
timestamp 1649977179
transform 1 0 30084 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_327
timestamp 1649977179
transform 1 0 31188 0 -1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1649977179
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_75_337
timestamp 1649977179
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_349
timestamp 1649977179
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_361
timestamp 1649977179
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_75_373
timestamp 1649977179
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1649977179
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1649977179
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_75_395
timestamp 1649977179
transform 1 0 37444 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_75_403
timestamp 1649977179
transform 1 0 38180 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_6
timestamp 1649977179
transform 1 0 1656 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_12
timestamp 1649977179
transform 1 0 2208 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_24
timestamp 1649977179
transform 1 0 3312 0 1 43520
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_76_29
timestamp 1649977179
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_41
timestamp 1649977179
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_53
timestamp 1649977179
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_65
timestamp 1649977179
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1649977179
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1649977179
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_85
timestamp 1649977179
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_97
timestamp 1649977179
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_109
timestamp 1649977179
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_121
timestamp 1649977179
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1649977179
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1649977179
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_141
timestamp 1649977179
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_153
timestamp 1649977179
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_165
timestamp 1649977179
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_177
timestamp 1649977179
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1649977179
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1649977179
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_197
timestamp 1649977179
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_209
timestamp 1649977179
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_221
timestamp 1649977179
transform 1 0 21436 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_76_229
timestamp 1649977179
transform 1 0 22172 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_233
timestamp 1649977179
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1649977179
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1649977179
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_253
timestamp 1649977179
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_265
timestamp 1649977179
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_76_277
timestamp 1649977179
transform 1 0 26588 0 1 43520
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_76_282
timestamp 1649977179
transform 1 0 27048 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_294
timestamp 1649977179
transform 1 0 28152 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_76_306
timestamp 1649977179
transform 1 0 29256 0 1 43520
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_76_309
timestamp 1649977179
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_321
timestamp 1649977179
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_333
timestamp 1649977179
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_76_345
timestamp 1649977179
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1649977179
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1649977179
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_76_368
timestamp 1649977179
transform 1 0 34960 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_76_380
timestamp 1649977179
transform 1 0 36064 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_383
timestamp 1649977179
transform 1 0 36340 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_389
timestamp 1649977179
transform 1 0 36892 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_403
timestamp 1649977179
transform 1 0 38180 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_6
timestamp 1649977179
transform 1 0 1656 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_12
timestamp 1649977179
transform 1 0 2208 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_18
timestamp 1649977179
transform 1 0 2760 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_24
timestamp 1649977179
transform 1 0 3312 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_36
timestamp 1649977179
transform 1 0 4416 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_77_48
timestamp 1649977179
transform 1 0 5520 0 -1 44608
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_77_57
timestamp 1649977179
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_69
timestamp 1649977179
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_81
timestamp 1649977179
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_93
timestamp 1649977179
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1649977179
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1649977179
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_113
timestamp 1649977179
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_125
timestamp 1649977179
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_137
timestamp 1649977179
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_149
timestamp 1649977179
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1649977179
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1649977179
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_169
timestamp 1649977179
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_181
timestamp 1649977179
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_193
timestamp 1649977179
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_205
timestamp 1649977179
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1649977179
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1649977179
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_77_231
timestamp 1649977179
transform 1 0 22356 0 -1 44608
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_77_240
timestamp 1649977179
transform 1 0 23184 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_252
timestamp 1649977179
transform 1 0 24288 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_264
timestamp 1649977179
transform 1 0 25392 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_276
timestamp 1649977179
transform 1 0 26496 0 -1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_77_281
timestamp 1649977179
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_293
timestamp 1649977179
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_305
timestamp 1649977179
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_317
timestamp 1649977179
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1649977179
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1649977179
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_77_337
timestamp 1649977179
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_351
timestamp 1649977179
transform 1 0 33396 0 -1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_77_363
timestamp 1649977179
transform 1 0 34500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_77_375
timestamp 1649977179
transform 1 0 35604 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_378
timestamp 1649977179
transform 1 0 35880 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_384
timestamp 1649977179
transform 1 0 36432 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_77_395
timestamp 1649977179
transform 1 0 37444 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_403
timestamp 1649977179
transform 1 0 38180 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_3
timestamp 1649977179
transform 1 0 1380 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_11
timestamp 1649977179
transform 1 0 2116 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_18
timestamp 1649977179
transform 1 0 2760 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_24
timestamp 1649977179
transform 1 0 3312 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_31
timestamp 1649977179
transform 1 0 3956 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_43
timestamp 1649977179
transform 1 0 5060 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_55
timestamp 1649977179
transform 1 0 6164 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_67
timestamp 1649977179
transform 1 0 7268 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_79
timestamp 1649977179
transform 1 0 8372 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1649977179
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_85
timestamp 1649977179
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_97
timestamp 1649977179
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_109
timestamp 1649977179
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_121
timestamp 1649977179
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1649977179
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1649977179
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_141
timestamp 1649977179
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_153
timestamp 1649977179
transform 1 0 15180 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_78_161
timestamp 1649977179
transform 1 0 15916 0 1 44608
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_78_165
timestamp 1649977179
transform 1 0 16284 0 1 44608
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_78_171
timestamp 1649977179
transform 1 0 16836 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_185
timestamp 1649977179
transform 1 0 18124 0 1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_78_193
timestamp 1649977179
transform 1 0 18860 0 1 44608
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_78_197
timestamp 1649977179
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_209
timestamp 1649977179
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_221
timestamp 1649977179
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_233
timestamp 1649977179
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1649977179
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1649977179
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_253
timestamp 1649977179
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_265
timestamp 1649977179
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_277
timestamp 1649977179
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_289
timestamp 1649977179
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1649977179
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1649977179
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_78_309
timestamp 1649977179
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_321
timestamp 1649977179
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_78_333
timestamp 1649977179
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_347
timestamp 1649977179
transform 1 0 33028 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_360
timestamp 1649977179
transform 1 0 34224 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_78_365
timestamp 1649977179
transform 1 0 34684 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_78_370
timestamp 1649977179
transform 1 0 35144 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_376
timestamp 1649977179
transform 1 0 35696 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_382
timestamp 1649977179
transform 1 0 36248 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_388
timestamp 1649977179
transform 1 0 36800 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_395
timestamp 1649977179
transform 1 0 37444 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_403
timestamp 1649977179
transform 1 0 38180 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_3
timestamp 1649977179
transform 1 0 1380 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_11
timestamp 1649977179
transform 1 0 2116 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_18
timestamp 1649977179
transform 1 0 2760 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_22
timestamp 1649977179
transform 1 0 3128 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_25
timestamp 1649977179
transform 1 0 3404 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_31
timestamp 1649977179
transform 1 0 3956 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_37
timestamp 1649977179
transform 1 0 4508 0 -1 45696
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_79_43
timestamp 1649977179
transform 1 0 5060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_55
timestamp 1649977179
transform 1 0 6164 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_57
timestamp 1649977179
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_69
timestamp 1649977179
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_81
timestamp 1649977179
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_93
timestamp 1649977179
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1649977179
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1649977179
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_113
timestamp 1649977179
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_79_125
timestamp 1649977179
transform 1 0 12604 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_79_130
timestamp 1649977179
transform 1 0 13064 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_79_140
timestamp 1649977179
transform 1 0 13984 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_146
timestamp 1649977179
transform 1 0 14536 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_79_154
timestamp 1649977179
transform 1 0 15272 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_157
timestamp 1649977179
transform 1 0 15548 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_161
timestamp 1649977179
transform 1 0 15916 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_164
timestamp 1649977179
transform 1 0 16192 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_169
timestamp 1649977179
transform 1 0 16652 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_177
timestamp 1649977179
transform 1 0 17388 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_79_184
timestamp 1649977179
transform 1 0 18032 0 -1 45696
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_79_192
timestamp 1649977179
transform 1 0 18768 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_204
timestamp 1649977179
transform 1 0 19872 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_216
timestamp 1649977179
transform 1 0 20976 0 -1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_79_225
timestamp 1649977179
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_237
timestamp 1649977179
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_249
timestamp 1649977179
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_261
timestamp 1649977179
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1649977179
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1649977179
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_281
timestamp 1649977179
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_293
timestamp 1649977179
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_305
timestamp 1649977179
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_79_317
timestamp 1649977179
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1649977179
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1649977179
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_79_337
timestamp 1649977179
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_349
timestamp 1649977179
transform 1 0 33212 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_353
timestamp 1649977179
transform 1 0 33580 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_356
timestamp 1649977179
transform 1 0 33856 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_362
timestamp 1649977179
transform 1 0 34408 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_368
timestamp 1649977179
transform 1 0 34960 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_79_372
timestamp 1649977179
transform 1 0 35328 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_79_375
timestamp 1649977179
transform 1 0 35604 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_381
timestamp 1649977179
transform 1 0 36156 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_388
timestamp 1649977179
transform 1 0 36800 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_395
timestamp 1649977179
transform 1 0 37444 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_403
timestamp 1649977179
transform 1 0 38180 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_7
timestamp 1649977179
transform 1 0 1748 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_15
timestamp 1649977179
transform 1 0 2484 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_23
timestamp 1649977179
transform 1 0 3220 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1649977179
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_29
timestamp 1649977179
transform 1 0 3772 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_80_35
timestamp 1649977179
transform 1 0 4324 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_43
timestamp 1649977179
transform 1 0 5060 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_49
timestamp 1649977179
transform 1 0 5612 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_80_59
timestamp 1649977179
transform 1 0 6532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_71
timestamp 1649977179
transform 1 0 7636 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_79
timestamp 1649977179
transform 1 0 8372 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_83
timestamp 1649977179
transform 1 0 8740 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_87
timestamp 1649977179
transform 1 0 9108 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_99
timestamp 1649977179
transform 1 0 10212 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_80_111
timestamp 1649977179
transform 1 0 11316 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_115
timestamp 1649977179
transform 1 0 11684 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_119
timestamp 1649977179
transform 1 0 12052 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_122
timestamp 1649977179
transform 1 0 12328 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_128
timestamp 1649977179
transform 1 0 12880 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_135
timestamp 1649977179
transform 1 0 13524 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1649977179
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_80_141
timestamp 1649977179
transform 1 0 14076 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_80_146
timestamp 1649977179
transform 1 0 14536 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_154
timestamp 1649977179
transform 1 0 15272 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_80_164
timestamp 1649977179
transform 1 0 16192 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_80_177
timestamp 1649977179
transform 1 0 17388 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_80_188
timestamp 1649977179
transform 1 0 18400 0 1 45696
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_80_199
timestamp 1649977179
transform 1 0 19412 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_211
timestamp 1649977179
transform 1 0 20516 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_223
timestamp 1649977179
transform 1 0 21620 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_235
timestamp 1649977179
transform 1 0 22724 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_247
timestamp 1649977179
transform 1 0 23828 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1649977179
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_255
timestamp 1649977179
transform 1 0 24564 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_267
timestamp 1649977179
transform 1 0 25668 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_279
timestamp 1649977179
transform 1 0 26772 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_291
timestamp 1649977179
transform 1 0 27876 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_303
timestamp 1649977179
transform 1 0 28980 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1649977179
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_80_311
timestamp 1649977179
transform 1 0 29716 0 1 45696
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_80_323
timestamp 1649977179
transform 1 0 30820 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_335
timestamp 1649977179
transform 1 0 31924 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_341
timestamp 1649977179
transform 1 0 32476 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_347
timestamp 1649977179
transform 1 0 33028 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_353
timestamp 1649977179
transform 1 0 33580 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_357
timestamp 1649977179
transform 1 0 33948 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_360
timestamp 1649977179
transform 1 0 34224 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_365
timestamp 1649977179
transform 1 0 34684 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_369
timestamp 1649977179
transform 1 0 35052 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_80_373
timestamp 1649977179
transform 1 0 35420 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_381
timestamp 1649977179
transform 1 0 36156 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_389
timestamp 1649977179
transform 1 0 36892 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_403
timestamp 1649977179
transform 1 0 38180 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_3
timestamp 1649977179
transform 1 0 1380 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_7
timestamp 1649977179
transform 1 0 1748 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_15
timestamp 1649977179
transform 1 0 2484 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_23
timestamp 1649977179
transform 1 0 3220 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_31
timestamp 1649977179
transform 1 0 3956 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_38
timestamp 1649977179
transform 1 0 4600 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_42
timestamp 1649977179
transform 1 0 4968 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_45
timestamp 1649977179
transform 1 0 5244 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_49
timestamp 1649977179
transform 1 0 5612 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_52
timestamp 1649977179
transform 1 0 5888 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_60
timestamp 1649977179
transform 1 0 6624 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_66
timestamp 1649977179
transform 1 0 7176 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_72
timestamp 1649977179
transform 1 0 7728 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_77
timestamp 1649977179
transform 1 0 8188 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_83
timestamp 1649977179
transform 1 0 8740 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_90
timestamp 1649977179
transform 1 0 9384 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_81_100
timestamp 1649977179
transform 1 0 10304 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_81_108
timestamp 1649977179
transform 1 0 11040 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_81_113
timestamp 1649977179
transform 1 0 11500 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_118
timestamp 1649977179
transform 1 0 11960 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_126
timestamp 1649977179
transform 1 0 12696 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_129
timestamp 1649977179
transform 1 0 12972 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_142
timestamp 1649977179
transform 1 0 14168 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_155
timestamp 1649977179
transform 1 0 15364 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_163
timestamp 1649977179
transform 1 0 16100 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1649977179
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_169
timestamp 1649977179
transform 1 0 16652 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_173
timestamp 1649977179
transform 1 0 17020 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_183
timestamp 1649977179
transform 1 0 17940 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_191
timestamp 1649977179
transform 1 0 18676 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_195
timestamp 1649977179
transform 1 0 19044 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_203
timestamp 1649977179
transform 1 0 19780 0 -1 46784
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_81_206
timestamp 1649977179
transform 1 0 20056 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_81_220
timestamp 1649977179
transform 1 0 21344 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_228
timestamp 1649977179
transform 1 0 22080 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_235
timestamp 1649977179
transform 1 0 22724 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_81_241
timestamp 1649977179
transform 1 0 23276 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_247
timestamp 1649977179
transform 1 0 23828 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_250
timestamp 1649977179
transform 1 0 24104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_254
timestamp 1649977179
transform 1 0 24472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_258
timestamp 1649977179
transform 1 0 24840 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_264
timestamp 1649977179
transform 1 0 25392 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_270
timestamp 1649977179
transform 1 0 25944 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_278
timestamp 1649977179
transform 1 0 26680 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_81_281
timestamp 1649977179
transform 1 0 26956 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_289
timestamp 1649977179
transform 1 0 27692 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_293
timestamp 1649977179
transform 1 0 28060 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_300
timestamp 1649977179
transform 1 0 28704 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_306
timestamp 1649977179
transform 1 0 29256 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_310
timestamp 1649977179
transform 1 0 29624 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_314
timestamp 1649977179
transform 1 0 29992 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_320
timestamp 1649977179
transform 1 0 30544 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_326
timestamp 1649977179
transform 1 0 31096 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_332
timestamp 1649977179
transform 1 0 31648 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_337
timestamp 1649977179
transform 1 0 32108 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_345
timestamp 1649977179
transform 1 0 32844 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_81_356
timestamp 1649977179
transform 1 0 33856 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_363
timestamp 1649977179
transform 1 0 34500 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_367
timestamp 1649977179
transform 1 0 34868 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_372
timestamp 1649977179
transform 1 0 35328 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_380
timestamp 1649977179
transform 1 0 36064 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_388
timestamp 1649977179
transform 1 0 36800 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_403
timestamp 1649977179
transform 1 0 38180 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_5
timestamp 1649977179
transform 1 0 1564 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_13
timestamp 1649977179
transform 1 0 2300 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_21
timestamp 1649977179
transform 1 0 3036 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_27
timestamp 1649977179
transform 1 0 3588 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_33
timestamp 1649977179
transform 1 0 4140 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_41
timestamp 1649977179
transform 1 0 4876 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_49
timestamp 1649977179
transform 1 0 5612 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_55
timestamp 1649977179
transform 1 0 6164 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_57
timestamp 1649977179
transform 1 0 6348 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_62
timestamp 1649977179
transform 1 0 6808 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_76
timestamp 1649977179
transform 1 0 8096 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_85
timestamp 1649977179
transform 1 0 8924 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_90
timestamp 1649977179
transform 1 0 9384 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_98
timestamp 1649977179
transform 1 0 10120 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_104
timestamp 1649977179
transform 1 0 10672 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_108
timestamp 1649977179
transform 1 0 11040 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_113
timestamp 1649977179
transform 1 0 11500 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_117
timestamp 1649977179
transform 1 0 11868 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_121
timestamp 1649977179
transform 1 0 12236 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_128
timestamp 1649977179
transform 1 0 12880 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_136
timestamp 1649977179
transform 1 0 13616 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_82_141
timestamp 1649977179
transform 1 0 14076 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_153
timestamp 1649977179
transform 1 0 15180 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_159
timestamp 1649977179
transform 1 0 15732 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_164
timestamp 1649977179
transform 1 0 16192 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_179
timestamp 1649977179
transform 1 0 17572 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_82_187
timestamp 1649977179
transform 1 0 18308 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1649977179
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_82_197
timestamp 1649977179
transform 1 0 19228 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_82_202
timestamp 1649977179
transform 1 0 19688 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_209
timestamp 1649977179
transform 1 0 20332 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_217
timestamp 1649977179
transform 1 0 21068 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_223
timestamp 1649977179
transform 1 0 21620 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_225
timestamp 1649977179
transform 1 0 21804 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_229
timestamp 1649977179
transform 1 0 22172 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_234
timestamp 1649977179
transform 1 0 22632 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_248
timestamp 1649977179
transform 1 0 23920 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_263
timestamp 1649977179
transform 1 0 25300 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_82_273
timestamp 1649977179
transform 1 0 26220 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_279
timestamp 1649977179
transform 1 0 26772 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_285
timestamp 1649977179
transform 1 0 27324 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_293
timestamp 1649977179
transform 1 0 28060 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_301
timestamp 1649977179
transform 1 0 28796 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_307
timestamp 1649977179
transform 1 0 29348 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_82_312
timestamp 1649977179
transform 1 0 29808 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_322
timestamp 1649977179
transform 1 0 30728 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_330
timestamp 1649977179
transform 1 0 31464 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_341
timestamp 1649977179
transform 1 0 32476 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_345
timestamp 1649977179
transform 1 0 32844 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_356
timestamp 1649977179
transform 1 0 33856 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_365
timestamp 1649977179
transform 1 0 34684 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_82_377
timestamp 1649977179
transform 1 0 35788 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_383
timestamp 1649977179
transform 1 0 36340 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_388
timestamp 1649977179
transform 1 0 36800 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_403
timestamp 1649977179
transform 1 0 38180 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1649977179
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1649977179
transform -1 0 38824 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1649977179
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1649977179
transform -1 0 38824 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1649977179
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1649977179
transform -1 0 38824 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1649977179
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1649977179
transform -1 0 38824 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1649977179
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1649977179
transform -1 0 38824 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1649977179
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1649977179
transform -1 0 38824 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1649977179
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1649977179
transform -1 0 38824 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1649977179
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1649977179
transform -1 0 38824 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1649977179
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1649977179
transform -1 0 38824 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1649977179
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1649977179
transform -1 0 38824 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1649977179
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1649977179
transform -1 0 38824 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1649977179
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1649977179
transform -1 0 38824 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1649977179
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1649977179
transform -1 0 38824 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1649977179
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1649977179
transform -1 0 38824 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1649977179
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1649977179
transform -1 0 38824 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1649977179
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1649977179
transform -1 0 38824 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1649977179
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1649977179
transform -1 0 38824 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1649977179
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1649977179
transform -1 0 38824 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1649977179
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1649977179
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1649977179
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1649977179
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1649977179
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1649977179
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1649977179
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1649977179
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1649977179
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1649977179
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1649977179
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1649977179
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1649977179
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1649977179
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1649977179
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1649977179
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1649977179
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1649977179
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1649977179
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1649977179
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1649977179
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1649977179
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1649977179
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1649977179
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1649977179
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1649977179
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1649977179
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1649977179
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1649977179
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1649977179
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1649977179
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1649977179
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1649977179
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1649977179
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1649977179
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1649977179
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1649977179
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1649977179
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1649977179
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1649977179
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1649977179
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1649977179
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1649977179
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1649977179
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1649977179
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1649977179
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1649977179
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1649977179
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1649977179
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1649977179
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1649977179
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1649977179
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1649977179
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1649977179
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1649977179
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1649977179
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1649977179
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1649977179
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1649977179
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1649977179
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1649977179
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1649977179
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1649977179
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1649977179
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1649977179
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1649977179
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1649977179
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1649977179
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1649977179
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1649977179
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1649977179
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1649977179
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1649977179
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1649977179
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1649977179
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1649977179
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1649977179
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1649977179
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1649977179
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1649977179
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1649977179
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1649977179
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1649977179
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1649977179
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1649977179
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1649977179
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1649977179
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1649977179
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1649977179
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1649977179
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1649977179
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1649977179
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1649977179
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1649977179
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1649977179
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1649977179
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1649977179
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1649977179
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1649977179
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1649977179
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1649977179
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1649977179
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1649977179
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1649977179
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1649977179
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1649977179
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1649977179
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1649977179
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1649977179
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1649977179
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1649977179
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1649977179
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1649977179
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1649977179
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1649977179
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1649977179
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1649977179
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1649977179
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1649977179
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1649977179
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1649977179
transform 1 0 6256 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1649977179
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1649977179
transform 1 0 11408 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1649977179
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1649977179
transform 1 0 16560 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1649977179
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1649977179
transform 1 0 21712 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1649977179
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1649977179
transform 1 0 26864 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1649977179
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1649977179
transform 1 0 32016 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1649977179
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1649977179
transform 1 0 37168 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_8  _109_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 24748 0 1 29376
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_6  _110_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17756 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _111_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10212 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _112_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _113_
timestamp 1649977179
transform 1 0 23184 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _114_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 22908 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _115_
timestamp 1649977179
transform -1 0 22632 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _116_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 22264 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _117_
timestamp 1649977179
transform 1 0 21804 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _118_
timestamp 1649977179
transform -1 0 21896 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _119_
timestamp 1649977179
transform -1 0 27416 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1649977179
transform -1 0 27600 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _121_
timestamp 1649977179
transform -1 0 16192 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _122_
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _123_
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _124_
timestamp 1649977179
transform -1 0 10948 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _125_
timestamp 1649977179
transform 1 0 9016 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1649977179
transform 1 0 8372 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _127_
timestamp 1649977179
transform -1 0 27324 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1649977179
transform -1 0 27324 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _129_
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1649977179
transform -1 0 23920 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _131_
timestamp 1649977179
transform 1 0 15364 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _132_
timestamp 1649977179
transform 1 0 14536 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1649977179
transform -1 0 14536 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _134_
timestamp 1649977179
transform -1 0 2392 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1649977179
transform 1 0 2668 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _136_
timestamp 1649977179
transform 1 0 13340 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1649977179
transform 1 0 13248 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _138_
timestamp 1649977179
transform -1 0 17388 0 1 45696
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _139_
timestamp 1649977179
transform 1 0 17020 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _140_
timestamp 1649977179
transform 1 0 7544 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _141_
timestamp 1649977179
transform 1 0 6900 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _142_
timestamp 1649977179
transform -1 0 17940 0 -1 46784
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _143_
timestamp 1649977179
transform -1 0 18032 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _144_
timestamp 1649977179
transform 1 0 27876 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _145_
timestamp 1649977179
transform 1 0 27324 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _146_
timestamp 1649977179
transform 1 0 5060 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _147_
timestamp 1649977179
transform 1 0 4968 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _148_
timestamp 1649977179
transform -1 0 38180 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _149_
timestamp 1649977179
transform 1 0 37812 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _150_
timestamp 1649977179
transform 1 0 23000 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _151_
timestamp 1649977179
transform -1 0 22724 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _152_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20700 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _153_
timestamp 1649977179
transform -1 0 29440 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1649977179
transform -1 0 29808 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _155_
timestamp 1649977179
transform 1 0 21896 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _156_
timestamp 1649977179
transform 1 0 21344 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _157_
timestamp 1649977179
transform 1 0 27508 0 -1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1649977179
transform -1 0 27416 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _159_
timestamp 1649977179
transform 1 0 22448 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _160_
timestamp 1649977179
transform -1 0 22540 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _161_
timestamp 1649977179
transform -1 0 21988 0 1 41344
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1649977179
transform -1 0 22632 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _163_
timestamp 1649977179
transform -1 0 28796 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1649977179
transform -1 0 28796 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _165_
timestamp 1649977179
transform 1 0 23644 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _166_
timestamp 1649977179
transform -1 0 23276 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _167_
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _168_
timestamp 1649977179
transform -1 0 19320 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _169_
timestamp 1649977179
transform -1 0 28888 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 1649977179
transform -1 0 29532 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _171_
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _172_
timestamp 1649977179
transform 1 0 19412 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  _173_
timestamp 1649977179
transform 1 0 18124 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _174_
timestamp 1649977179
transform 1 0 21160 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _175_
timestamp 1649977179
transform -1 0 21344 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _176_
timestamp 1649977179
transform -1 0 20516 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _177_
timestamp 1649977179
transform -1 0 20332 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _178_
timestamp 1649977179
transform 1 0 20424 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _179_
timestamp 1649977179
transform 1 0 19872 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _180_
timestamp 1649977179
transform 1 0 12788 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _181_
timestamp 1649977179
transform 1 0 12512 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _182_
timestamp 1649977179
transform -1 0 23000 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _183_
timestamp 1649977179
transform -1 0 23644 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _184_
timestamp 1649977179
transform -1 0 26496 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _185_
timestamp 1649977179
transform -1 0 26772 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _186_
timestamp 1649977179
transform 1 0 13616 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1649977179
transform 1 0 13340 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _188_
timestamp 1649977179
transform 1 0 21896 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _189_
timestamp 1649977179
transform -1 0 22356 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _190_
timestamp 1649977179
transform 1 0 20792 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _191_
timestamp 1649977179
transform 1 0 20240 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _192_
timestamp 1649977179
transform -1 0 21436 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _193_
timestamp 1649977179
transform -1 0 21344 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _194_
timestamp 1649977179
transform 1 0 18032 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__mux2_1  _195_
timestamp 1649977179
transform -1 0 27784 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 1649977179
transform -1 0 27508 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _197_
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _198_
timestamp 1649977179
transform -1 0 22080 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _199_
timestamp 1649977179
transform -1 0 23276 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _200_
timestamp 1649977179
transform 1 0 23092 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _201_
timestamp 1649977179
transform 1 0 22172 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _202_
timestamp 1649977179
transform -1 0 22448 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _203_
timestamp 1649977179
transform -1 0 27600 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _204_
timestamp 1649977179
transform -1 0 27784 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _205_
timestamp 1649977179
transform -1 0 15180 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _206_
timestamp 1649977179
transform -1 0 16100 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _207_
timestamp 1649977179
transform 1 0 23920 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _208_
timestamp 1649977179
transform -1 0 23552 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _209_
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _210_
timestamp 1649977179
transform -1 0 27140 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _211_
timestamp 1649977179
transform -1 0 18032 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _212_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17572 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _213_
timestamp 1649977179
transform -1 0 25392 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _214_
timestamp 1649977179
transform -1 0 26036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _215_
timestamp 1649977179
transform 1 0 13432 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _216_
timestamp 1649977179
transform 1 0 12788 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _217_
timestamp 1649977179
transform 1 0 25484 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _218_
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _219_
timestamp 1649977179
transform 1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _220_
timestamp 1649977179
transform -1 0 4968 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _221_
timestamp 1649977179
transform 1 0 5152 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _222_
timestamp 1649977179
transform -1 0 4784 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _223_
timestamp 1649977179
transform 1 0 4876 0 -1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _224_
timestamp 1649977179
transform -1 0 4600 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _225_
timestamp 1649977179
transform 1 0 4600 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _226_
timestamp 1649977179
transform -1 0 26496 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _227_
timestamp 1649977179
transform -1 0 27140 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _228_
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _229_
timestamp 1649977179
transform 1 0 5612 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _230_
timestamp 1649977179
transform -1 0 4600 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _231_
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _232_
timestamp 1649977179
transform 1 0 27416 0 1 42432
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _233_
timestamp 1649977179
transform 1 0 26220 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _234_
timestamp 1649977179
transform 1 0 27048 0 -1 43520
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _235_
timestamp 1649977179
transform -1 0 26588 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _236_
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _237_
timestamp 1649977179
transform 1 0 3312 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _238_
timestamp 1649977179
transform 1 0 2852 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _239_
timestamp 1649977179
transform 1 0 2668 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _240_
timestamp 1649977179
transform -1 0 6900 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _241_
timestamp 1649977179
transform 1 0 7268 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _242_
timestamp 1649977179
transform -1 0 2392 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _243_
timestamp 1649977179
transform 1 0 2116 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _244_
timestamp 1649977179
transform 1 0 25208 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _245_
timestamp 1649977179
transform -1 0 33856 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _246_
timestamp 1649977179
transform 1 0 33580 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _247_
timestamp 1649977179
transform -1 0 33856 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _248_
timestamp 1649977179
transform -1 0 34500 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _249_
timestamp 1649977179
transform -1 0 15548 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _250_
timestamp 1649977179
transform 1 0 15456 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _251_
timestamp 1649977179
transform -1 0 31648 0 -1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _252_
timestamp 1649977179
transform -1 0 32384 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _253_
timestamp 1649977179
transform -1 0 34316 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _254_
timestamp 1649977179
transform -1 0 34960 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _255_
timestamp 1649977179
transform -1 0 34224 0 1 44608
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _256_
timestamp 1649977179
transform -1 0 34960 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _257_
timestamp 1649977179
transform 1 0 20332 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _258_
timestamp 1649977179
transform -1 0 20700 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _259_
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _260_
timestamp 1649977179
transform -1 0 16652 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _261_
timestamp 1649977179
transform 1 0 33764 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _262_
timestamp 1649977179
transform -1 0 34224 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _263_
timestamp 1649977179
transform 1 0 20332 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _264_
timestamp 1649977179
transform -1 0 20700 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _265_
timestamp 1649977179
transform 1 0 22264 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _266_
timestamp 1649977179
transform 1 0 22356 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _267_
timestamp 1649977179
transform 1 0 15088 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _268_
timestamp 1649977179
transform 1 0 14536 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _269_
timestamp 1649977179
transform -1 0 9568 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _270_
timestamp 1649977179
transform -1 0 12420 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _271_
timestamp 1649977179
transform -1 0 18308 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _272_
timestamp 1649977179
transform 1 0 17848 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _273_
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _274_
timestamp 1649977179
transform -1 0 34868 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _275_
timestamp 1649977179
transform 1 0 11224 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _276_
timestamp 1649977179
transform 1 0 10580 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _277_
timestamp 1649977179
transform -1 0 22172 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _278_
timestamp 1649977179
transform -1 0 22264 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_1  _279_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 22908 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _280_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21436 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _281_
timestamp 1649977179
transform -1 0 23000 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _282_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21804 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _283_
timestamp 1649977179
transform 1 0 22356 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _284_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22724 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _285_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22632 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _286_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18032 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _287_
timestamp 1649977179
transform -1 0 24932 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _288_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21344 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _289_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 23920 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _290_
timestamp 1649977179
transform -1 0 23092 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__a31o_1  _291_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22264 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _292_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21528 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _293_
timestamp 1649977179
transform -1 0 22816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _294_
timestamp 1649977179
transform 1 0 21804 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _295_
timestamp 1649977179
transform -1 0 23184 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _296_
timestamp 1649977179
transform -1 0 24932 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _297_
timestamp 1649977179
transform 1 0 24748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _298_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14996 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _299_
timestamp 1649977179
transform -1 0 16928 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _300_
timestamp 1649977179
transform -1 0 22080 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _301_
timestamp 1649977179
transform 1 0 20608 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _302_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13892 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _303_
timestamp 1649977179
transform 1 0 15364 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfstp_1  _304_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14168 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _304__260 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 14812 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _305_
timestamp 1649977179
transform 1 0 15364 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  _306__259
timestamp 1649977179
transform -1 0 19872 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_1  _306_
timestamp 1649977179
transform 1 0 19320 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__dfstp_1  _307_
timestamp 1649977179
transform 1 0 20240 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_i_clk opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14720 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_i_clk
timestamp 1649977179
transform 1 0 12972 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_i_clk
timestamp 1649977179
transform 1 0 12972 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15456 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1649977179
transform -1 0 17388 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1
timestamp 1649977179
transform -1 0 2300 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1649977179
transform 1 0 9016 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform 1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1649977179
transform 1 0 35144 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 37168 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform -1 0 1656 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1649977179
transform -1 0 1656 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1649977179
transform -1 0 6808 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1649977179
transform -1 0 1656 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform -1 0 21344 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1649977179
transform -1 0 38180 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform 1 0 35052 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 4600 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1649977179
transform -1 0 2300 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform -1 0 2944 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform -1 0 1656 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1649977179
transform -1 0 38180 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform -1 0 11040 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1649977179
transform 1 0 37260 0 -1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1649977179
transform 1 0 1932 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform 1 0 37904 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1649977179
transform 1 0 14260 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1649977179
transform -1 0 38180 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1649977179
transform -1 0 11776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1649977179
transform -1 0 2300 0 -1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1649977179
transform 1 0 37904 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1649977179
transform -1 0 2300 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1649977179
transform -1 0 38180 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1649977179
transform -1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input32
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input33
timestamp 1649977179
transform -1 0 2300 0 -1 41344
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform 1 0 37904 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input35
timestamp 1649977179
transform -1 0 2300 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform -1 0 1656 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform 1 0 37904 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform 1 0 37904 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1649977179
transform 1 0 33580 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform -1 0 1656 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform 1 0 37904 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1649977179
transform -1 0 38180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform -1 0 19044 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input44
timestamp 1649977179
transform 1 0 37260 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1649977179
transform 1 0 29716 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1649977179
transform 1 0 37904 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1649977179
transform 1 0 19412 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1649977179
transform -1 0 6624 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1649977179
transform -1 0 12880 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1649977179
transform 1 0 28428 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input51
timestamp 1649977179
transform 1 0 23000 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1649977179
transform 1 0 37904 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1649977179
transform 1 0 37904 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1649977179
transform -1 0 1656 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1649977179
transform -1 0 7452 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1649977179
transform -1 0 1656 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input57
timestamp 1649977179
transform -1 0 38180 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input58
timestamp 1649977179
transform -1 0 2300 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1649977179
transform 1 0 4508 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1649977179
transform -1 0 1656 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1649977179
transform 1 0 20056 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input62
timestamp 1649977179
transform 1 0 16652 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1649977179
transform 1 0 2116 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1649977179
transform 1 0 2116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input65
timestamp 1649977179
transform 1 0 37260 0 1 45696
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1649977179
transform -1 0 16008 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input67
timestamp 1649977179
transform 1 0 32936 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1649977179
transform -1 0 22080 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input69
timestamp 1649977179
transform -1 0 2300 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1649977179
transform -1 0 1656 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1649977179
transform -1 0 15548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1649977179
transform -1 0 1656 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1649977179
transform 1 0 18124 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1649977179
transform -1 0 34500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1649977179
transform 1 0 1748 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input76
timestamp 1649977179
transform 1 0 1748 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input77
timestamp 1649977179
transform 1 0 1380 0 -1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1649977179
transform -1 0 13248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input79
timestamp 1649977179
transform 1 0 37904 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input80
timestamp 1649977179
transform 1 0 36524 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input81
timestamp 1649977179
transform 1 0 2852 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input82
timestamp 1649977179
transform 1 0 23276 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input83
timestamp 1649977179
transform -1 0 2300 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1649977179
transform -1 0 1656 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1649977179
transform -1 0 2300 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input86
timestamp 1649977179
transform 1 0 13248 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input87
timestamp 1649977179
transform -1 0 38180 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1649977179
transform 1 0 35696 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1649977179
transform 1 0 37904 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1649977179
transform 1 0 31004 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input91
timestamp 1649977179
transform 1 0 1748 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1649977179
transform -1 0 9384 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input93
timestamp 1649977179
transform 1 0 37904 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input94
timestamp 1649977179
transform 1 0 18768 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input95
timestamp 1649977179
transform 1 0 37168 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input96
timestamp 1649977179
transform -1 0 1656 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 1649977179
transform 1 0 32752 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input98
timestamp 1649977179
transform 1 0 1748 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input99
timestamp 1649977179
transform 1 0 7176 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input100
timestamp 1649977179
transform 1 0 37904 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input101
timestamp 1649977179
transform -1 0 1656 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input102
timestamp 1649977179
transform 1 0 34868 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input103
timestamp 1649977179
transform -1 0 36064 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input104
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input105
timestamp 1649977179
transform 1 0 3956 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input106
timestamp 1649977179
transform 1 0 28428 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input107
timestamp 1649977179
transform 1 0 37904 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input108
timestamp 1649977179
transform -1 0 38180 0 1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input109
timestamp 1649977179
transform 1 0 29716 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input110
timestamp 1649977179
transform -1 0 36064 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input111
timestamp 1649977179
transform -1 0 2300 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input112
timestamp 1649977179
transform 1 0 11684 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input113
timestamp 1649977179
transform 1 0 1748 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input114
timestamp 1649977179
transform -1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input115
timestamp 1649977179
transform -1 0 38180 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input116
timestamp 1649977179
transform 1 0 24380 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input117
timestamp 1649977179
transform 1 0 37904 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input118
timestamp 1649977179
transform 1 0 2668 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input119
timestamp 1649977179
transform 1 0 5244 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input120
timestamp 1649977179
transform 1 0 3772 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input121
timestamp 1649977179
transform 1 0 2852 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input122
timestamp 1649977179
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input123
timestamp 1649977179
transform 1 0 37904 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input124
timestamp 1649977179
transform 1 0 21988 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input125
timestamp 1649977179
transform 1 0 37260 0 1 46784
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input126
timestamp 1649977179
transform 1 0 37260 0 1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input127
timestamp 1649977179
transform -1 0 11960 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input128
timestamp 1649977179
transform 1 0 5520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input129
timestamp 1649977179
transform 1 0 37904 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input130
timestamp 1649977179
transform -1 0 38180 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input131
timestamp 1649977179
transform 1 0 1748 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input132
timestamp 1649977179
transform 1 0 37904 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input133
timestamp 1649977179
transform 1 0 27600 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input134
timestamp 1649977179
transform -1 0 1656 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input135
timestamp 1649977179
transform 1 0 37904 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input136
timestamp 1649977179
transform 1 0 34224 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input137
timestamp 1649977179
transform -1 0 38180 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input138
timestamp 1649977179
transform -1 0 32844 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input139
timestamp 1649977179
transform -1 0 1656 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input140
timestamp 1649977179
transform -1 0 1656 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input141
timestamp 1649977179
transform 1 0 28244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input142
timestamp 1649977179
transform -1 0 3864 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input143
timestamp 1649977179
transform 1 0 33396 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input144
timestamp 1649977179
transform -1 0 1656 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input145
timestamp 1649977179
transform -1 0 2760 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input146
timestamp 1649977179
transform -1 0 1656 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input147
timestamp 1649977179
transform -1 0 2300 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input148
timestamp 1649977179
transform 1 0 8464 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input149
timestamp 1649977179
transform -1 0 4048 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input150
timestamp 1649977179
transform 1 0 22448 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input151
timestamp 1649977179
transform -1 0 12236 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input152
timestamp 1649977179
transform -1 0 23644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input153
timestamp 1649977179
transform 1 0 29532 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input154
timestamp 1649977179
transform 1 0 37904 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input155
timestamp 1649977179
transform -1 0 1656 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input156
timestamp 1649977179
transform 1 0 37904 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input157
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input158
timestamp 1649977179
transform 1 0 15916 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input159
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input160
timestamp 1649977179
transform -1 0 38180 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input161
timestamp 1649977179
transform 1 0 27600 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input162
timestamp 1649977179
transform -1 0 26220 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input163
timestamp 1649977179
transform 1 0 24564 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input164
timestamp 1649977179
transform -1 0 1656 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input165
timestamp 1649977179
transform -1 0 2760 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input166
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input167
timestamp 1649977179
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input168
timestamp 1649977179
transform -1 0 2300 0 1 38080
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input169
timestamp 1649977179
transform 1 0 37904 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output170
timestamp 1649977179
transform -1 0 2484 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output171
timestamp 1649977179
transform 1 0 37076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output172
timestamp 1649977179
transform -1 0 5612 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output173
timestamp 1649977179
transform -1 0 1748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output174
timestamp 1649977179
transform -1 0 10028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output175
timestamp 1649977179
transform 1 0 37812 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output176
timestamp 1649977179
transform -1 0 16100 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output177
timestamp 1649977179
transform -1 0 1748 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output178
timestamp 1649977179
transform 1 0 37812 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output179
timestamp 1649977179
transform -1 0 33948 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output180
timestamp 1649977179
transform -1 0 1748 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output181
timestamp 1649977179
transform -1 0 3220 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output182
timestamp 1649977179
transform -1 0 8188 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output183
timestamp 1649977179
transform 1 0 37812 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output184
timestamp 1649977179
transform 1 0 28428 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output185
timestamp 1649977179
transform 1 0 37812 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output186
timestamp 1649977179
transform 1 0 37812 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output187
timestamp 1649977179
transform 1 0 37812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output188
timestamp 1649977179
transform -1 0 10764 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1649977179
transform 1 0 27692 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output190
timestamp 1649977179
transform -1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1649977179
transform 1 0 26956 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output192
timestamp 1649977179
transform 1 0 31004 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1649977179
transform -1 0 1748 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1649977179
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1649977179
transform 1 0 37812 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1649977179
transform -1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1649977179
transform -1 0 1748 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1649977179
transform -1 0 17204 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1649977179
transform -1 0 1748 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output200
timestamp 1649977179
transform 1 0 17940 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1649977179
transform -1 0 1748 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1649977179
transform -1 0 1748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output203
timestamp 1649977179
transform 1 0 37812 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1649977179
transform 1 0 30360 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output205
timestamp 1649977179
transform 1 0 37444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1649977179
transform -1 0 10120 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1649977179
transform -1 0 3956 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output208
timestamp 1649977179
transform 1 0 35696 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1649977179
transform 1 0 25576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1649977179
transform 1 0 14904 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output211
timestamp 1649977179
transform -1 0 1748 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1649977179
transform -1 0 1748 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1649977179
transform 1 0 31096 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output214
timestamp 1649977179
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1649977179
transform 1 0 37812 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 1649977179
transform -1 0 1748 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output217
timestamp 1649977179
transform 1 0 32108 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1649977179
transform 1 0 36524 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output219
timestamp 1649977179
transform 1 0 24564 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1649977179
transform 1 0 37812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1649977179
transform 1 0 37812 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1649977179
transform 1 0 36432 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1649977179
transform 1 0 22264 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 1649977179
transform -1 0 1748 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output226
timestamp 1649977179
transform 1 0 37812 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1649977179
transform 1 0 37812 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 1649977179
transform -1 0 1748 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output229
timestamp 1649977179
transform 1 0 37812 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1649977179
transform 1 0 37812 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 1649977179
transform 1 0 34868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 1649977179
transform 1 0 35788 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 1649977179
transform 1 0 37812 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output234
timestamp 1649977179
transform 1 0 20700 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output235
timestamp 1649977179
transform -1 0 4876 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output236
timestamp 1649977179
transform 1 0 37812 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output237
timestamp 1649977179
transform 1 0 20700 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output238
timestamp 1649977179
transform -1 0 1748 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output239
timestamp 1649977179
transform -1 0 1748 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output240
timestamp 1649977179
transform -1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output241
timestamp 1649977179
transform 1 0 37812 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output242
timestamp 1649977179
transform 1 0 37812 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output243
timestamp 1649977179
transform 1 0 34960 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output244
timestamp 1649977179
transform -1 0 16192 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output245
timestamp 1649977179
transform -1 0 13340 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output246
timestamp 1649977179
transform -1 0 1748 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output247
timestamp 1649977179
transform -1 0 1748 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output248
timestamp 1649977179
transform 1 0 37812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output249
timestamp 1649977179
transform -1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output250
timestamp 1649977179
transform 1 0 36340 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output251
timestamp 1649977179
transform -1 0 6900 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output252
timestamp 1649977179
transform -1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output253
timestamp 1649977179
transform 1 0 37812 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output254
timestamp 1649977179
transform 1 0 36432 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output255
timestamp 1649977179
transform 1 0 37812 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output256
timestamp 1649977179
transform 1 0 37812 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output257
timestamp 1649977179
transform -1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output258
timestamp 1649977179
transform 1 0 37812 0 1 26112
box -38 -48 406 592
<< labels >>
flabel metal3 s 0 47608 800 47728 0 FreeSans 480 0 0 0 c_wb_4_burst
port 0 nsew signal tristate
flabel metal2 s 38658 0 38714 800 0 FreeSans 224 90 0 0 c_wb_8_burst
port 1 nsew signal tristate
flabel metal3 s 0 34008 800 34128 0 FreeSans 480 0 0 0 c_wb_ack_cmp
port 2 nsew signal input
flabel metal2 s 5170 0 5226 800 0 FreeSans 224 90 0 0 c_wb_adr[0]
port 3 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 c_wb_adr[10]
port 4 nsew signal tristate
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 c_wb_adr[11]
port 5 nsew signal tristate
flabel metal3 s 39200 27208 40000 27328 0 FreeSans 480 0 0 0 c_wb_adr[12]
port 6 nsew signal tristate
flabel metal2 s 15474 49200 15530 50000 0 FreeSans 224 90 0 0 c_wb_adr[13]
port 7 nsew signal tristate
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 c_wb_adr[14]
port 8 nsew signal tristate
flabel metal3 s 39200 15648 40000 15768 0 FreeSans 480 0 0 0 c_wb_adr[15]
port 9 nsew signal tristate
flabel metal2 s 33506 0 33562 800 0 FreeSans 224 90 0 0 c_wb_adr[16]
port 10 nsew signal tristate
flabel metal3 s 0 36728 800 36848 0 FreeSans 480 0 0 0 c_wb_adr[17]
port 11 nsew signal tristate
flabel metal3 s 0 49648 800 49768 0 FreeSans 480 0 0 0 c_wb_adr[18]
port 12 nsew signal tristate
flabel metal2 s 7746 49200 7802 50000 0 FreeSans 224 90 0 0 c_wb_adr[19]
port 13 nsew signal tristate
flabel metal3 s 39200 36048 40000 36168 0 FreeSans 480 0 0 0 c_wb_adr[1]
port 14 nsew signal tristate
flabel metal2 s 27710 49200 27766 50000 0 FreeSans 224 90 0 0 c_wb_adr[20]
port 15 nsew signal tristate
flabel metal3 s 39200 29928 40000 30048 0 FreeSans 480 0 0 0 c_wb_adr[21]
port 16 nsew signal tristate
flabel metal3 s 39200 27888 40000 28008 0 FreeSans 480 0 0 0 c_wb_adr[22]
port 17 nsew signal tristate
flabel metal3 s 39200 6128 40000 6248 0 FreeSans 480 0 0 0 c_wb_adr[23]
port 18 nsew signal tristate
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 c_wb_adr[2]
port 19 nsew signal tristate
flabel metal2 s 27066 49200 27122 50000 0 FreeSans 224 90 0 0 c_wb_adr[3]
port 20 nsew signal tristate
flabel metal3 s 0 6128 800 6248 0 FreeSans 480 0 0 0 c_wb_adr[4]
port 21 nsew signal tristate
flabel metal2 s 26422 49200 26478 50000 0 FreeSans 224 90 0 0 c_wb_adr[5]
port 22 nsew signal tristate
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 c_wb_adr[6]
port 23 nsew signal tristate
flabel metal3 s 0 34688 800 34808 0 FreeSans 480 0 0 0 c_wb_adr[7]
port 24 nsew signal tristate
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 c_wb_adr[8]
port 25 nsew signal tristate
flabel metal3 s 39200 23808 40000 23928 0 FreeSans 480 0 0 0 c_wb_adr[9]
port 26 nsew signal tristate
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 c_wb_cyc
port 27 nsew signal tristate
flabel metal2 s 8390 49200 8446 50000 0 FreeSans 224 90 0 0 c_wb_err_cmp
port 28 nsew signal input
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 c_wb_i_dat_cmp[0]
port 29 nsew signal input
flabel metal2 s 35438 49200 35494 50000 0 FreeSans 224 90 0 0 c_wb_i_dat_cmp[10]
port 30 nsew signal input
flabel metal3 s 39200 45568 40000 45688 0 FreeSans 480 0 0 0 c_wb_i_dat_cmp[11]
port 31 nsew signal input
flabel metal3 s 0 17008 800 17128 0 FreeSans 480 0 0 0 c_wb_i_dat_cmp[12]
port 32 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 c_wb_i_dat_cmp[13]
port 33 nsew signal input
flabel metal2 s 6458 49200 6514 50000 0 FreeSans 224 90 0 0 c_wb_i_dat_cmp[14]
port 34 nsew signal input
flabel metal3 s 0 44208 800 44328 0 FreeSans 480 0 0 0 c_wb_i_dat_cmp[15]
port 35 nsew signal input
flabel metal2 s 21270 0 21326 800 0 FreeSans 224 90 0 0 c_wb_i_dat_cmp[1]
port 36 nsew signal input
flabel metal3 s 39200 31288 40000 31408 0 FreeSans 480 0 0 0 c_wb_i_dat_cmp[2]
port 37 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 c_wb_i_dat_cmp[3]
port 38 nsew signal input
flabel metal2 s 3882 49200 3938 50000 0 FreeSans 224 90 0 0 c_wb_i_dat_cmp[4]
port 39 nsew signal input
flabel metal3 s 0 8168 800 8288 0 FreeSans 480 0 0 0 c_wb_i_dat_cmp[5]
port 40 nsew signal input
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 c_wb_i_dat_cmp[6]
port 41 nsew signal input
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 c_wb_i_dat_cmp[7]
port 42 nsew signal input
flabel metal3 s 0 31288 800 31408 0 FreeSans 480 0 0 0 c_wb_i_dat_cmp[8]
port 43 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 c_wb_i_dat_cmp[9]
port 44 nsew signal input
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 c_wb_o_dat[0]
port 45 nsew signal tristate
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 c_wb_o_dat[10]
port 46 nsew signal tristate
flabel metal3 s 0 35368 800 35488 0 FreeSans 480 0 0 0 c_wb_o_dat[11]
port 47 nsew signal tristate
flabel metal2 s 17406 49200 17462 50000 0 FreeSans 224 90 0 0 c_wb_o_dat[12]
port 48 nsew signal tristate
flabel metal3 s 0 5448 800 5568 0 FreeSans 480 0 0 0 c_wb_o_dat[13]
port 49 nsew signal tristate
flabel metal3 s 0 29248 800 29368 0 FreeSans 480 0 0 0 c_wb_o_dat[14]
port 50 nsew signal tristate
flabel metal3 s 39200 4768 40000 4888 0 FreeSans 480 0 0 0 c_wb_o_dat[15]
port 51 nsew signal tristate
flabel metal2 s 30286 49200 30342 50000 0 FreeSans 224 90 0 0 c_wb_o_dat[1]
port 52 nsew signal tristate
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 c_wb_o_dat[2]
port 53 nsew signal tristate
flabel metal2 s 9678 49200 9734 50000 0 FreeSans 224 90 0 0 c_wb_o_dat[3]
port 54 nsew signal tristate
flabel metal2 s 662 49200 718 50000 0 FreeSans 224 90 0 0 c_wb_o_dat[4]
port 55 nsew signal tristate
flabel metal3 s 39200 1368 40000 1488 0 FreeSans 480 0 0 0 c_wb_o_dat[5]
port 56 nsew signal tristate
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 c_wb_o_dat[6]
port 57 nsew signal tristate
flabel metal2 s 14830 49200 14886 50000 0 FreeSans 224 90 0 0 c_wb_o_dat[7]
port 58 nsew signal tristate
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 c_wb_o_dat[8]
port 59 nsew signal tristate
flabel metal3 s 0 45568 800 45688 0 FreeSans 480 0 0 0 c_wb_o_dat[9]
port 60 nsew signal tristate
flabel metal2 s 30930 49200 30986 50000 0 FreeSans 224 90 0 0 c_wb_sel[0]
port 61 nsew signal tristate
flabel metal2 s 18050 0 18106 800 0 FreeSans 224 90 0 0 c_wb_sel[1]
port 62 nsew signal tristate
flabel metal3 s 39200 38768 40000 38888 0 FreeSans 480 0 0 0 c_wb_stb
port 63 nsew signal tristate
flabel metal3 s 0 38768 800 38888 0 FreeSans 480 0 0 0 c_wb_we
port 64 nsew signal tristate
flabel metal3 s 39200 22448 40000 22568 0 FreeSans 480 0 0 0 cc_wb_4_burst
port 65 nsew signal input
flabel metal2 s 10966 49200 11022 50000 0 FreeSans 224 90 0 0 cc_wb_8_burst
port 66 nsew signal input
flabel metal2 s 38014 49200 38070 50000 0 FreeSans 224 90 0 0 cc_wb_adr[0]
port 67 nsew signal input
flabel metal2 s 1950 49200 2006 50000 0 FreeSans 224 90 0 0 cc_wb_adr[10]
port 68 nsew signal input
flabel metal3 s 39200 28568 40000 28688 0 FreeSans 480 0 0 0 cc_wb_adr[11]
port 69 nsew signal input
flabel metal2 s 14186 49200 14242 50000 0 FreeSans 224 90 0 0 cc_wb_adr[12]
port 70 nsew signal input
flabel metal3 s 39200 12248 40000 12368 0 FreeSans 480 0 0 0 cc_wb_adr[13]
port 71 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 cc_wb_adr[14]
port 72 nsew signal input
flabel metal3 s 0 37408 800 37528 0 FreeSans 480 0 0 0 cc_wb_adr[15]
port 73 nsew signal input
flabel metal3 s 39200 17688 40000 17808 0 FreeSans 480 0 0 0 cc_wb_adr[16]
port 74 nsew signal input
flabel metal3 s 0 3408 800 3528 0 FreeSans 480 0 0 0 cc_wb_adr[17]
port 75 nsew signal input
flabel metal3 s 39200 4088 40000 4208 0 FreeSans 480 0 0 0 cc_wb_adr[18]
port 76 nsew signal input
flabel metal2 s 36726 0 36782 800 0 FreeSans 224 90 0 0 cc_wb_adr[19]
port 77 nsew signal input
flabel metal3 s 39200 11568 40000 11688 0 FreeSans 480 0 0 0 cc_wb_adr[1]
port 78 nsew signal input
flabel metal3 s 0 40808 800 40928 0 FreeSans 480 0 0 0 cc_wb_adr[20]
port 79 nsew signal input
flabel metal3 s 39200 25168 40000 25288 0 FreeSans 480 0 0 0 cc_wb_adr[21]
port 80 nsew signal input
flabel metal3 s 0 7488 800 7608 0 FreeSans 480 0 0 0 cc_wb_adr[22]
port 81 nsew signal input
flabel metal3 s 0 24488 800 24608 0 FreeSans 480 0 0 0 cc_wb_adr[23]
port 82 nsew signal input
flabel metal3 s 39200 10208 40000 10328 0 FreeSans 480 0 0 0 cc_wb_adr[2]
port 83 nsew signal input
flabel metal3 s 39200 40808 40000 40928 0 FreeSans 480 0 0 0 cc_wb_adr[3]
port 84 nsew signal input
flabel metal2 s 33506 49200 33562 50000 0 FreeSans 224 90 0 0 cc_wb_adr[4]
port 85 nsew signal input
flabel metal3 s 0 42848 800 42968 0 FreeSans 480 0 0 0 cc_wb_adr[5]
port 86 nsew signal input
flabel metal3 s 39200 32648 40000 32768 0 FreeSans 480 0 0 0 cc_wb_adr[6]
port 87 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 cc_wb_adr[7]
port 88 nsew signal input
flabel metal2 s 18694 49200 18750 50000 0 FreeSans 224 90 0 0 cc_wb_adr[8]
port 89 nsew signal input
flabel metal3 s 39200 8 40000 128 0 FreeSans 480 0 0 0 cc_wb_adr[9]
port 90 nsew signal input
flabel metal2 s 29642 49200 29698 50000 0 FreeSans 224 90 0 0 cc_wb_cyc
port 91 nsew signal input
flabel metal3 s 39200 40128 40000 40248 0 FreeSans 480 0 0 0 cc_wb_o_dat[0]
port 92 nsew signal input
flabel metal2 s 19338 49200 19394 50000 0 FreeSans 224 90 0 0 cc_wb_o_dat[10]
port 93 nsew signal input
flabel metal2 s 5814 49200 5870 50000 0 FreeSans 224 90 0 0 cc_wb_o_dat[11]
port 94 nsew signal input
flabel metal2 s 12898 49200 12954 50000 0 FreeSans 224 90 0 0 cc_wb_o_dat[12]
port 95 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 cc_wb_o_dat[13]
port 96 nsew signal input
flabel metal2 s 23202 49200 23258 50000 0 FreeSans 224 90 0 0 cc_wb_o_dat[14]
port 97 nsew signal input
flabel metal3 s 39200 17008 40000 17128 0 FreeSans 480 0 0 0 cc_wb_o_dat[15]
port 98 nsew signal input
flabel metal3 s 39200 34008 40000 34128 0 FreeSans 480 0 0 0 cc_wb_o_dat[1]
port 99 nsew signal input
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 cc_wb_o_dat[2]
port 100 nsew signal input
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 cc_wb_o_dat[3]
port 101 nsew signal input
flabel metal3 s 0 42168 800 42288 0 FreeSans 480 0 0 0 cc_wb_o_dat[4]
port 102 nsew signal input
flabel metal3 s 39200 46928 40000 47048 0 FreeSans 480 0 0 0 cc_wb_o_dat[5]
port 103 nsew signal input
flabel metal3 s 0 688 800 808 0 FreeSans 480 0 0 0 cc_wb_o_dat[6]
port 104 nsew signal input
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 cc_wb_o_dat[7]
port 105 nsew signal input
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 cc_wb_o_dat[8]
port 106 nsew signal input
flabel metal2 s 19982 49200 20038 50000 0 FreeSans 224 90 0 0 cc_wb_o_dat[9]
port 107 nsew signal input
flabel metal2 s 16118 49200 16174 50000 0 FreeSans 224 90 0 0 cc_wb_sel[0]
port 108 nsew signal input
flabel metal3 s 0 48288 800 48408 0 FreeSans 480 0 0 0 cc_wb_sel[1]
port 109 nsew signal input
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 cc_wb_stb
port 110 nsew signal input
flabel metal2 s 39302 49200 39358 50000 0 FreeSans 224 90 0 0 cc_wb_we
port 111 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 cw_ack
port 112 nsew signal input
flabel metal2 s 32862 49200 32918 50000 0 FreeSans 224 90 0 0 cw_clk
port 113 nsew signal input
flabel metal2 s 21270 49200 21326 50000 0 FreeSans 224 90 0 0 cw_err
port 114 nsew signal input
flabel metal3 s 0 19728 800 19848 0 FreeSans 480 0 0 0 cw_io_i[0]
port 115 nsew signal input
flabel metal3 s 0 32648 800 32768 0 FreeSans 480 0 0 0 cw_io_i[10]
port 116 nsew signal input
flabel metal2 s 15474 0 15530 800 0 FreeSans 224 90 0 0 cw_io_i[11]
port 117 nsew signal input
flabel metal3 s 0 4768 800 4888 0 FreeSans 480 0 0 0 cw_io_i[12]
port 118 nsew signal input
flabel metal2 s 18050 49200 18106 50000 0 FreeSans 224 90 0 0 cw_io_i[13]
port 119 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 cw_io_i[14]
port 120 nsew signal input
flabel metal3 s 0 40128 800 40248 0 FreeSans 480 0 0 0 cw_io_i[15]
port 121 nsew signal input
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 cw_io_i[1]
port 122 nsew signal input
flabel metal3 s 0 39448 800 39568 0 FreeSans 480 0 0 0 cw_io_i[2]
port 123 nsew signal input
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 cw_io_i[3]
port 124 nsew signal input
flabel metal3 s 39200 29248 40000 29368 0 FreeSans 480 0 0 0 cw_io_i[4]
port 125 nsew signal input
flabel metal2 s 38658 49200 38714 50000 0 FreeSans 224 90 0 0 cw_io_i[5]
port 126 nsew signal input
flabel metal3 s 0 48968 800 49088 0 FreeSans 480 0 0 0 cw_io_i[6]
port 127 nsew signal input
flabel metal2 s 23202 0 23258 800 0 FreeSans 224 90 0 0 cw_io_i[7]
port 128 nsew signal input
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 cw_io_i[8]
port 129 nsew signal input
flabel metal3 s 0 28568 800 28688 0 FreeSans 480 0 0 0 cw_io_i[9]
port 130 nsew signal input
flabel metal2 s 31574 49200 31630 50000 0 FreeSans 224 90 0 0 cw_rst
port 131 nsew signal tristate
flabel metal3 s 39200 48288 40000 48408 0 FreeSans 480 0 0 0 cw_rst_z
port 132 nsew signal tristate
flabel metal3 s 0 2728 800 2848 0 FreeSans 480 0 0 0 i_clk
port 133 nsew signal input
flabel metal3 s 0 1368 800 1488 0 FreeSans 480 0 0 0 i_irq
port 134 nsew signal input
flabel metal2 s 13542 49200 13598 50000 0 FreeSans 224 90 0 0 i_rst
port 135 nsew signal input
flabel metal3 s 39200 9528 40000 9648 0 FreeSans 480 0 0 0 ic_split_clock
port 136 nsew signal input
flabel metal2 s 24490 0 24546 800 0 FreeSans 224 90 0 0 irq_s
port 137 nsew signal tristate
flabel metal3 s 39200 30608 40000 30728 0 FreeSans 480 0 0 0 la_cw_ack
port 138 nsew signal input
flabel metal2 s 36082 0 36138 800 0 FreeSans 224 90 0 0 la_cw_io_i[0]
port 139 nsew signal input
flabel metal3 s 39200 42168 40000 42288 0 FreeSans 480 0 0 0 la_cw_io_i[10]
port 140 nsew signal input
flabel metal2 s 30930 0 30986 800 0 FreeSans 224 90 0 0 la_cw_io_i[11]
port 141 nsew signal input
flabel metal2 s 18 49200 74 50000 0 FreeSans 224 90 0 0 la_cw_io_i[12]
port 142 nsew signal input
flabel metal2 s 9034 49200 9090 50000 0 FreeSans 224 90 0 0 la_cw_io_i[13]
port 143 nsew signal input
flabel metal3 s 39200 10888 40000 11008 0 FreeSans 480 0 0 0 la_cw_io_i[14]
port 144 nsew signal input
flabel metal2 s 18694 0 18750 800 0 FreeSans 224 90 0 0 la_cw_io_i[15]
port 145 nsew signal input
flabel metal3 s 39200 16328 40000 16448 0 FreeSans 480 0 0 0 la_cw_io_i[1]
port 146 nsew signal input
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 la_cw_io_i[2]
port 147 nsew signal input
flabel metal2 s 32218 0 32274 800 0 FreeSans 224 90 0 0 la_cw_io_i[3]
port 148 nsew signal input
flabel metal3 s 0 23808 800 23928 0 FreeSans 480 0 0 0 la_cw_io_i[4]
port 149 nsew signal input
flabel metal2 s 7102 49200 7158 50000 0 FreeSans 224 90 0 0 la_cw_io_i[5]
port 150 nsew signal input
flabel metal3 s 39200 21768 40000 21888 0 FreeSans 480 0 0 0 la_cw_io_i[6]
port 151 nsew signal input
flabel metal3 s 0 22448 800 22568 0 FreeSans 480 0 0 0 la_cw_io_i[7]
port 152 nsew signal input
flabel metal2 s 34794 49200 34850 50000 0 FreeSans 224 90 0 0 la_cw_io_i[8]
port 153 nsew signal input
flabel metal3 s 39200 688 40000 808 0 FreeSans 480 0 0 0 la_cw_io_i[9]
port 154 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 la_cw_ovr
port 155 nsew signal input
flabel metal3 s 39200 7488 40000 7608 0 FreeSans 480 0 0 0 m_cw_ack
port 156 nsew signal tristate
flabel metal3 s 39200 44208 40000 44328 0 FreeSans 480 0 0 0 m_cw_err
port 157 nsew signal tristate
flabel metal2 s 37370 49200 37426 50000 0 FreeSans 224 90 0 0 m_cw_io_i[0]
port 158 nsew signal tristate
flabel metal2 s 22558 49200 22614 50000 0 FreeSans 224 90 0 0 m_cw_io_i[10]
port 159 nsew signal tristate
flabel metal3 s 0 26528 800 26648 0 FreeSans 480 0 0 0 m_cw_io_i[11]
port 160 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 m_cw_io_i[12]
port 161 nsew signal tristate
flabel metal3 s 39200 23128 40000 23248 0 FreeSans 480 0 0 0 m_cw_io_i[13]
port 162 nsew signal tristate
flabel metal3 s 39200 21088 40000 21208 0 FreeSans 480 0 0 0 m_cw_io_i[14]
port 163 nsew signal tristate
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 m_cw_io_i[15]
port 164 nsew signal tristate
flabel metal3 s 39200 18368 40000 18488 0 FreeSans 480 0 0 0 m_cw_io_i[1]
port 165 nsew signal tristate
flabel metal3 s 39200 8168 40000 8288 0 FreeSans 480 0 0 0 m_cw_io_i[2]
port 166 nsew signal tristate
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 m_cw_io_i[3]
port 167 nsew signal tristate
flabel metal3 s 39200 47608 40000 47728 0 FreeSans 480 0 0 0 m_cw_io_i[4]
port 168 nsew signal tristate
flabel metal3 s 39200 37408 40000 37528 0 FreeSans 480 0 0 0 m_cw_io_i[5]
port 169 nsew signal tristate
flabel metal2 s 20626 0 20682 800 0 FreeSans 224 90 0 0 m_cw_io_i[6]
port 170 nsew signal tristate
flabel metal2 s 4526 49200 4582 50000 0 FreeSans 224 90 0 0 m_cw_io_i[7]
port 171 nsew signal tristate
flabel metal3 s 39200 5448 40000 5568 0 FreeSans 480 0 0 0 m_cw_io_i[8]
port 172 nsew signal tristate
flabel metal2 s 20626 49200 20682 50000 0 FreeSans 224 90 0 0 m_cw_io_i[9]
port 173 nsew signal tristate
flabel metal3 s 0 29928 800 30048 0 FreeSans 480 0 0 0 s_rst
port 174 nsew signal tristate
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 u_wb_4_burst
port 175 nsew signal input
flabel metal2 s 28354 49200 28410 50000 0 FreeSans 224 90 0 0 u_wb_8_burst
port 176 nsew signal input
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 u_wb_ack
port 177 nsew signal tristate
flabel metal3 s 39200 35368 40000 35488 0 FreeSans 480 0 0 0 u_wb_ack_cc
port 178 nsew signal input
flabel metal2 s 13542 0 13598 800 0 FreeSans 224 90 0 0 u_wb_ack_clk
port 179 nsew signal tristate
flabel metal3 s 39200 44888 40000 45008 0 FreeSans 480 0 0 0 u_wb_ack_mxed
port 180 nsew signal tristate
flabel metal3 s 39200 14288 40000 14408 0 FreeSans 480 0 0 0 u_wb_adr[0]
port 181 nsew signal input
flabel metal2 s 29642 0 29698 800 0 FreeSans 224 90 0 0 u_wb_adr[10]
port 182 nsew signal input
flabel metal3 s 39200 46248 40000 46368 0 FreeSans 480 0 0 0 u_wb_adr[11]
port 183 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 u_wb_adr[12]
port 184 nsew signal input
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 u_wb_adr[13]
port 185 nsew signal input
flabel metal3 s 0 46928 800 47048 0 FreeSans 480 0 0 0 u_wb_adr[14]
port 186 nsew signal input
flabel metal2 s 38014 0 38070 800 0 FreeSans 224 90 0 0 u_wb_adr[15]
port 187 nsew signal input
flabel metal3 s 39200 8848 40000 8968 0 FreeSans 480 0 0 0 u_wb_adr[16]
port 188 nsew signal input
flabel metal2 s 23846 49200 23902 50000 0 FreeSans 224 90 0 0 u_wb_adr[17]
port 189 nsew signal input
flabel metal3 s 39200 33328 40000 33448 0 FreeSans 480 0 0 0 u_wb_adr[18]
port 190 nsew signal input
flabel metal2 s 2594 49200 2650 50000 0 FreeSans 224 90 0 0 u_wb_adr[19]
port 191 nsew signal input
flabel metal2 s 5170 49200 5226 50000 0 FreeSans 224 90 0 0 u_wb_adr[1]
port 192 nsew signal input
flabel metal2 s 3238 49200 3294 50000 0 FreeSans 224 90 0 0 u_wb_adr[20]
port 193 nsew signal input
flabel metal2 s 1306 0 1362 800 0 FreeSans 224 90 0 0 u_wb_adr[21]
port 194 nsew signal input
flabel metal2 s 7746 0 7802 800 0 FreeSans 224 90 0 0 u_wb_adr[22]
port 195 nsew signal input
flabel metal3 s 39200 20408 40000 20528 0 FreeSans 480 0 0 0 u_wb_adr[23]
port 196 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 u_wb_adr[2]
port 197 nsew signal input
flabel metal2 s 36082 49200 36138 50000 0 FreeSans 224 90 0 0 u_wb_adr[3]
port 198 nsew signal input
flabel metal3 s 39200 43528 40000 43648 0 FreeSans 480 0 0 0 u_wb_adr[4]
port 199 nsew signal input
flabel metal2 s 11610 49200 11666 50000 0 FreeSans 224 90 0 0 u_wb_adr[5]
port 200 nsew signal input
flabel metal2 s 5814 0 5870 800 0 FreeSans 224 90 0 0 u_wb_adr[6]
port 201 nsew signal input
flabel metal3 s 39200 24488 40000 24608 0 FreeSans 480 0 0 0 u_wb_adr[7]
port 202 nsew signal input
flabel metal3 s 39200 42848 40000 42968 0 FreeSans 480 0 0 0 u_wb_adr[8]
port 203 nsew signal input
flabel metal3 s 0 41488 800 41608 0 FreeSans 480 0 0 0 u_wb_adr[9]
port 204 nsew signal input
flabel metal3 s 39200 31968 40000 32088 0 FreeSans 480 0 0 0 u_wb_cyc
port 205 nsew signal input
flabel metal3 s 39200 13608 40000 13728 0 FreeSans 480 0 0 0 u_wb_err
port 206 nsew signal tristate
flabel metal2 s 27066 0 27122 800 0 FreeSans 224 90 0 0 u_wb_err_cc
port 207 nsew signal input
flabel metal3 s 39200 48968 40000 49088 0 FreeSans 480 0 0 0 u_wb_i_dat[0]
port 208 nsew signal tristate
flabel metal2 s 16762 49200 16818 50000 0 FreeSans 224 90 0 0 u_wb_i_dat[10]
port 209 nsew signal tristate
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 u_wb_i_dat[11]
port 210 nsew signal tristate
flabel metal3 s 0 25848 800 25968 0 FreeSans 480 0 0 0 u_wb_i_dat[12]
port 211 nsew signal tristate
flabel metal3 s 0 19048 800 19168 0 FreeSans 480 0 0 0 u_wb_i_dat[13]
port 212 nsew signal tristate
flabel metal3 s 39200 12928 40000 13048 0 FreeSans 480 0 0 0 u_wb_i_dat[14]
port 213 nsew signal tristate
flabel metal3 s 0 36048 800 36168 0 FreeSans 480 0 0 0 u_wb_i_dat[15]
port 214 nsew signal tristate
flabel metal3 s 39200 2048 40000 2168 0 FreeSans 480 0 0 0 u_wb_i_dat[1]
port 215 nsew signal tristate
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 u_wb_i_dat[2]
port 216 nsew signal tristate
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 u_wb_i_dat[3]
port 217 nsew signal tristate
flabel metal3 s 39200 19728 40000 19848 0 FreeSans 480 0 0 0 u_wb_i_dat[4]
port 218 nsew signal tristate
flabel metal2 s 36726 49200 36782 50000 0 FreeSans 224 90 0 0 u_wb_i_dat[5]
port 219 nsew signal tristate
flabel metal3 s 39200 39448 40000 39568 0 FreeSans 480 0 0 0 u_wb_i_dat[6]
port 220 nsew signal tristate
flabel metal3 s 39200 2728 40000 2848 0 FreeSans 480 0 0 0 u_wb_i_dat[7]
port 221 nsew signal tristate
flabel metal2 s 3238 0 3294 800 0 FreeSans 224 90 0 0 u_wb_i_dat[8]
port 222 nsew signal tristate
flabel metal3 s 39200 25848 40000 25968 0 FreeSans 480 0 0 0 u_wb_i_dat[9]
port 223 nsew signal tristate
flabel metal2 s 662 0 718 800 0 FreeSans 224 90 0 0 u_wb_i_dat_cc[0]
port 224 nsew signal input
flabel metal3 s 39200 41488 40000 41608 0 FreeSans 480 0 0 0 u_wb_i_dat_cc[10]
port 225 nsew signal input
flabel metal2 s 34150 49200 34206 50000 0 FreeSans 224 90 0 0 u_wb_i_dat_cc[11]
port 226 nsew signal input
flabel metal3 s 39200 6808 40000 6928 0 FreeSans 480 0 0 0 u_wb_i_dat_cc[12]
port 227 nsew signal input
flabel metal2 s 32218 49200 32274 50000 0 FreeSans 224 90 0 0 u_wb_i_dat_cc[13]
port 228 nsew signal input
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 u_wb_i_dat_cc[14]
port 229 nsew signal input
flabel metal3 s 0 21768 800 21888 0 FreeSans 480 0 0 0 u_wb_i_dat_cc[15]
port 230 nsew signal input
flabel metal2 s 27710 0 27766 800 0 FreeSans 224 90 0 0 u_wb_i_dat_cc[1]
port 231 nsew signal input
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 u_wb_i_dat_cc[2]
port 232 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 u_wb_i_dat_cc[3]
port 233 nsew signal input
flabel metal3 s 0 27888 800 28008 0 FreeSans 480 0 0 0 u_wb_i_dat_cc[4]
port 234 nsew signal input
flabel metal3 s 0 44888 800 45008 0 FreeSans 480 0 0 0 u_wb_i_dat_cc[5]
port 235 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 u_wb_i_dat_cc[6]
port 236 nsew signal input
flabel metal3 s 0 21088 800 21208 0 FreeSans 480 0 0 0 u_wb_i_dat_cc[7]
port 237 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 u_wb_i_dat_cc[8]
port 238 nsew signal input
flabel metal2 s 2594 0 2650 800 0 FreeSans 224 90 0 0 u_wb_i_dat_cc[9]
port 239 nsew signal input
flabel metal2 s 21914 49200 21970 50000 0 FreeSans 224 90 0 0 u_wb_o_dat[0]
port 240 nsew signal input
flabel metal2 s 12254 49200 12310 50000 0 FreeSans 224 90 0 0 u_wb_o_dat[10]
port 241 nsew signal input
flabel metal2 s 22558 0 22614 800 0 FreeSans 224 90 0 0 u_wb_o_dat[11]
port 242 nsew signal input
flabel metal2 s 28998 49200 29054 50000 0 FreeSans 224 90 0 0 u_wb_o_dat[12]
port 243 nsew signal input
flabel metal3 s 39200 14968 40000 15088 0 FreeSans 480 0 0 0 u_wb_o_dat[13]
port 244 nsew signal input
flabel metal3 s 0 33328 800 33448 0 FreeSans 480 0 0 0 u_wb_o_dat[14]
port 245 nsew signal input
flabel metal3 s 39200 38088 40000 38208 0 FreeSans 480 0 0 0 u_wb_o_dat[15]
port 246 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 u_wb_o_dat[1]
port 247 nsew signal input
flabel metal2 s 16118 0 16174 800 0 FreeSans 224 90 0 0 u_wb_o_dat[2]
port 248 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 u_wb_o_dat[3]
port 249 nsew signal input
flabel metal3 s 39200 36728 40000 36848 0 FreeSans 480 0 0 0 u_wb_o_dat[4]
port 250 nsew signal input
flabel metal2 s 25778 0 25834 800 0 FreeSans 224 90 0 0 u_wb_o_dat[5]
port 251 nsew signal input
flabel metal2 s 25778 49200 25834 50000 0 FreeSans 224 90 0 0 u_wb_o_dat[6]
port 252 nsew signal input
flabel metal2 s 24490 49200 24546 50000 0 FreeSans 224 90 0 0 u_wb_o_dat[7]
port 253 nsew signal input
flabel metal3 s 0 43528 800 43648 0 FreeSans 480 0 0 0 u_wb_o_dat[8]
port 254 nsew signal input
flabel metal2 s 1306 49200 1362 50000 0 FreeSans 224 90 0 0 u_wb_o_dat[9]
port 255 nsew signal input
flabel metal2 s 31574 0 31630 800 0 FreeSans 224 90 0 0 u_wb_sel[0]
port 256 nsew signal input
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 u_wb_sel[1]
port 257 nsew signal input
flabel metal3 s 0 38088 800 38208 0 FreeSans 480 0 0 0 u_wb_stb
port 258 nsew signal input
flabel metal3 s 39200 26528 40000 26648 0 FreeSans 480 0 0 0 u_wb_we
port 259 nsew signal input
flabel metal4 s 4208 2128 4528 47376 0 FreeSans 1920 90 0 0 vccd1
port 260 nsew power bidirectional
flabel metal4 s 34928 2128 35248 47376 0 FreeSans 1920 90 0 0 vccd1
port 260 nsew power bidirectional
flabel metal4 s 19568 2128 19888 47376 0 FreeSans 1920 90 0 0 vssd1
port 261 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 50000
<< end >>
