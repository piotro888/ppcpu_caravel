magic
tech sky130B
magscale 1 2
timestamp 1663005167
<< viali >>
rect 37289 37417 37323 37451
rect 9689 37349 9723 37383
rect 1961 37281 1995 37315
rect 2421 37281 2455 37315
rect 5825 37281 5859 37315
rect 6377 37281 6411 37315
rect 7113 37281 7147 37315
rect 7573 37281 7607 37315
rect 10149 37281 10183 37315
rect 11989 37281 12023 37315
rect 14105 37281 14139 37315
rect 23673 37281 23707 37315
rect 26341 37281 26375 37315
rect 36645 37281 36679 37315
rect 2697 37213 2731 37247
rect 4169 37213 4203 37247
rect 5549 37213 5583 37247
rect 7849 37213 7883 37247
rect 10425 37213 10459 37247
rect 12265 37213 12299 37247
rect 13369 37213 13403 37247
rect 14657 37213 14691 37247
rect 15301 37213 15335 37247
rect 15945 37213 15979 37247
rect 17141 37213 17175 37247
rect 17877 37213 17911 37247
rect 18705 37213 18739 37247
rect 19349 37213 19383 37247
rect 20085 37213 20119 37247
rect 20821 37213 20855 37247
rect 22293 37213 22327 37247
rect 23213 37213 23247 37247
rect 24593 37213 24627 37247
rect 25237 37213 25271 37247
rect 25881 37213 25915 37247
rect 26985 37213 27019 37247
rect 27813 37213 27847 37247
rect 28457 37213 28491 37247
rect 28917 37213 28951 37247
rect 29745 37213 29779 37247
rect 30389 37213 30423 37247
rect 31033 37213 31067 37247
rect 31493 37213 31527 37247
rect 32321 37213 32355 37247
rect 32965 37213 32999 37247
rect 33609 37213 33643 37247
rect 34069 37213 34103 37247
rect 34897 37213 34931 37247
rect 35541 37213 35575 37247
rect 36185 37213 36219 37247
rect 37841 37213 37875 37247
rect 3985 37077 4019 37111
rect 13553 37077 13587 37111
rect 14841 37077 14875 37111
rect 15485 37077 15519 37111
rect 16129 37077 16163 37111
rect 17325 37077 17359 37111
rect 18061 37077 18095 37111
rect 18521 37077 18555 37111
rect 19533 37077 19567 37111
rect 20269 37077 20303 37111
rect 21005 37077 21039 37111
rect 22477 37077 22511 37111
rect 23029 37077 23063 37111
rect 24409 37077 24443 37111
rect 25053 37077 25087 37111
rect 25697 37077 25731 37111
rect 27169 37077 27203 37111
rect 27629 37077 27663 37111
rect 28273 37077 28307 37111
rect 29561 37077 29595 37111
rect 30205 37077 30239 37111
rect 30849 37077 30883 37111
rect 32137 37077 32171 37111
rect 32781 37077 32815 37111
rect 33425 37077 33459 37111
rect 34713 37077 34747 37111
rect 35357 37077 35391 37111
rect 36001 37077 36035 37111
rect 38025 37077 38059 37111
rect 14933 36873 14967 36907
rect 15577 36873 15611 36907
rect 16129 36873 16163 36907
rect 17049 36873 17083 36907
rect 17785 36873 17819 36907
rect 18613 36873 18647 36907
rect 19257 36873 19291 36907
rect 19993 36873 20027 36907
rect 20729 36873 20763 36907
rect 24225 36873 24259 36907
rect 24869 36873 24903 36907
rect 25513 36873 25547 36907
rect 26985 36873 27019 36907
rect 27629 36873 27663 36907
rect 30021 36873 30055 36907
rect 30665 36873 30699 36907
rect 32229 36873 32263 36907
rect 32689 36873 32723 36907
rect 34529 36873 34563 36907
rect 36277 36873 36311 36907
rect 37289 36873 37323 36907
rect 2697 36737 2731 36771
rect 3157 36737 3191 36771
rect 4629 36737 4663 36771
rect 6837 36737 6871 36771
rect 8309 36737 8343 36771
rect 9781 36737 9815 36771
rect 11529 36737 11563 36771
rect 12817 36737 12851 36771
rect 13737 36737 13771 36771
rect 14197 36737 14231 36771
rect 21833 36737 21867 36771
rect 22477 36737 22511 36771
rect 26157 36737 26191 36771
rect 31309 36737 31343 36771
rect 34989 36737 35023 36771
rect 35633 36737 35667 36771
rect 36461 36737 36495 36771
rect 37841 36737 37875 36771
rect 3433 36669 3467 36703
rect 4905 36669 4939 36703
rect 7113 36669 7147 36703
rect 8585 36669 8619 36703
rect 10057 36669 10091 36703
rect 11805 36669 11839 36703
rect 35817 36601 35851 36635
rect 38025 36601 38059 36635
rect 13001 36533 13035 36567
rect 14381 36533 14415 36567
rect 22017 36533 22051 36567
rect 25973 36533 26007 36567
rect 29377 36533 29411 36567
rect 31125 36533 31159 36567
rect 35173 36533 35207 36567
rect 4537 36329 4571 36363
rect 4997 36329 5031 36363
rect 7389 36329 7423 36363
rect 8217 36329 8251 36363
rect 10333 36329 10367 36363
rect 11345 36329 11379 36363
rect 11897 36329 11931 36363
rect 12633 36329 12667 36363
rect 35357 36329 35391 36363
rect 5641 36193 5675 36227
rect 6101 36193 6135 36227
rect 9045 36193 9079 36227
rect 34805 36193 34839 36227
rect 38117 36193 38151 36227
rect 6377 36125 6411 36159
rect 9321 36125 9355 36159
rect 35817 36125 35851 36159
rect 37841 36125 37875 36159
rect 36461 36057 36495 36091
rect 36001 35989 36035 36023
rect 8953 35785 8987 35819
rect 35633 35785 35667 35819
rect 36185 35785 36219 35819
rect 37841 35649 37875 35683
rect 36645 35581 36679 35615
rect 38025 35513 38059 35547
rect 35081 35445 35115 35479
rect 37289 35445 37323 35479
rect 36829 35037 36863 35071
rect 37749 35037 37783 35071
rect 37933 35037 37967 35071
rect 35725 34901 35759 34935
rect 36277 34901 36311 34935
rect 37013 34901 37047 34935
rect 37565 34901 37599 34935
rect 35449 34697 35483 34731
rect 36093 34697 36127 34731
rect 37473 34697 37507 34731
rect 35909 34561 35943 34595
rect 36553 34561 36587 34595
rect 37749 34561 37783 34595
rect 37841 34561 37875 34595
rect 37933 34561 37967 34595
rect 38117 34561 38151 34595
rect 36645 34493 36679 34527
rect 37841 34153 37875 34187
rect 36001 34017 36035 34051
rect 37197 34017 37231 34051
rect 37381 34017 37415 34051
rect 36277 33949 36311 33983
rect 37473 33949 37507 33983
rect 35449 33813 35483 33847
rect 36185 33813 36219 33847
rect 36645 33813 36679 33847
rect 36737 33609 36771 33643
rect 37289 33609 37323 33643
rect 37933 33609 37967 33643
rect 36553 33473 36587 33507
rect 37749 33473 37783 33507
rect 37657 33405 37691 33439
rect 34989 33269 35023 33303
rect 36001 33269 36035 33303
rect 37289 33065 37323 33099
rect 35909 32997 35943 33031
rect 36553 32997 36587 33031
rect 35265 32929 35299 32963
rect 35541 32861 35575 32895
rect 36369 32861 36403 32895
rect 37105 32861 37139 32895
rect 37841 32861 37875 32895
rect 35449 32793 35483 32827
rect 38025 32725 38059 32759
rect 34805 32521 34839 32555
rect 35173 32521 35207 32555
rect 35817 32521 35851 32555
rect 35633 32385 35667 32419
rect 37841 32385 37875 32419
rect 34529 32317 34563 32351
rect 34713 32317 34747 32351
rect 37289 32249 37323 32283
rect 33885 32181 33919 32215
rect 38025 32181 38059 32215
rect 35357 31977 35391 32011
rect 38117 31977 38151 32011
rect 34161 31909 34195 31943
rect 34897 31909 34931 31943
rect 33609 31841 33643 31875
rect 34713 31773 34747 31807
rect 33793 31705 33827 31739
rect 33701 31637 33735 31671
rect 37841 31297 37875 31331
rect 34897 31161 34931 31195
rect 38025 31161 38059 31195
rect 34253 31093 34287 31127
rect 37841 30685 37875 30719
rect 33149 30549 33183 30583
rect 38025 30549 38059 30583
rect 32597 30277 32631 30311
rect 33425 30209 33459 30243
rect 34069 30209 34103 30243
rect 37841 30209 37875 30243
rect 32321 30141 32355 30175
rect 32505 30141 32539 30175
rect 32965 30073 32999 30107
rect 33609 30073 33643 30107
rect 34253 30005 34287 30039
rect 38025 30005 38059 30039
rect 33517 29801 33551 29835
rect 31677 29665 31711 29699
rect 32873 29665 32907 29699
rect 31953 29597 31987 29631
rect 33149 29597 33183 29631
rect 37841 29597 37875 29631
rect 31861 29529 31895 29563
rect 33977 29529 34011 29563
rect 32321 29461 32355 29495
rect 33057 29461 33091 29495
rect 38025 29461 38059 29495
rect 31125 29257 31159 29291
rect 31493 29257 31527 29291
rect 32321 29257 32355 29291
rect 32137 29121 32171 29155
rect 32781 29121 32815 29155
rect 30849 29053 30883 29087
rect 31033 29053 31067 29087
rect 32965 28985 32999 29019
rect 33609 28985 33643 29019
rect 31401 28645 31435 28679
rect 30205 28577 30239 28611
rect 30297 28577 30331 28611
rect 31861 28577 31895 28611
rect 30389 28509 30423 28543
rect 31217 28509 31251 28543
rect 37841 28509 37875 28543
rect 30757 28373 30791 28407
rect 32413 28373 32447 28407
rect 38025 28373 38059 28407
rect 28273 28169 28307 28203
rect 29653 28169 29687 28203
rect 31493 28169 31527 28203
rect 28181 28033 28215 28067
rect 30573 28033 30607 28067
rect 37841 28033 37875 28067
rect 29377 27965 29411 27999
rect 29561 27965 29595 27999
rect 30757 27897 30791 27931
rect 30021 27829 30055 27863
rect 38025 27829 38059 27863
rect 28733 27625 28767 27659
rect 30113 27557 30147 27591
rect 30573 27489 30607 27523
rect 29929 27421 29963 27455
rect 37841 27421 37875 27455
rect 38025 27285 38059 27319
rect 28917 27081 28951 27115
rect 29285 27081 29319 27115
rect 29929 27081 29963 27115
rect 29745 26945 29779 26979
rect 37841 26945 37875 26979
rect 28641 26877 28675 26911
rect 28825 26877 28859 26911
rect 30389 26877 30423 26911
rect 38025 26741 38059 26775
rect 27997 26401 28031 26435
rect 28181 26333 28215 26367
rect 28089 26265 28123 26299
rect 29561 26265 29595 26299
rect 28549 26197 28583 26231
rect 27353 25993 27387 26027
rect 29009 25993 29043 26027
rect 27261 25925 27295 25959
rect 29469 25925 29503 25959
rect 28181 25857 28215 25891
rect 28825 25857 28859 25891
rect 37841 25857 37875 25891
rect 27169 25789 27203 25823
rect 28365 25721 28399 25755
rect 38025 25721 38059 25755
rect 27721 25653 27755 25687
rect 27905 25449 27939 25483
rect 27353 25313 27387 25347
rect 27537 25245 27571 25279
rect 28365 25245 28399 25279
rect 37841 25245 37875 25279
rect 27445 25109 27479 25143
rect 28549 25109 28583 25143
rect 38025 25109 38059 25143
rect 37841 24769 37875 24803
rect 26249 24565 26283 24599
rect 27997 24565 28031 24599
rect 38025 24565 38059 24599
rect 26801 24361 26835 24395
rect 26157 24293 26191 24327
rect 25513 24225 25547 24259
rect 25789 24157 25823 24191
rect 26617 24157 26651 24191
rect 37841 24157 37875 24191
rect 25697 24021 25731 24055
rect 38025 24021 38059 24055
rect 25237 23817 25271 23851
rect 25605 23817 25639 23851
rect 26065 23681 26099 23715
rect 24961 23613 24995 23647
rect 25145 23613 25179 23647
rect 23581 23545 23615 23579
rect 26249 23477 26283 23511
rect 36829 23273 36863 23307
rect 24501 23137 24535 23171
rect 24685 23137 24719 23171
rect 23029 23069 23063 23103
rect 24777 23069 24811 23103
rect 25605 23069 25639 23103
rect 37013 23069 37047 23103
rect 37841 23069 37875 23103
rect 23121 22933 23155 22967
rect 25145 22933 25179 22967
rect 25789 22933 25823 22967
rect 26249 22933 26283 22967
rect 38025 22933 38059 22967
rect 23765 22729 23799 22763
rect 24133 22729 24167 22763
rect 36369 22729 36403 22763
rect 36737 22729 36771 22763
rect 24593 22593 24627 22627
rect 37841 22593 37875 22627
rect 23489 22525 23523 22559
rect 23673 22525 23707 22559
rect 36093 22525 36127 22559
rect 36277 22525 36311 22559
rect 37289 22525 37323 22559
rect 24777 22457 24811 22491
rect 25237 22389 25271 22423
rect 35449 22389 35483 22423
rect 38025 22389 38059 22423
rect 22477 21981 22511 22015
rect 37841 21981 37875 22015
rect 22293 21845 22327 21879
rect 23489 21845 23523 21879
rect 24501 21845 24535 21879
rect 38025 21845 38059 21879
rect 23029 21641 23063 21675
rect 23397 21641 23431 21675
rect 23857 21505 23891 21539
rect 37473 21505 37507 21539
rect 38117 21505 38151 21539
rect 22753 21437 22787 21471
rect 22937 21437 22971 21471
rect 24041 21301 24075 21335
rect 37933 21301 37967 21335
rect 22385 21097 22419 21131
rect 23765 21097 23799 21131
rect 22293 21029 22327 21063
rect 21925 20893 21959 20927
rect 22937 20893 22971 20927
rect 23029 20893 23063 20927
rect 23213 20757 23247 20791
rect 22201 20553 22235 20587
rect 23765 20553 23799 20587
rect 23213 20417 23247 20451
rect 37841 20417 37875 20451
rect 22293 20349 22327 20383
rect 22385 20349 22419 20383
rect 38025 20281 38059 20315
rect 21833 20213 21867 20247
rect 23029 20213 23063 20247
rect 19901 20009 19935 20043
rect 20545 19873 20579 19907
rect 20821 19805 20855 19839
rect 21833 19805 21867 19839
rect 37841 19805 37875 19839
rect 20729 19669 20763 19703
rect 21189 19669 21223 19703
rect 22017 19669 22051 19703
rect 38025 19669 38059 19703
rect 21281 19465 21315 19499
rect 19625 19397 19659 19431
rect 21097 19329 21131 19363
rect 37841 19329 37875 19363
rect 20545 19261 20579 19295
rect 19349 19125 19383 19159
rect 38025 19125 38059 19159
rect 19809 18785 19843 18819
rect 19993 18717 20027 18751
rect 20913 18717 20947 18751
rect 37841 18717 37875 18751
rect 20085 18581 20119 18615
rect 20453 18581 20487 18615
rect 21097 18581 21131 18615
rect 38025 18581 38059 18615
rect 18245 18377 18279 18411
rect 19441 18377 19475 18411
rect 19809 18377 19843 18411
rect 20269 18241 20303 18275
rect 18061 18173 18095 18207
rect 18153 18173 18187 18207
rect 19165 18173 19199 18207
rect 19349 18173 19383 18207
rect 18613 18037 18647 18071
rect 20453 18037 20487 18071
rect 18613 17833 18647 17867
rect 19993 17833 20027 17867
rect 19349 17629 19383 17663
rect 37841 17629 37875 17663
rect 37289 17561 37323 17595
rect 19533 17493 19567 17527
rect 38025 17493 38059 17527
rect 18153 17153 18187 17187
rect 37841 17153 37875 17187
rect 18337 16949 18371 16983
rect 37289 16949 37323 16983
rect 38025 16949 38059 16983
rect 18337 16745 18371 16779
rect 20913 16745 20947 16779
rect 17785 16609 17819 16643
rect 17877 16609 17911 16643
rect 20453 16541 20487 16575
rect 37841 16541 37875 16575
rect 17969 16473 18003 16507
rect 19257 16473 19291 16507
rect 20177 16473 20211 16507
rect 37289 16405 37323 16439
rect 38025 16405 38059 16439
rect 17509 16201 17543 16235
rect 17141 16065 17175 16099
rect 17969 16065 18003 16099
rect 37841 16065 37875 16099
rect 16957 15997 16991 16031
rect 17049 15997 17083 16031
rect 18153 15861 18187 15895
rect 37289 15861 37323 15895
rect 38025 15861 38059 15895
rect 17877 15657 17911 15691
rect 16773 15589 16807 15623
rect 16221 15521 16255 15555
rect 16405 15453 16439 15487
rect 17233 15453 17267 15487
rect 16313 15317 16347 15351
rect 17417 15317 17451 15351
rect 15761 15113 15795 15147
rect 17325 15113 17359 15147
rect 15669 14977 15703 15011
rect 16681 14977 16715 15011
rect 37841 14977 37875 15011
rect 15577 14909 15611 14943
rect 16129 14841 16163 14875
rect 16865 14841 16899 14875
rect 38025 14841 38059 14875
rect 37289 14773 37323 14807
rect 16497 14569 16531 14603
rect 15393 14501 15427 14535
rect 14841 14433 14875 14467
rect 15025 14365 15059 14399
rect 15853 14365 15887 14399
rect 37841 14365 37875 14399
rect 14933 14229 14967 14263
rect 16037 14229 16071 14263
rect 37289 14229 37323 14263
rect 38025 14229 38059 14263
rect 14933 14025 14967 14059
rect 15485 14025 15519 14059
rect 12357 13889 12391 13923
rect 37289 13889 37323 13923
rect 37841 13889 37875 13923
rect 12081 13821 12115 13855
rect 38025 13685 38059 13719
rect 12081 13481 12115 13515
rect 15485 13481 15519 13515
rect 12265 13413 12299 13447
rect 12541 13345 12575 13379
rect 14289 13345 14323 13379
rect 14473 13277 14507 13311
rect 15301 13277 15335 13311
rect 37841 13277 37875 13311
rect 13001 13141 13035 13175
rect 14381 13141 14415 13175
rect 14841 13141 14875 13175
rect 37289 13141 37323 13175
rect 38025 13141 38059 13175
rect 12633 12937 12667 12971
rect 13553 12937 13587 12971
rect 13921 12937 13955 12971
rect 14381 12801 14415 12835
rect 13369 12733 13403 12767
rect 13461 12733 13495 12767
rect 15025 12733 15059 12767
rect 14565 12665 14599 12699
rect 12817 12257 12851 12291
rect 14749 12257 14783 12291
rect 13001 12189 13035 12223
rect 14105 12189 14139 12223
rect 37841 12189 37875 12223
rect 12909 12121 12943 12155
rect 13369 12053 13403 12087
rect 14289 12053 14323 12087
rect 37289 12053 37323 12087
rect 38025 12053 38059 12087
rect 12173 11849 12207 11883
rect 13001 11849 13035 11883
rect 13369 11849 13403 11883
rect 13829 11713 13863 11747
rect 37841 11713 37875 11747
rect 12817 11645 12851 11679
rect 12909 11645 12943 11679
rect 14013 11509 14047 11543
rect 37289 11509 37323 11543
rect 38025 11509 38059 11543
rect 11989 11305 12023 11339
rect 13185 11237 13219 11271
rect 14289 11237 14323 11271
rect 38025 11237 38059 11271
rect 12633 11169 12667 11203
rect 12817 11101 12851 11135
rect 14105 11101 14139 11135
rect 37289 11101 37323 11135
rect 37841 11101 37875 11135
rect 11345 11033 11379 11067
rect 12725 11033 12759 11067
rect 10425 10761 10459 10795
rect 11897 10761 11931 10795
rect 9873 10693 9907 10727
rect 11805 10625 11839 10659
rect 12725 10625 12759 10659
rect 12909 10625 12943 10659
rect 13093 10625 13127 10659
rect 13737 10625 13771 10659
rect 37841 10625 37875 10659
rect 10977 10557 11011 10591
rect 11713 10557 11747 10591
rect 14289 10489 14323 10523
rect 12265 10421 12299 10455
rect 13553 10421 13587 10455
rect 14749 10421 14783 10455
rect 37289 10421 37323 10455
rect 38025 10421 38059 10455
rect 10793 10149 10827 10183
rect 9597 10081 9631 10115
rect 10149 10081 10183 10115
rect 11253 10081 11287 10115
rect 13093 10081 13127 10115
rect 14105 10081 14139 10115
rect 10425 10013 10459 10047
rect 11529 10013 11563 10047
rect 12909 9945 12943 9979
rect 10333 9877 10367 9911
rect 12541 9877 12575 9911
rect 13001 9877 13035 9911
rect 9321 9605 9355 9639
rect 11989 9605 12023 9639
rect 12541 9537 12575 9571
rect 37841 9537 37875 9571
rect 9137 9469 9171 9503
rect 9229 9469 9263 9503
rect 10149 9469 10183 9503
rect 10425 9469 10459 9503
rect 12817 9469 12851 9503
rect 9689 9401 9723 9435
rect 37289 9401 37323 9435
rect 38025 9401 38059 9435
rect 9597 9129 9631 9163
rect 12633 8993 12667 9027
rect 10057 8925 10091 8959
rect 10333 8925 10367 8959
rect 12357 8925 12391 8959
rect 37841 8925 37875 8959
rect 37289 8857 37323 8891
rect 38025 8789 38059 8823
rect 9229 8585 9263 8619
rect 9597 8585 9631 8619
rect 10057 8517 10091 8551
rect 37841 8449 37875 8483
rect 8401 8381 8435 8415
rect 8953 8381 8987 8415
rect 9137 8381 9171 8415
rect 37289 8381 37323 8415
rect 10609 8313 10643 8347
rect 38025 8313 38059 8347
rect 8953 8041 8987 8075
rect 8401 7973 8435 8007
rect 7849 7905 7883 7939
rect 9505 7905 9539 7939
rect 9781 7905 9815 7939
rect 8033 7837 8067 7871
rect 37841 7837 37875 7871
rect 7941 7701 7975 7735
rect 37289 7701 37323 7735
rect 38025 7701 38059 7735
rect 8217 7497 8251 7531
rect 10425 7497 10459 7531
rect 7389 7293 7423 7327
rect 7941 7293 7975 7327
rect 8125 7293 8159 7327
rect 9137 7293 9171 7327
rect 9413 7293 9447 7327
rect 8585 7225 8619 7259
rect 6561 6817 6595 6851
rect 7205 6817 7239 6851
rect 7849 6817 7883 6851
rect 9229 6817 9263 6851
rect 8033 6749 8067 6783
rect 8953 6749 8987 6783
rect 10241 6749 10275 6783
rect 10517 6749 10551 6783
rect 37289 6749 37323 6783
rect 37841 6749 37875 6783
rect 7941 6681 7975 6715
rect 8401 6613 8435 6647
rect 38025 6613 38059 6647
rect 7113 6409 7147 6443
rect 8033 6409 8067 6443
rect 8401 6409 8435 6443
rect 10149 6409 10183 6443
rect 37289 6409 37323 6443
rect 7941 6273 7975 6307
rect 8861 6273 8895 6307
rect 37841 6273 37875 6307
rect 7757 6205 7791 6239
rect 9137 6205 9171 6239
rect 38025 6069 38059 6103
rect 8309 5865 8343 5899
rect 37289 5865 37323 5899
rect 7757 5729 7791 5763
rect 7113 5661 7147 5695
rect 7941 5661 7975 5695
rect 8953 5661 8987 5695
rect 9229 5661 9263 5695
rect 37841 5661 37875 5695
rect 7849 5525 7883 5559
rect 38025 5525 38059 5559
rect 8309 5321 8343 5355
rect 9413 5321 9447 5355
rect 7113 5253 7147 5287
rect 7941 5253 7975 5287
rect 8861 5253 8895 5287
rect 7849 5185 7883 5219
rect 37289 5185 37323 5219
rect 37841 5185 37875 5219
rect 7757 5117 7791 5151
rect 38025 4981 38059 5015
rect 36829 4437 36863 4471
rect 37565 4437 37599 4471
rect 38025 4437 38059 4471
rect 38025 4165 38059 4199
rect 37841 4097 37875 4131
rect 37289 3961 37323 3995
rect 34713 3893 34747 3927
rect 36185 3893 36219 3927
rect 36645 3893 36679 3927
rect 35081 3553 35115 3587
rect 36553 3553 36587 3587
rect 34805 3485 34839 3519
rect 36277 3485 36311 3519
rect 37841 3485 37875 3519
rect 5273 3349 5307 3383
rect 30297 3349 30331 3383
rect 31953 3349 31987 3383
rect 33241 3349 33275 3383
rect 38025 3349 38059 3383
rect 4813 3145 4847 3179
rect 9229 3145 9263 3179
rect 14381 3145 14415 3179
rect 22017 3145 22051 3179
rect 23029 3145 23063 3179
rect 26157 3145 26191 3179
rect 29101 3145 29135 3179
rect 37933 3145 37967 3179
rect 4169 3009 4203 3043
rect 4629 3009 4663 3043
rect 8585 3009 8619 3043
rect 9045 3009 9079 3043
rect 13737 3009 13771 3043
rect 14197 3009 14231 3043
rect 21833 3009 21867 3043
rect 22477 3009 22511 3043
rect 25513 3009 25547 3043
rect 25973 3009 26007 3043
rect 28917 3009 28951 3043
rect 29561 3009 29595 3043
rect 30665 3009 30699 3043
rect 32413 3009 32447 3043
rect 33701 3009 33735 3043
rect 34989 3009 35023 3043
rect 36461 3009 36495 3043
rect 37841 3009 37875 3043
rect 30389 2941 30423 2975
rect 32137 2941 32171 2975
rect 33425 2941 33459 2975
rect 34713 2941 34747 2975
rect 3341 2805 3375 2839
rect 5825 2805 5859 2839
rect 6745 2805 6779 2839
rect 7481 2805 7515 2839
rect 9781 2805 9815 2839
rect 10425 2805 10459 2839
rect 10977 2805 11011 2839
rect 11897 2805 11931 2839
rect 12633 2805 12667 2839
rect 14933 2805 14967 2839
rect 15577 2805 15611 2839
rect 16129 2805 16163 2839
rect 17049 2805 17083 2839
rect 17785 2805 17819 2839
rect 18613 2805 18647 2839
rect 19257 2805 19291 2839
rect 19993 2805 20027 2839
rect 20729 2805 20763 2839
rect 24225 2805 24259 2839
rect 24869 2805 24903 2839
rect 26985 2805 27019 2839
rect 27629 2805 27663 2839
rect 36645 2805 36679 2839
rect 5181 2601 5215 2635
rect 5825 2601 5859 2635
rect 8217 2601 8251 2635
rect 9505 2601 9539 2635
rect 10333 2601 10367 2635
rect 12909 2601 12943 2635
rect 13553 2601 13587 2635
rect 14841 2601 14875 2635
rect 15485 2601 15519 2635
rect 16129 2601 16163 2635
rect 17325 2601 17359 2635
rect 18061 2601 18095 2635
rect 18521 2601 18555 2635
rect 20085 2601 20119 2635
rect 20821 2601 20855 2635
rect 23213 2601 23247 2635
rect 24593 2601 24627 2635
rect 25237 2601 25271 2635
rect 25881 2601 25915 2635
rect 27169 2601 27203 2635
rect 27813 2601 27847 2635
rect 28457 2601 28491 2635
rect 36553 2601 36587 2635
rect 3249 2533 3283 2567
rect 7021 2533 7055 2567
rect 7757 2533 7791 2567
rect 12173 2533 12207 2567
rect 19533 2533 19567 2567
rect 33609 2533 33643 2567
rect 30205 2465 30239 2499
rect 32413 2465 32447 2499
rect 34989 2465 35023 2499
rect 36001 2465 36035 2499
rect 37289 2465 37323 2499
rect 1961 2397 1995 2431
rect 2421 2397 2455 2431
rect 3065 2397 3099 2431
rect 4169 2397 4203 2431
rect 4997 2397 5031 2431
rect 5641 2397 5675 2431
rect 6837 2397 6871 2431
rect 7573 2397 7607 2431
rect 8401 2397 8435 2431
rect 8953 2397 8987 2431
rect 9689 2397 9723 2431
rect 10149 2397 10183 2431
rect 10793 2397 10827 2431
rect 11989 2397 12023 2431
rect 12725 2397 12759 2431
rect 13369 2397 13403 2431
rect 14105 2397 14139 2431
rect 14657 2397 14691 2431
rect 15301 2397 15335 2431
rect 15945 2397 15979 2431
rect 17141 2397 17175 2431
rect 17877 2397 17911 2431
rect 18705 2397 18739 2431
rect 19349 2397 19383 2431
rect 20269 2397 20303 2431
rect 21005 2397 21039 2431
rect 22569 2397 22603 2431
rect 23029 2397 23063 2431
rect 23673 2397 23707 2431
rect 24409 2397 24443 2431
rect 25053 2397 25087 2431
rect 25697 2397 25731 2431
rect 26341 2397 26375 2431
rect 26985 2397 27019 2431
rect 27629 2397 27663 2431
rect 28273 2397 28307 2431
rect 28917 2397 28951 2431
rect 30481 2397 30515 2431
rect 30941 2397 30975 2431
rect 32137 2397 32171 2431
rect 34713 2397 34747 2431
rect 36737 2397 36771 2431
rect 37565 2397 37599 2431
rect 2605 2261 2639 2295
rect 3985 2261 4019 2295
rect 10977 2261 11011 2295
rect 22385 2261 22419 2295
rect 31493 2261 31527 2295
rect 34069 2261 34103 2295
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 36170 37408 36176 37460
rect 36228 37448 36234 37460
rect 37277 37451 37335 37457
rect 37277 37448 37289 37451
rect 36228 37420 37289 37448
rect 36228 37408 36234 37420
rect 37277 37417 37289 37420
rect 37323 37417 37335 37451
rect 37277 37411 37335 37417
rect 9677 37383 9735 37389
rect 9677 37349 9689 37383
rect 9723 37380 9735 37383
rect 10410 37380 10416 37392
rect 9723 37352 10416 37380
rect 9723 37349 9735 37352
rect 9677 37343 9735 37349
rect 1949 37315 2007 37321
rect 1949 37281 1961 37315
rect 1995 37312 2007 37315
rect 2314 37312 2320 37324
rect 1995 37284 2320 37312
rect 1995 37281 2007 37284
rect 1949 37275 2007 37281
rect 2314 37272 2320 37284
rect 2372 37312 2378 37324
rect 2409 37315 2467 37321
rect 2409 37312 2421 37315
rect 2372 37284 2421 37312
rect 2372 37272 2378 37284
rect 2409 37281 2421 37284
rect 2455 37281 2467 37315
rect 2409 37275 2467 37281
rect 5258 37272 5264 37324
rect 5316 37312 5322 37324
rect 5813 37315 5871 37321
rect 5813 37312 5825 37315
rect 5316 37284 5825 37312
rect 5316 37272 5322 37284
rect 5813 37281 5825 37284
rect 5859 37312 5871 37315
rect 6365 37315 6423 37321
rect 6365 37312 6377 37315
rect 5859 37284 6377 37312
rect 5859 37281 5871 37284
rect 5813 37275 5871 37281
rect 6365 37281 6377 37284
rect 6411 37281 6423 37315
rect 6365 37275 6423 37281
rect 7101 37315 7159 37321
rect 7101 37281 7113 37315
rect 7147 37312 7159 37315
rect 7466 37312 7472 37324
rect 7147 37284 7472 37312
rect 7147 37281 7159 37284
rect 7101 37275 7159 37281
rect 7466 37272 7472 37284
rect 7524 37312 7530 37324
rect 10152 37321 10180 37352
rect 10410 37340 10416 37352
rect 10468 37340 10474 37392
rect 7561 37315 7619 37321
rect 7561 37312 7573 37315
rect 7524 37284 7573 37312
rect 7524 37272 7530 37284
rect 7561 37281 7573 37284
rect 7607 37281 7619 37315
rect 7561 37275 7619 37281
rect 10137 37315 10195 37321
rect 10137 37281 10149 37315
rect 10183 37281 10195 37315
rect 10137 37275 10195 37281
rect 11882 37272 11888 37324
rect 11940 37312 11946 37324
rect 11977 37315 12035 37321
rect 11977 37312 11989 37315
rect 11940 37284 11989 37312
rect 11940 37272 11946 37284
rect 11977 37281 11989 37284
rect 12023 37281 12035 37315
rect 14093 37315 14151 37321
rect 14093 37312 14105 37315
rect 11977 37275 12035 37281
rect 13372 37284 14105 37312
rect 13372 37256 13400 37284
rect 14093 37281 14105 37284
rect 14139 37281 14151 37315
rect 23661 37315 23719 37321
rect 23661 37312 23673 37315
rect 14093 37275 14151 37281
rect 23216 37284 23673 37312
rect 2682 37244 2688 37256
rect 2643 37216 2688 37244
rect 2682 37204 2688 37216
rect 2740 37204 2746 37256
rect 4157 37247 4215 37253
rect 4157 37213 4169 37247
rect 4203 37244 4215 37247
rect 4982 37244 4988 37256
rect 4203 37216 4988 37244
rect 4203 37213 4215 37216
rect 4157 37207 4215 37213
rect 4982 37204 4988 37216
rect 5040 37204 5046 37256
rect 5537 37247 5595 37253
rect 5537 37213 5549 37247
rect 5583 37244 5595 37247
rect 6546 37244 6552 37256
rect 5583 37216 6552 37244
rect 5583 37213 5595 37216
rect 5537 37207 5595 37213
rect 6546 37204 6552 37216
rect 6604 37204 6610 37256
rect 7837 37247 7895 37253
rect 7837 37213 7849 37247
rect 7883 37244 7895 37247
rect 8018 37244 8024 37256
rect 7883 37216 8024 37244
rect 7883 37213 7895 37216
rect 7837 37207 7895 37213
rect 8018 37204 8024 37216
rect 8076 37204 8082 37256
rect 10410 37244 10416 37256
rect 10371 37216 10416 37244
rect 10410 37204 10416 37216
rect 10468 37204 10474 37256
rect 12158 37204 12164 37256
rect 12216 37244 12222 37256
rect 12253 37247 12311 37253
rect 12253 37244 12265 37247
rect 12216 37216 12265 37244
rect 12216 37204 12222 37216
rect 12253 37213 12265 37216
rect 12299 37213 12311 37247
rect 13354 37244 13360 37256
rect 13315 37216 13360 37244
rect 12253 37207 12311 37213
rect 13354 37204 13360 37216
rect 13412 37204 13418 37256
rect 14645 37247 14703 37253
rect 14645 37213 14657 37247
rect 14691 37244 14703 37247
rect 14826 37244 14832 37256
rect 14691 37216 14832 37244
rect 14691 37213 14703 37216
rect 14645 37207 14703 37213
rect 14826 37204 14832 37216
rect 14884 37204 14890 37256
rect 15289 37247 15347 37253
rect 15289 37213 15301 37247
rect 15335 37244 15347 37247
rect 15562 37244 15568 37256
rect 15335 37216 15568 37244
rect 15335 37213 15347 37216
rect 15289 37207 15347 37213
rect 15562 37204 15568 37216
rect 15620 37204 15626 37256
rect 15933 37247 15991 37253
rect 15933 37213 15945 37247
rect 15979 37244 15991 37247
rect 16298 37244 16304 37256
rect 15979 37216 16304 37244
rect 15979 37213 15991 37216
rect 15933 37207 15991 37213
rect 16298 37204 16304 37216
rect 16356 37204 16362 37256
rect 17034 37204 17040 37256
rect 17092 37244 17098 37256
rect 17129 37247 17187 37253
rect 17129 37244 17141 37247
rect 17092 37216 17141 37244
rect 17092 37204 17098 37216
rect 17129 37213 17141 37216
rect 17175 37213 17187 37247
rect 17129 37207 17187 37213
rect 17770 37204 17776 37256
rect 17828 37244 17834 37256
rect 17865 37247 17923 37253
rect 17865 37244 17877 37247
rect 17828 37216 17877 37244
rect 17828 37204 17834 37216
rect 17865 37213 17877 37216
rect 17911 37213 17923 37247
rect 17865 37207 17923 37213
rect 18506 37204 18512 37256
rect 18564 37244 18570 37256
rect 18693 37247 18751 37253
rect 18693 37244 18705 37247
rect 18564 37216 18705 37244
rect 18564 37204 18570 37216
rect 18693 37213 18705 37216
rect 18739 37213 18751 37247
rect 18693 37207 18751 37213
rect 19242 37204 19248 37256
rect 19300 37244 19306 37256
rect 19337 37247 19395 37253
rect 19337 37244 19349 37247
rect 19300 37216 19349 37244
rect 19300 37204 19306 37216
rect 19337 37213 19349 37216
rect 19383 37213 19395 37247
rect 19337 37207 19395 37213
rect 19978 37204 19984 37256
rect 20036 37244 20042 37256
rect 20073 37247 20131 37253
rect 20073 37244 20085 37247
rect 20036 37216 20085 37244
rect 20036 37204 20042 37216
rect 20073 37213 20085 37216
rect 20119 37213 20131 37247
rect 20073 37207 20131 37213
rect 20714 37204 20720 37256
rect 20772 37244 20778 37256
rect 20809 37247 20867 37253
rect 20809 37244 20821 37247
rect 20772 37216 20821 37244
rect 20772 37204 20778 37216
rect 20809 37213 20821 37216
rect 20855 37213 20867 37247
rect 22278 37244 22284 37256
rect 22239 37216 22284 37244
rect 20809 37207 20867 37213
rect 22278 37204 22284 37216
rect 22336 37204 22342 37256
rect 22922 37204 22928 37256
rect 22980 37244 22986 37256
rect 23216 37253 23244 37284
rect 23661 37281 23673 37284
rect 23707 37281 23719 37315
rect 23661 37275 23719 37281
rect 25130 37272 25136 37324
rect 25188 37312 25194 37324
rect 26329 37315 26387 37321
rect 26329 37312 26341 37315
rect 25188 37284 26341 37312
rect 25188 37272 25194 37284
rect 23201 37247 23259 37253
rect 23201 37244 23213 37247
rect 22980 37216 23213 37244
rect 22980 37204 22986 37216
rect 23201 37213 23213 37216
rect 23247 37213 23259 37247
rect 24578 37244 24584 37256
rect 24539 37216 24584 37244
rect 23201 37207 23259 37213
rect 24578 37204 24584 37216
rect 24636 37204 24642 37256
rect 24854 37204 24860 37256
rect 24912 37244 24918 37256
rect 25884 37253 25912 37284
rect 26329 37281 26341 37284
rect 26375 37281 26387 37315
rect 26329 37275 26387 37281
rect 34698 37272 34704 37324
rect 34756 37312 34762 37324
rect 36633 37315 36691 37321
rect 36633 37312 36645 37315
rect 34756 37284 36645 37312
rect 34756 37272 34762 37284
rect 25225 37247 25283 37253
rect 25225 37244 25237 37247
rect 24912 37216 25237 37244
rect 24912 37204 24918 37216
rect 25225 37213 25237 37216
rect 25271 37213 25283 37247
rect 25225 37207 25283 37213
rect 25869 37247 25927 37253
rect 25869 37213 25881 37247
rect 25915 37213 25927 37247
rect 25869 37207 25927 37213
rect 26602 37204 26608 37256
rect 26660 37244 26666 37256
rect 26970 37244 26976 37256
rect 26660 37216 26976 37244
rect 26660 37204 26666 37216
rect 26970 37204 26976 37216
rect 27028 37204 27034 37256
rect 27338 37204 27344 37256
rect 27396 37244 27402 37256
rect 27614 37244 27620 37256
rect 27396 37216 27620 37244
rect 27396 37204 27402 37216
rect 27614 37204 27620 37216
rect 27672 37244 27678 37256
rect 27801 37247 27859 37253
rect 27801 37244 27813 37247
rect 27672 37216 27813 37244
rect 27672 37204 27678 37216
rect 27801 37213 27813 37216
rect 27847 37213 27859 37247
rect 27801 37207 27859 37213
rect 28074 37204 28080 37256
rect 28132 37244 28138 37256
rect 28445 37247 28503 37253
rect 28445 37244 28457 37247
rect 28132 37216 28457 37244
rect 28132 37204 28138 37216
rect 28445 37213 28457 37216
rect 28491 37244 28503 37247
rect 28905 37247 28963 37253
rect 28905 37244 28917 37247
rect 28491 37216 28917 37244
rect 28491 37213 28503 37216
rect 28445 37207 28503 37213
rect 28905 37213 28917 37216
rect 28951 37213 28963 37247
rect 28905 37207 28963 37213
rect 29362 37204 29368 37256
rect 29420 37244 29426 37256
rect 29733 37247 29791 37253
rect 29733 37244 29745 37247
rect 29420 37216 29745 37244
rect 29420 37204 29426 37216
rect 29733 37213 29745 37216
rect 29779 37213 29791 37247
rect 29733 37207 29791 37213
rect 30006 37204 30012 37256
rect 30064 37244 30070 37256
rect 30377 37247 30435 37253
rect 30377 37244 30389 37247
rect 30064 37216 30389 37244
rect 30064 37204 30070 37216
rect 30377 37213 30389 37216
rect 30423 37213 30435 37247
rect 30377 37207 30435 37213
rect 30466 37204 30472 37256
rect 30524 37244 30530 37256
rect 31021 37247 31079 37253
rect 31021 37244 31033 37247
rect 30524 37216 31033 37244
rect 30524 37204 30530 37216
rect 31021 37213 31033 37216
rect 31067 37244 31079 37247
rect 31481 37247 31539 37253
rect 31481 37244 31493 37247
rect 31067 37216 31493 37244
rect 31067 37213 31079 37216
rect 31021 37207 31079 37213
rect 31481 37213 31493 37216
rect 31527 37213 31539 37247
rect 31481 37207 31539 37213
rect 31754 37204 31760 37256
rect 31812 37244 31818 37256
rect 32214 37244 32220 37256
rect 31812 37216 32220 37244
rect 31812 37204 31818 37216
rect 32214 37204 32220 37216
rect 32272 37244 32278 37256
rect 32309 37247 32367 37253
rect 32309 37244 32321 37247
rect 32272 37216 32321 37244
rect 32272 37204 32278 37216
rect 32309 37213 32321 37216
rect 32355 37213 32367 37247
rect 32309 37207 32367 37213
rect 32490 37204 32496 37256
rect 32548 37244 32554 37256
rect 32953 37247 33011 37253
rect 32953 37244 32965 37247
rect 32548 37216 32965 37244
rect 32548 37204 32554 37216
rect 32953 37213 32965 37216
rect 32999 37213 33011 37247
rect 32953 37207 33011 37213
rect 33226 37204 33232 37256
rect 33284 37244 33290 37256
rect 33597 37247 33655 37253
rect 33597 37244 33609 37247
rect 33284 37216 33609 37244
rect 33284 37204 33290 37216
rect 33597 37213 33609 37216
rect 33643 37244 33655 37247
rect 34057 37247 34115 37253
rect 34057 37244 34069 37247
rect 33643 37216 34069 37244
rect 33643 37213 33655 37216
rect 33597 37207 33655 37213
rect 34057 37213 34069 37216
rect 34103 37213 34115 37247
rect 34057 37207 34115 37213
rect 34514 37204 34520 37256
rect 34572 37244 34578 37256
rect 35544 37253 35572 37284
rect 36633 37281 36645 37284
rect 36679 37281 36691 37315
rect 36633 37275 36691 37281
rect 34885 37247 34943 37253
rect 34885 37244 34897 37247
rect 34572 37216 34897 37244
rect 34572 37204 34578 37216
rect 34885 37213 34897 37216
rect 34931 37213 34943 37247
rect 34885 37207 34943 37213
rect 35529 37247 35587 37253
rect 35529 37213 35541 37247
rect 35575 37213 35587 37247
rect 35529 37207 35587 37213
rect 35894 37204 35900 37256
rect 35952 37244 35958 37256
rect 36173 37247 36231 37253
rect 36173 37244 36185 37247
rect 35952 37216 36185 37244
rect 35952 37204 35958 37216
rect 36173 37213 36185 37216
rect 36219 37213 36231 37247
rect 36173 37207 36231 37213
rect 36446 37204 36452 37256
rect 36504 37244 36510 37256
rect 37829 37247 37887 37253
rect 37829 37244 37841 37247
rect 36504 37216 37841 37244
rect 36504 37204 36510 37216
rect 37829 37213 37841 37216
rect 37875 37213 37887 37247
rect 37829 37207 37887 37213
rect 3786 37068 3792 37120
rect 3844 37108 3850 37120
rect 3973 37111 4031 37117
rect 3973 37108 3985 37111
rect 3844 37080 3985 37108
rect 3844 37068 3850 37080
rect 3973 37077 3985 37080
rect 4019 37077 4031 37111
rect 13538 37108 13544 37120
rect 13499 37080 13544 37108
rect 3973 37071 4031 37077
rect 13538 37068 13544 37080
rect 13596 37068 13602 37120
rect 14829 37111 14887 37117
rect 14829 37077 14841 37111
rect 14875 37108 14887 37111
rect 15010 37108 15016 37120
rect 14875 37080 15016 37108
rect 14875 37077 14887 37080
rect 14829 37071 14887 37077
rect 15010 37068 15016 37080
rect 15068 37068 15074 37120
rect 15473 37111 15531 37117
rect 15473 37077 15485 37111
rect 15519 37108 15531 37111
rect 15746 37108 15752 37120
rect 15519 37080 15752 37108
rect 15519 37077 15531 37080
rect 15473 37071 15531 37077
rect 15746 37068 15752 37080
rect 15804 37068 15810 37120
rect 16117 37111 16175 37117
rect 16117 37077 16129 37111
rect 16163 37108 16175 37111
rect 16390 37108 16396 37120
rect 16163 37080 16396 37108
rect 16163 37077 16175 37080
rect 16117 37071 16175 37077
rect 16390 37068 16396 37080
rect 16448 37068 16454 37120
rect 17313 37111 17371 37117
rect 17313 37077 17325 37111
rect 17359 37108 17371 37111
rect 17862 37108 17868 37120
rect 17359 37080 17868 37108
rect 17359 37077 17371 37080
rect 17313 37071 17371 37077
rect 17862 37068 17868 37080
rect 17920 37068 17926 37120
rect 18046 37108 18052 37120
rect 18007 37080 18052 37108
rect 18046 37068 18052 37080
rect 18104 37068 18110 37120
rect 18230 37068 18236 37120
rect 18288 37108 18294 37120
rect 18509 37111 18567 37117
rect 18509 37108 18521 37111
rect 18288 37080 18521 37108
rect 18288 37068 18294 37080
rect 18509 37077 18521 37080
rect 18555 37077 18567 37111
rect 18509 37071 18567 37077
rect 19426 37068 19432 37120
rect 19484 37108 19490 37120
rect 19521 37111 19579 37117
rect 19521 37108 19533 37111
rect 19484 37080 19533 37108
rect 19484 37068 19490 37080
rect 19521 37077 19533 37080
rect 19567 37077 19579 37111
rect 19521 37071 19579 37077
rect 20257 37111 20315 37117
rect 20257 37077 20269 37111
rect 20303 37108 20315 37111
rect 20530 37108 20536 37120
rect 20303 37080 20536 37108
rect 20303 37077 20315 37080
rect 20257 37071 20315 37077
rect 20530 37068 20536 37080
rect 20588 37068 20594 37120
rect 20806 37068 20812 37120
rect 20864 37108 20870 37120
rect 20993 37111 21051 37117
rect 20993 37108 21005 37111
rect 20864 37080 21005 37108
rect 20864 37068 20870 37080
rect 20993 37077 21005 37080
rect 21039 37077 21051 37111
rect 20993 37071 21051 37077
rect 22186 37068 22192 37120
rect 22244 37108 22250 37120
rect 22465 37111 22523 37117
rect 22465 37108 22477 37111
rect 22244 37080 22477 37108
rect 22244 37068 22250 37080
rect 22465 37077 22477 37080
rect 22511 37077 22523 37111
rect 22465 37071 22523 37077
rect 22830 37068 22836 37120
rect 22888 37108 22894 37120
rect 23017 37111 23075 37117
rect 23017 37108 23029 37111
rect 22888 37080 23029 37108
rect 22888 37068 22894 37080
rect 23017 37077 23029 37080
rect 23063 37077 23075 37111
rect 23017 37071 23075 37077
rect 23750 37068 23756 37120
rect 23808 37108 23814 37120
rect 24397 37111 24455 37117
rect 24397 37108 24409 37111
rect 23808 37080 24409 37108
rect 23808 37068 23814 37080
rect 24397 37077 24409 37080
rect 24443 37077 24455 37111
rect 24397 37071 24455 37077
rect 24762 37068 24768 37120
rect 24820 37108 24826 37120
rect 25041 37111 25099 37117
rect 25041 37108 25053 37111
rect 24820 37080 25053 37108
rect 24820 37068 24826 37080
rect 25041 37077 25053 37080
rect 25087 37077 25099 37111
rect 25041 37071 25099 37077
rect 25314 37068 25320 37120
rect 25372 37108 25378 37120
rect 25685 37111 25743 37117
rect 25685 37108 25697 37111
rect 25372 37080 25697 37108
rect 25372 37068 25378 37080
rect 25685 37077 25697 37080
rect 25731 37077 25743 37111
rect 25685 37071 25743 37077
rect 27157 37111 27215 37117
rect 27157 37077 27169 37111
rect 27203 37108 27215 37111
rect 27338 37108 27344 37120
rect 27203 37080 27344 37108
rect 27203 37077 27215 37080
rect 27157 37071 27215 37077
rect 27338 37068 27344 37080
rect 27396 37068 27402 37120
rect 27522 37068 27528 37120
rect 27580 37108 27586 37120
rect 27617 37111 27675 37117
rect 27617 37108 27629 37111
rect 27580 37080 27629 37108
rect 27580 37068 27586 37080
rect 27617 37077 27629 37080
rect 27663 37077 27675 37111
rect 28258 37108 28264 37120
rect 28219 37080 28264 37108
rect 27617 37071 27675 37077
rect 28258 37068 28264 37080
rect 28316 37068 28322 37120
rect 28718 37068 28724 37120
rect 28776 37108 28782 37120
rect 29549 37111 29607 37117
rect 29549 37108 29561 37111
rect 28776 37080 29561 37108
rect 28776 37068 28782 37080
rect 29549 37077 29561 37080
rect 29595 37077 29607 37111
rect 29549 37071 29607 37077
rect 29638 37068 29644 37120
rect 29696 37108 29702 37120
rect 30193 37111 30251 37117
rect 30193 37108 30205 37111
rect 29696 37080 30205 37108
rect 29696 37068 29702 37080
rect 30193 37077 30205 37080
rect 30239 37077 30251 37111
rect 30193 37071 30251 37077
rect 30374 37068 30380 37120
rect 30432 37108 30438 37120
rect 30837 37111 30895 37117
rect 30837 37108 30849 37111
rect 30432 37080 30849 37108
rect 30432 37068 30438 37080
rect 30837 37077 30849 37080
rect 30883 37077 30895 37111
rect 32122 37108 32128 37120
rect 32083 37080 32128 37108
rect 30837 37071 30895 37077
rect 32122 37068 32128 37080
rect 32180 37068 32186 37120
rect 32582 37068 32588 37120
rect 32640 37108 32646 37120
rect 32769 37111 32827 37117
rect 32769 37108 32781 37111
rect 32640 37080 32781 37108
rect 32640 37068 32646 37080
rect 32769 37077 32781 37080
rect 32815 37077 32827 37111
rect 33410 37108 33416 37120
rect 33371 37080 33416 37108
rect 32769 37071 32827 37077
rect 33410 37068 33416 37080
rect 33468 37068 33474 37120
rect 33778 37068 33784 37120
rect 33836 37108 33842 37120
rect 34701 37111 34759 37117
rect 34701 37108 34713 37111
rect 33836 37080 34713 37108
rect 33836 37068 33842 37080
rect 34701 37077 34713 37080
rect 34747 37077 34759 37111
rect 34701 37071 34759 37077
rect 34790 37068 34796 37120
rect 34848 37108 34854 37120
rect 35345 37111 35403 37117
rect 35345 37108 35357 37111
rect 34848 37080 35357 37108
rect 34848 37068 34854 37080
rect 35345 37077 35357 37080
rect 35391 37077 35403 37111
rect 35345 37071 35403 37077
rect 35526 37068 35532 37120
rect 35584 37108 35590 37120
rect 35989 37111 36047 37117
rect 35989 37108 36001 37111
rect 35584 37080 36001 37108
rect 35584 37068 35590 37080
rect 35989 37077 36001 37080
rect 36035 37077 36047 37111
rect 38010 37108 38016 37120
rect 37971 37080 38016 37108
rect 35989 37071 36047 37077
rect 38010 37068 38016 37080
rect 38068 37068 38074 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 14826 36864 14832 36916
rect 14884 36904 14890 36916
rect 14921 36907 14979 36913
rect 14921 36904 14933 36907
rect 14884 36876 14933 36904
rect 14884 36864 14890 36876
rect 14921 36873 14933 36876
rect 14967 36873 14979 36907
rect 15562 36904 15568 36916
rect 15523 36876 15568 36904
rect 14921 36867 14979 36873
rect 15562 36864 15568 36876
rect 15620 36864 15626 36916
rect 16117 36907 16175 36913
rect 16117 36873 16129 36907
rect 16163 36904 16175 36907
rect 16298 36904 16304 36916
rect 16163 36876 16304 36904
rect 16163 36873 16175 36876
rect 16117 36867 16175 36873
rect 16298 36864 16304 36876
rect 16356 36864 16362 36916
rect 17034 36904 17040 36916
rect 16995 36876 17040 36904
rect 17034 36864 17040 36876
rect 17092 36864 17098 36916
rect 17770 36904 17776 36916
rect 17731 36876 17776 36904
rect 17770 36864 17776 36876
rect 17828 36864 17834 36916
rect 18506 36864 18512 36916
rect 18564 36904 18570 36916
rect 18601 36907 18659 36913
rect 18601 36904 18613 36907
rect 18564 36876 18613 36904
rect 18564 36864 18570 36876
rect 18601 36873 18613 36876
rect 18647 36873 18659 36907
rect 19242 36904 19248 36916
rect 19203 36876 19248 36904
rect 18601 36867 18659 36873
rect 19242 36864 19248 36876
rect 19300 36864 19306 36916
rect 19978 36904 19984 36916
rect 19939 36876 19984 36904
rect 19978 36864 19984 36876
rect 20036 36864 20042 36916
rect 20714 36904 20720 36916
rect 20675 36876 20720 36904
rect 20714 36864 20720 36876
rect 20772 36864 20778 36916
rect 23658 36864 23664 36916
rect 23716 36904 23722 36916
rect 24213 36907 24271 36913
rect 24213 36904 24225 36907
rect 23716 36876 24225 36904
rect 23716 36864 23722 36876
rect 24213 36873 24225 36876
rect 24259 36904 24271 36907
rect 24578 36904 24584 36916
rect 24259 36876 24584 36904
rect 24259 36873 24271 36876
rect 24213 36867 24271 36873
rect 24578 36864 24584 36876
rect 24636 36864 24642 36916
rect 24854 36904 24860 36916
rect 24815 36876 24860 36904
rect 24854 36864 24860 36876
rect 24912 36864 24918 36916
rect 25501 36907 25559 36913
rect 25501 36873 25513 36907
rect 25547 36904 25559 36907
rect 25866 36904 25872 36916
rect 25547 36876 25872 36904
rect 25547 36873 25559 36876
rect 25501 36867 25559 36873
rect 25866 36864 25872 36876
rect 25924 36864 25930 36916
rect 26970 36904 26976 36916
rect 26931 36876 26976 36904
rect 26970 36864 26976 36876
rect 27028 36864 27034 36916
rect 27614 36904 27620 36916
rect 27575 36876 27620 36904
rect 27614 36864 27620 36876
rect 27672 36864 27678 36916
rect 29546 36864 29552 36916
rect 29604 36904 29610 36916
rect 30006 36904 30012 36916
rect 29604 36876 30012 36904
rect 29604 36864 29610 36876
rect 30006 36864 30012 36876
rect 30064 36864 30070 36916
rect 30653 36907 30711 36913
rect 30653 36873 30665 36907
rect 30699 36904 30711 36907
rect 31018 36904 31024 36916
rect 30699 36876 31024 36904
rect 30699 36873 30711 36876
rect 30653 36867 30711 36873
rect 31018 36864 31024 36876
rect 31076 36864 31082 36916
rect 32214 36904 32220 36916
rect 32175 36876 32220 36904
rect 32214 36864 32220 36876
rect 32272 36864 32278 36916
rect 32490 36864 32496 36916
rect 32548 36904 32554 36916
rect 32677 36907 32735 36913
rect 32677 36904 32689 36907
rect 32548 36876 32689 36904
rect 32548 36864 32554 36876
rect 32677 36873 32689 36876
rect 32723 36873 32735 36907
rect 34514 36904 34520 36916
rect 34475 36876 34520 36904
rect 32677 36867 32735 36873
rect 34514 36864 34520 36876
rect 34572 36864 34578 36916
rect 36262 36904 36268 36916
rect 36223 36876 36268 36904
rect 36262 36864 36268 36876
rect 36320 36864 36326 36916
rect 36906 36864 36912 36916
rect 36964 36904 36970 36916
rect 37277 36907 37335 36913
rect 37277 36904 37289 36907
rect 36964 36876 37289 36904
rect 36964 36864 36970 36876
rect 37277 36873 37289 36876
rect 37323 36873 37335 36907
rect 37277 36867 37335 36873
rect 2685 36771 2743 36777
rect 2685 36737 2697 36771
rect 2731 36768 2743 36771
rect 3050 36768 3056 36780
rect 2731 36740 3056 36768
rect 2731 36737 2743 36740
rect 2685 36731 2743 36737
rect 3050 36728 3056 36740
rect 3108 36768 3114 36780
rect 3145 36771 3203 36777
rect 3145 36768 3157 36771
rect 3108 36740 3157 36768
rect 3108 36728 3114 36740
rect 3145 36737 3157 36740
rect 3191 36737 3203 36771
rect 4614 36768 4620 36780
rect 4575 36740 4620 36768
rect 3145 36731 3203 36737
rect 4614 36728 4620 36740
rect 4672 36728 4678 36780
rect 6730 36728 6736 36780
rect 6788 36768 6794 36780
rect 6825 36771 6883 36777
rect 6825 36768 6837 36771
rect 6788 36740 6837 36768
rect 6788 36728 6794 36740
rect 6825 36737 6837 36740
rect 6871 36737 6883 36771
rect 6825 36731 6883 36737
rect 8202 36728 8208 36780
rect 8260 36768 8266 36780
rect 8297 36771 8355 36777
rect 8297 36768 8309 36771
rect 8260 36740 8309 36768
rect 8260 36728 8266 36740
rect 8297 36737 8309 36740
rect 8343 36737 8355 36771
rect 8297 36731 8355 36737
rect 9674 36728 9680 36780
rect 9732 36768 9738 36780
rect 9769 36771 9827 36777
rect 9769 36768 9781 36771
rect 9732 36740 9781 36768
rect 9732 36728 9738 36740
rect 9769 36737 9781 36740
rect 9815 36737 9827 36771
rect 9769 36731 9827 36737
rect 11146 36728 11152 36780
rect 11204 36768 11210 36780
rect 11517 36771 11575 36777
rect 11517 36768 11529 36771
rect 11204 36740 11529 36768
rect 11204 36728 11210 36740
rect 11517 36737 11529 36740
rect 11563 36737 11575 36771
rect 11517 36731 11575 36737
rect 12618 36728 12624 36780
rect 12676 36768 12682 36780
rect 12805 36771 12863 36777
rect 12805 36768 12817 36771
rect 12676 36740 12817 36768
rect 12676 36728 12682 36740
rect 12805 36737 12817 36740
rect 12851 36737 12863 36771
rect 12805 36731 12863 36737
rect 13725 36771 13783 36777
rect 13725 36737 13737 36771
rect 13771 36768 13783 36771
rect 14090 36768 14096 36780
rect 13771 36740 14096 36768
rect 13771 36737 13783 36740
rect 13725 36731 13783 36737
rect 14090 36728 14096 36740
rect 14148 36768 14154 36780
rect 14185 36771 14243 36777
rect 14185 36768 14197 36771
rect 14148 36740 14197 36768
rect 14148 36728 14154 36740
rect 14185 36737 14197 36740
rect 14231 36737 14243 36771
rect 14185 36731 14243 36737
rect 21450 36728 21456 36780
rect 21508 36768 21514 36780
rect 21821 36771 21879 36777
rect 21821 36768 21833 36771
rect 21508 36740 21833 36768
rect 21508 36728 21514 36740
rect 21821 36737 21833 36740
rect 21867 36768 21879 36771
rect 22465 36771 22523 36777
rect 22465 36768 22477 36771
rect 21867 36740 22477 36768
rect 21867 36737 21879 36740
rect 21821 36731 21879 36737
rect 22465 36737 22477 36740
rect 22511 36737 22523 36771
rect 25884 36768 25912 36864
rect 26145 36771 26203 36777
rect 26145 36768 26157 36771
rect 25884 36740 26157 36768
rect 22465 36731 22523 36737
rect 26145 36737 26157 36740
rect 26191 36737 26203 36771
rect 31036 36768 31064 36864
rect 36924 36836 36952 36864
rect 35636 36808 36952 36836
rect 35636 36777 35664 36808
rect 31297 36771 31355 36777
rect 31297 36768 31309 36771
rect 31036 36740 31309 36768
rect 26145 36731 26203 36737
rect 31297 36737 31309 36740
rect 31343 36737 31355 36771
rect 31297 36731 31355 36737
rect 34977 36771 35035 36777
rect 34977 36737 34989 36771
rect 35023 36737 35035 36771
rect 34977 36731 35035 36737
rect 35621 36771 35679 36777
rect 35621 36737 35633 36771
rect 35667 36737 35679 36771
rect 35621 36731 35679 36737
rect 3418 36700 3424 36712
rect 3379 36672 3424 36700
rect 3418 36660 3424 36672
rect 3476 36660 3482 36712
rect 4890 36700 4896 36712
rect 4851 36672 4896 36700
rect 4890 36660 4896 36672
rect 4948 36660 4954 36712
rect 7098 36700 7104 36712
rect 7059 36672 7104 36700
rect 7098 36660 7104 36672
rect 7156 36660 7162 36712
rect 8573 36703 8631 36709
rect 8573 36669 8585 36703
rect 8619 36700 8631 36703
rect 8846 36700 8852 36712
rect 8619 36672 8852 36700
rect 8619 36669 8631 36672
rect 8573 36663 8631 36669
rect 8846 36660 8852 36672
rect 8904 36660 8910 36712
rect 10042 36700 10048 36712
rect 10003 36672 10048 36700
rect 10042 36660 10048 36672
rect 10100 36660 10106 36712
rect 11793 36703 11851 36709
rect 11793 36669 11805 36703
rect 11839 36700 11851 36703
rect 11974 36700 11980 36712
rect 11839 36672 11980 36700
rect 11839 36669 11851 36672
rect 11793 36663 11851 36669
rect 11974 36660 11980 36672
rect 12032 36660 12038 36712
rect 34992 36700 35020 36731
rect 36170 36728 36176 36780
rect 36228 36768 36234 36780
rect 36449 36771 36507 36777
rect 36449 36768 36461 36771
rect 36228 36740 36461 36768
rect 36228 36728 36234 36740
rect 36449 36737 36461 36740
rect 36495 36737 36507 36771
rect 36449 36731 36507 36737
rect 36538 36728 36544 36780
rect 36596 36768 36602 36780
rect 37829 36771 37887 36777
rect 37829 36768 37841 36771
rect 36596 36740 37841 36768
rect 36596 36728 36602 36740
rect 37829 36737 37841 36740
rect 37875 36737 37887 36771
rect 37829 36731 37887 36737
rect 35342 36700 35348 36712
rect 34992 36672 35348 36700
rect 35342 36660 35348 36672
rect 35400 36700 35406 36712
rect 37642 36700 37648 36712
rect 35400 36672 37648 36700
rect 35400 36660 35406 36672
rect 37642 36660 37648 36672
rect 37700 36660 37706 36712
rect 35805 36635 35863 36641
rect 35805 36601 35817 36635
rect 35851 36632 35863 36635
rect 36354 36632 36360 36644
rect 35851 36604 36360 36632
rect 35851 36601 35863 36604
rect 35805 36595 35863 36601
rect 36354 36592 36360 36604
rect 36412 36592 36418 36644
rect 37182 36592 37188 36644
rect 37240 36632 37246 36644
rect 38013 36635 38071 36641
rect 38013 36632 38025 36635
rect 37240 36604 38025 36632
rect 37240 36592 37246 36604
rect 38013 36601 38025 36604
rect 38059 36601 38071 36635
rect 38013 36595 38071 36601
rect 12986 36564 12992 36576
rect 12947 36536 12992 36564
rect 12986 36524 12992 36536
rect 13044 36524 13050 36576
rect 14369 36567 14427 36573
rect 14369 36533 14381 36567
rect 14415 36564 14427 36567
rect 14826 36564 14832 36576
rect 14415 36536 14832 36564
rect 14415 36533 14427 36536
rect 14369 36527 14427 36533
rect 14826 36524 14832 36536
rect 14884 36524 14890 36576
rect 22005 36567 22063 36573
rect 22005 36533 22017 36567
rect 22051 36564 22063 36567
rect 22186 36564 22192 36576
rect 22051 36536 22192 36564
rect 22051 36533 22063 36536
rect 22005 36527 22063 36533
rect 22186 36524 22192 36536
rect 22244 36524 22250 36576
rect 25774 36524 25780 36576
rect 25832 36564 25838 36576
rect 25961 36567 26019 36573
rect 25961 36564 25973 36567
rect 25832 36536 25973 36564
rect 25832 36524 25838 36536
rect 25961 36533 25973 36536
rect 26007 36533 26019 36567
rect 29362 36564 29368 36576
rect 29323 36536 29368 36564
rect 25961 36527 26019 36533
rect 29362 36524 29368 36536
rect 29420 36524 29426 36576
rect 31110 36564 31116 36576
rect 31071 36536 31116 36564
rect 31110 36524 31116 36536
rect 31168 36524 31174 36576
rect 35161 36567 35219 36573
rect 35161 36533 35173 36567
rect 35207 36564 35219 36567
rect 37458 36564 37464 36576
rect 35207 36536 37464 36564
rect 35207 36533 35219 36536
rect 35161 36527 35219 36533
rect 37458 36524 37464 36536
rect 37516 36524 37522 36576
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 4525 36363 4583 36369
rect 4525 36329 4537 36363
rect 4571 36360 4583 36363
rect 4614 36360 4620 36372
rect 4571 36332 4620 36360
rect 4571 36329 4583 36332
rect 4525 36323 4583 36329
rect 4614 36320 4620 36332
rect 4672 36320 4678 36372
rect 4706 36320 4712 36372
rect 4764 36360 4770 36372
rect 4982 36360 4988 36372
rect 4764 36332 4988 36360
rect 4764 36320 4770 36332
rect 4982 36320 4988 36332
rect 5040 36320 5046 36372
rect 6730 36320 6736 36372
rect 6788 36360 6794 36372
rect 7377 36363 7435 36369
rect 7377 36360 7389 36363
rect 6788 36332 7389 36360
rect 6788 36320 6794 36332
rect 7377 36329 7389 36332
rect 7423 36329 7435 36363
rect 8202 36360 8208 36372
rect 8163 36332 8208 36360
rect 7377 36323 7435 36329
rect 8202 36320 8208 36332
rect 8260 36320 8266 36372
rect 9674 36320 9680 36372
rect 9732 36360 9738 36372
rect 10321 36363 10379 36369
rect 10321 36360 10333 36363
rect 9732 36332 10333 36360
rect 9732 36320 9738 36332
rect 10321 36329 10333 36332
rect 10367 36329 10379 36363
rect 10321 36323 10379 36329
rect 11146 36320 11152 36372
rect 11204 36360 11210 36372
rect 11333 36363 11391 36369
rect 11333 36360 11345 36363
rect 11204 36332 11345 36360
rect 11204 36320 11210 36332
rect 11333 36329 11345 36332
rect 11379 36329 11391 36363
rect 11882 36360 11888 36372
rect 11843 36332 11888 36360
rect 11333 36323 11391 36329
rect 11882 36320 11888 36332
rect 11940 36320 11946 36372
rect 12618 36360 12624 36372
rect 12579 36332 12624 36360
rect 12618 36320 12624 36332
rect 12676 36320 12682 36372
rect 35342 36360 35348 36372
rect 35303 36332 35348 36360
rect 35342 36320 35348 36332
rect 35400 36320 35406 36372
rect 5629 36227 5687 36233
rect 5629 36193 5641 36227
rect 5675 36224 5687 36227
rect 5994 36224 6000 36236
rect 5675 36196 6000 36224
rect 5675 36193 5687 36196
rect 5629 36187 5687 36193
rect 5994 36184 6000 36196
rect 6052 36224 6058 36236
rect 6089 36227 6147 36233
rect 6089 36224 6101 36227
rect 6052 36196 6101 36224
rect 6052 36184 6058 36196
rect 6089 36193 6101 36196
rect 6135 36193 6147 36227
rect 6089 36187 6147 36193
rect 8938 36184 8944 36236
rect 8996 36224 9002 36236
rect 9033 36227 9091 36233
rect 9033 36224 9045 36227
rect 8996 36196 9045 36224
rect 8996 36184 9002 36196
rect 9033 36193 9045 36196
rect 9079 36193 9091 36227
rect 9033 36187 9091 36193
rect 34793 36227 34851 36233
rect 34793 36193 34805 36227
rect 34839 36224 34851 36227
rect 38102 36224 38108 36236
rect 34839 36196 38108 36224
rect 34839 36193 34851 36196
rect 34793 36187 34851 36193
rect 38102 36184 38108 36196
rect 38160 36184 38166 36236
rect 6362 36156 6368 36168
rect 6323 36128 6368 36156
rect 6362 36116 6368 36128
rect 6420 36116 6426 36168
rect 9214 36116 9220 36168
rect 9272 36156 9278 36168
rect 9309 36159 9367 36165
rect 9309 36156 9321 36159
rect 9272 36128 9321 36156
rect 9272 36116 9278 36128
rect 9309 36125 9321 36128
rect 9355 36125 9367 36159
rect 9309 36119 9367 36125
rect 35805 36159 35863 36165
rect 35805 36125 35817 36159
rect 35851 36156 35863 36159
rect 36170 36156 36176 36168
rect 35851 36128 36176 36156
rect 35851 36125 35863 36128
rect 35805 36119 35863 36125
rect 36170 36116 36176 36128
rect 36228 36116 36234 36168
rect 37826 36156 37832 36168
rect 37787 36128 37832 36156
rect 37826 36116 37832 36128
rect 37884 36116 37890 36168
rect 36446 36088 36452 36100
rect 36407 36060 36452 36088
rect 36446 36048 36452 36060
rect 36504 36048 36510 36100
rect 35986 36020 35992 36032
rect 35947 35992 35992 36020
rect 35986 35980 35992 35992
rect 36044 35980 36050 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 8938 35816 8944 35828
rect 8899 35788 8944 35816
rect 8938 35776 8944 35788
rect 8996 35776 9002 35828
rect 28810 35776 28816 35828
rect 28868 35816 28874 35828
rect 29362 35816 29368 35828
rect 28868 35788 29368 35816
rect 28868 35776 28874 35788
rect 29362 35776 29368 35788
rect 29420 35776 29426 35828
rect 35621 35819 35679 35825
rect 35621 35785 35633 35819
rect 35667 35816 35679 35819
rect 35802 35816 35808 35828
rect 35667 35788 35808 35816
rect 35667 35785 35679 35788
rect 35621 35779 35679 35785
rect 35802 35776 35808 35788
rect 35860 35776 35866 35828
rect 36170 35816 36176 35828
rect 36131 35788 36176 35816
rect 36170 35776 36176 35788
rect 36228 35776 36234 35828
rect 36722 35640 36728 35692
rect 36780 35680 36786 35692
rect 37829 35683 37887 35689
rect 37829 35680 37841 35683
rect 36780 35652 37841 35680
rect 36780 35640 36786 35652
rect 37829 35649 37841 35652
rect 37875 35649 37887 35683
rect 37829 35643 37887 35649
rect 36633 35615 36691 35621
rect 36633 35581 36645 35615
rect 36679 35612 36691 35615
rect 37642 35612 37648 35624
rect 36679 35584 37648 35612
rect 36679 35581 36691 35584
rect 36633 35575 36691 35581
rect 37642 35572 37648 35584
rect 37700 35572 37706 35624
rect 37090 35504 37096 35556
rect 37148 35544 37154 35556
rect 38013 35547 38071 35553
rect 38013 35544 38025 35547
rect 37148 35516 38025 35544
rect 37148 35504 37154 35516
rect 38013 35513 38025 35516
rect 38059 35513 38071 35547
rect 38013 35507 38071 35513
rect 35069 35479 35127 35485
rect 35069 35445 35081 35479
rect 35115 35476 35127 35479
rect 35894 35476 35900 35488
rect 35115 35448 35900 35476
rect 35115 35445 35127 35448
rect 35069 35439 35127 35445
rect 35894 35436 35900 35448
rect 35952 35476 35958 35488
rect 36446 35476 36452 35488
rect 35952 35448 36452 35476
rect 35952 35436 35958 35448
rect 36446 35436 36452 35448
rect 36504 35476 36510 35488
rect 37277 35479 37335 35485
rect 37277 35476 37289 35479
rect 36504 35448 37289 35476
rect 36504 35436 36510 35448
rect 37277 35445 37289 35448
rect 37323 35445 37335 35479
rect 37277 35439 37335 35445
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 36814 35068 36820 35080
rect 36775 35040 36820 35068
rect 36814 35028 36820 35040
rect 36872 35028 36878 35080
rect 37734 35068 37740 35080
rect 37695 35040 37740 35068
rect 37734 35028 37740 35040
rect 37792 35028 37798 35080
rect 37918 35068 37924 35080
rect 37879 35040 37924 35068
rect 37918 35028 37924 35040
rect 37976 35028 37982 35080
rect 38010 35000 38016 35012
rect 35728 34972 38016 35000
rect 35434 34892 35440 34944
rect 35492 34932 35498 34944
rect 35728 34941 35756 34972
rect 38010 34960 38016 34972
rect 38068 34960 38074 35012
rect 35713 34935 35771 34941
rect 35713 34932 35725 34935
rect 35492 34904 35725 34932
rect 35492 34892 35498 34904
rect 35713 34901 35725 34904
rect 35759 34901 35771 34935
rect 35713 34895 35771 34901
rect 35894 34892 35900 34944
rect 35952 34932 35958 34944
rect 36265 34935 36323 34941
rect 36265 34932 36277 34935
rect 35952 34904 36277 34932
rect 35952 34892 35958 34904
rect 36265 34901 36277 34904
rect 36311 34901 36323 34935
rect 36998 34932 37004 34944
rect 36959 34904 37004 34932
rect 36265 34895 36323 34901
rect 36998 34892 37004 34904
rect 37056 34892 37062 34944
rect 37550 34932 37556 34944
rect 37511 34904 37556 34932
rect 37550 34892 37556 34904
rect 37608 34892 37614 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 35434 34728 35440 34740
rect 35395 34700 35440 34728
rect 35434 34688 35440 34700
rect 35492 34688 35498 34740
rect 36081 34731 36139 34737
rect 36081 34697 36093 34731
rect 36127 34728 36139 34731
rect 36538 34728 36544 34740
rect 36127 34700 36544 34728
rect 36127 34697 36139 34700
rect 36081 34691 36139 34697
rect 36538 34688 36544 34700
rect 36596 34688 36602 34740
rect 37461 34731 37519 34737
rect 37461 34697 37473 34731
rect 37507 34728 37519 34731
rect 37826 34728 37832 34740
rect 37507 34700 37832 34728
rect 37507 34697 37519 34700
rect 37461 34691 37519 34697
rect 37826 34688 37832 34700
rect 37884 34688 37890 34740
rect 37550 34660 37556 34672
rect 35912 34632 37556 34660
rect 35912 34601 35940 34632
rect 37550 34620 37556 34632
rect 37608 34620 37614 34672
rect 38010 34660 38016 34672
rect 37844 34632 38016 34660
rect 35897 34595 35955 34601
rect 35897 34561 35909 34595
rect 35943 34561 35955 34595
rect 35897 34555 35955 34561
rect 35986 34552 35992 34604
rect 36044 34592 36050 34604
rect 36541 34595 36599 34601
rect 36541 34592 36553 34595
rect 36044 34564 36553 34592
rect 36044 34552 36050 34564
rect 36541 34561 36553 34564
rect 36587 34561 36599 34595
rect 36541 34555 36599 34561
rect 37642 34552 37648 34604
rect 37700 34592 37706 34604
rect 37844 34601 37872 34632
rect 38010 34620 38016 34632
rect 38068 34620 38074 34672
rect 37737 34595 37795 34601
rect 37737 34592 37749 34595
rect 37700 34564 37749 34592
rect 37700 34552 37706 34564
rect 37737 34561 37749 34564
rect 37783 34561 37795 34595
rect 37737 34555 37795 34561
rect 37829 34595 37887 34601
rect 37829 34561 37841 34595
rect 37875 34561 37887 34595
rect 37829 34555 37887 34561
rect 37918 34552 37924 34604
rect 37976 34592 37982 34604
rect 38105 34595 38163 34601
rect 37976 34564 38069 34592
rect 37976 34552 37982 34564
rect 38105 34561 38117 34595
rect 38151 34592 38163 34595
rect 38194 34592 38200 34604
rect 38151 34564 38200 34592
rect 38151 34561 38163 34564
rect 38105 34555 38163 34561
rect 38194 34552 38200 34564
rect 38252 34552 38258 34604
rect 36633 34527 36691 34533
rect 36633 34493 36645 34527
rect 36679 34524 36691 34527
rect 37936 34524 37964 34552
rect 36679 34496 37964 34524
rect 36679 34493 36691 34496
rect 36633 34487 36691 34493
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 37734 34144 37740 34196
rect 37792 34184 37798 34196
rect 37829 34187 37887 34193
rect 37829 34184 37841 34187
rect 37792 34156 37841 34184
rect 37792 34144 37798 34156
rect 37829 34153 37841 34156
rect 37875 34153 37887 34187
rect 37829 34147 37887 34153
rect 35894 34008 35900 34060
rect 35952 34048 35958 34060
rect 35989 34051 36047 34057
rect 35989 34048 36001 34051
rect 35952 34020 36001 34048
rect 35952 34008 35958 34020
rect 35989 34017 36001 34020
rect 36035 34048 36047 34051
rect 37185 34051 37243 34057
rect 37185 34048 37197 34051
rect 36035 34020 37197 34048
rect 36035 34017 36047 34020
rect 35989 34011 36047 34017
rect 37185 34017 37197 34020
rect 37231 34017 37243 34051
rect 37185 34011 37243 34017
rect 37369 34051 37427 34057
rect 37369 34017 37381 34051
rect 37415 34048 37427 34051
rect 38010 34048 38016 34060
rect 37415 34020 38016 34048
rect 37415 34017 37427 34020
rect 37369 34011 37427 34017
rect 38010 34008 38016 34020
rect 38068 34008 38074 34060
rect 36262 33980 36268 33992
rect 36223 33952 36268 33980
rect 36262 33940 36268 33952
rect 36320 33940 36326 33992
rect 37458 33980 37464 33992
rect 37419 33952 37464 33980
rect 37458 33940 37464 33952
rect 37516 33940 37522 33992
rect 35437 33847 35495 33853
rect 35437 33813 35449 33847
rect 35483 33844 35495 33847
rect 36173 33847 36231 33853
rect 36173 33844 36185 33847
rect 35483 33816 36185 33844
rect 35483 33813 35495 33816
rect 35437 33807 35495 33813
rect 36173 33813 36185 33816
rect 36219 33844 36231 33847
rect 36446 33844 36452 33856
rect 36219 33816 36452 33844
rect 36219 33813 36231 33816
rect 36173 33807 36231 33813
rect 36446 33804 36452 33816
rect 36504 33804 36510 33856
rect 36538 33804 36544 33856
rect 36596 33844 36602 33856
rect 36633 33847 36691 33853
rect 36633 33844 36645 33847
rect 36596 33816 36645 33844
rect 36596 33804 36602 33816
rect 36633 33813 36645 33816
rect 36679 33813 36691 33847
rect 36633 33807 36691 33813
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 36722 33640 36728 33652
rect 36683 33612 36728 33640
rect 36722 33600 36728 33612
rect 36780 33600 36786 33652
rect 37277 33643 37335 33649
rect 37277 33609 37289 33643
rect 37323 33640 37335 33643
rect 37458 33640 37464 33652
rect 37323 33612 37464 33640
rect 37323 33609 37335 33612
rect 37277 33603 37335 33609
rect 37458 33600 37464 33612
rect 37516 33600 37522 33652
rect 37921 33643 37979 33649
rect 37921 33609 37933 33643
rect 37967 33640 37979 33643
rect 38194 33640 38200 33652
rect 37967 33612 38200 33640
rect 37967 33609 37979 33612
rect 37921 33603 37979 33609
rect 38194 33600 38200 33612
rect 38252 33600 38258 33652
rect 36538 33504 36544 33516
rect 36499 33476 36544 33504
rect 36538 33464 36544 33476
rect 36596 33464 36602 33516
rect 37737 33507 37795 33513
rect 37737 33473 37749 33507
rect 37783 33504 37795 33507
rect 38010 33504 38016 33516
rect 37783 33476 38016 33504
rect 37783 33473 37795 33476
rect 37737 33467 37795 33473
rect 38010 33464 38016 33476
rect 38068 33464 38074 33516
rect 37642 33436 37648 33448
rect 37603 33408 37648 33436
rect 37642 33396 37648 33408
rect 37700 33396 37706 33448
rect 34514 33260 34520 33312
rect 34572 33300 34578 33312
rect 34977 33303 35035 33309
rect 34977 33300 34989 33303
rect 34572 33272 34989 33300
rect 34572 33260 34578 33272
rect 34977 33269 34989 33272
rect 35023 33269 35035 33303
rect 35986 33300 35992 33312
rect 35947 33272 35992 33300
rect 34977 33263 35035 33269
rect 35986 33260 35992 33272
rect 36044 33260 36050 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 37274 33096 37280 33108
rect 37235 33068 37280 33096
rect 37274 33056 37280 33068
rect 37332 33056 37338 33108
rect 35897 33031 35955 33037
rect 35897 32997 35909 33031
rect 35943 32997 35955 33031
rect 35897 32991 35955 32997
rect 36541 33031 36599 33037
rect 36541 32997 36553 33031
rect 36587 32997 36599 33031
rect 36541 32991 36599 32997
rect 34514 32920 34520 32972
rect 34572 32960 34578 32972
rect 35253 32963 35311 32969
rect 35253 32960 35265 32963
rect 34572 32932 35265 32960
rect 34572 32920 34578 32932
rect 35253 32929 35265 32932
rect 35299 32929 35311 32963
rect 35253 32923 35311 32929
rect 35526 32892 35532 32904
rect 35487 32864 35532 32892
rect 35526 32852 35532 32864
rect 35584 32852 35590 32904
rect 35912 32892 35940 32991
rect 36357 32895 36415 32901
rect 36357 32892 36369 32895
rect 35912 32864 36369 32892
rect 36357 32861 36369 32864
rect 36403 32861 36415 32895
rect 36556 32892 36584 32991
rect 37093 32895 37151 32901
rect 37093 32892 37105 32895
rect 36556 32864 37105 32892
rect 36357 32855 36415 32861
rect 37093 32861 37105 32864
rect 37139 32861 37151 32895
rect 37826 32892 37832 32904
rect 37787 32864 37832 32892
rect 37093 32855 37151 32861
rect 37826 32852 37832 32864
rect 37884 32852 37890 32904
rect 35434 32824 35440 32836
rect 35347 32796 35440 32824
rect 35434 32784 35440 32796
rect 35492 32824 35498 32836
rect 35986 32824 35992 32836
rect 35492 32796 35992 32824
rect 35492 32784 35498 32796
rect 35986 32784 35992 32796
rect 36044 32784 36050 32836
rect 38010 32756 38016 32768
rect 37971 32728 38016 32756
rect 38010 32716 38016 32728
rect 38068 32716 38074 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 34790 32552 34796 32564
rect 34751 32524 34796 32552
rect 34790 32512 34796 32524
rect 34848 32512 34854 32564
rect 35161 32555 35219 32561
rect 35161 32521 35173 32555
rect 35207 32521 35219 32555
rect 35161 32515 35219 32521
rect 35805 32555 35863 32561
rect 35805 32521 35817 32555
rect 35851 32552 35863 32555
rect 37826 32552 37832 32564
rect 35851 32524 37832 32552
rect 35851 32521 35863 32524
rect 35805 32515 35863 32521
rect 35176 32416 35204 32515
rect 37826 32512 37832 32524
rect 37884 32512 37890 32564
rect 35621 32419 35679 32425
rect 35621 32416 35633 32419
rect 35176 32388 35633 32416
rect 35621 32385 35633 32388
rect 35667 32385 35679 32419
rect 37826 32416 37832 32428
rect 37787 32388 37832 32416
rect 35621 32379 35679 32385
rect 37826 32376 37832 32388
rect 37884 32376 37890 32428
rect 34514 32348 34520 32360
rect 33888 32320 34520 32348
rect 31662 32172 31668 32224
rect 31720 32212 31726 32224
rect 33888 32221 33916 32320
rect 34514 32308 34520 32320
rect 34572 32308 34578 32360
rect 34698 32348 34704 32360
rect 34659 32320 34704 32348
rect 34698 32308 34704 32320
rect 34756 32308 34762 32360
rect 34532 32280 34560 32308
rect 37277 32283 37335 32289
rect 37277 32280 37289 32283
rect 34532 32252 37289 32280
rect 37277 32249 37289 32252
rect 37323 32280 37335 32283
rect 37642 32280 37648 32292
rect 37323 32252 37648 32280
rect 37323 32249 37335 32252
rect 37277 32243 37335 32249
rect 37642 32240 37648 32252
rect 37700 32240 37706 32292
rect 33873 32215 33931 32221
rect 33873 32212 33885 32215
rect 31720 32184 33885 32212
rect 31720 32172 31726 32184
rect 33873 32181 33885 32184
rect 33919 32181 33931 32215
rect 38010 32212 38016 32224
rect 37971 32184 38016 32212
rect 33873 32175 33931 32181
rect 38010 32172 38016 32184
rect 38068 32172 38074 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 34698 31968 34704 32020
rect 34756 32008 34762 32020
rect 35345 32011 35403 32017
rect 35345 32008 35357 32011
rect 34756 31980 35357 32008
rect 34756 31968 34762 31980
rect 35345 31977 35357 31980
rect 35391 31977 35403 32011
rect 35345 31971 35403 31977
rect 37734 31968 37740 32020
rect 37792 32008 37798 32020
rect 38102 32008 38108 32020
rect 37792 31980 38108 32008
rect 37792 31968 37798 31980
rect 38102 31968 38108 31980
rect 38160 31968 38166 32020
rect 34149 31943 34207 31949
rect 34149 31909 34161 31943
rect 34195 31909 34207 31943
rect 34149 31903 34207 31909
rect 34885 31943 34943 31949
rect 34885 31909 34897 31943
rect 34931 31940 34943 31943
rect 37826 31940 37832 31952
rect 34931 31912 37832 31940
rect 34931 31909 34943 31912
rect 34885 31903 34943 31909
rect 33594 31872 33600 31884
rect 33555 31844 33600 31872
rect 33594 31832 33600 31844
rect 33652 31832 33658 31884
rect 34164 31804 34192 31903
rect 37826 31900 37832 31912
rect 37884 31900 37890 31952
rect 34701 31807 34759 31813
rect 34701 31804 34713 31807
rect 34164 31776 34713 31804
rect 34701 31773 34713 31776
rect 34747 31773 34759 31807
rect 34701 31767 34759 31773
rect 33778 31736 33784 31748
rect 33739 31708 33784 31736
rect 33778 31696 33784 31708
rect 33836 31696 33842 31748
rect 33689 31671 33747 31677
rect 33689 31637 33701 31671
rect 33735 31668 33747 31671
rect 33962 31668 33968 31680
rect 33735 31640 33968 31668
rect 33735 31637 33747 31640
rect 33689 31631 33747 31637
rect 33962 31628 33968 31640
rect 34020 31628 34026 31680
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 34606 31288 34612 31340
rect 34664 31328 34670 31340
rect 37829 31331 37887 31337
rect 37829 31328 37841 31331
rect 34664 31300 37841 31328
rect 34664 31288 34670 31300
rect 37829 31297 37841 31300
rect 37875 31297 37887 31331
rect 37829 31291 37887 31297
rect 33594 31152 33600 31204
rect 33652 31192 33658 31204
rect 34885 31195 34943 31201
rect 34885 31192 34897 31195
rect 33652 31164 34897 31192
rect 33652 31152 33658 31164
rect 34885 31161 34897 31164
rect 34931 31192 34943 31195
rect 35894 31192 35900 31204
rect 34931 31164 35900 31192
rect 34931 31161 34943 31164
rect 34885 31155 34943 31161
rect 35894 31152 35900 31164
rect 35952 31152 35958 31204
rect 38010 31192 38016 31204
rect 37971 31164 38016 31192
rect 38010 31152 38016 31164
rect 38068 31152 38074 31204
rect 33962 31084 33968 31136
rect 34020 31124 34026 31136
rect 34241 31127 34299 31133
rect 34241 31124 34253 31127
rect 34020 31096 34253 31124
rect 34020 31084 34026 31096
rect 34241 31093 34253 31096
rect 34287 31093 34299 31127
rect 34241 31087 34299 31093
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 34514 30676 34520 30728
rect 34572 30716 34578 30728
rect 37829 30719 37887 30725
rect 37829 30716 37841 30719
rect 34572 30688 37841 30716
rect 34572 30676 34578 30688
rect 37829 30685 37841 30688
rect 37875 30685 37887 30719
rect 37829 30679 37887 30685
rect 32490 30540 32496 30592
rect 32548 30580 32554 30592
rect 33137 30583 33195 30589
rect 33137 30580 33149 30583
rect 32548 30552 33149 30580
rect 32548 30540 32554 30552
rect 33137 30549 33149 30552
rect 33183 30549 33195 30583
rect 38010 30580 38016 30592
rect 37971 30552 38016 30580
rect 33137 30543 33195 30549
rect 38010 30540 38016 30552
rect 38068 30540 38074 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 32582 30308 32588 30320
rect 32543 30280 32588 30308
rect 32582 30268 32588 30280
rect 32640 30268 32646 30320
rect 33413 30243 33471 30249
rect 33413 30240 33425 30243
rect 32968 30212 33425 30240
rect 32306 30172 32312 30184
rect 32267 30144 32312 30172
rect 32306 30132 32312 30144
rect 32364 30132 32370 30184
rect 32490 30172 32496 30184
rect 32451 30144 32496 30172
rect 32490 30132 32496 30144
rect 32548 30132 32554 30184
rect 32968 30113 32996 30212
rect 33413 30209 33425 30212
rect 33459 30209 33471 30243
rect 33413 30203 33471 30209
rect 33502 30200 33508 30252
rect 33560 30240 33566 30252
rect 34057 30243 34115 30249
rect 34057 30240 34069 30243
rect 33560 30212 34069 30240
rect 33560 30200 33566 30212
rect 34057 30209 34069 30212
rect 34103 30209 34115 30243
rect 34057 30203 34115 30209
rect 34146 30200 34152 30252
rect 34204 30240 34210 30252
rect 37829 30243 37887 30249
rect 37829 30240 37841 30243
rect 34204 30212 37841 30240
rect 34204 30200 34210 30212
rect 37829 30209 37841 30212
rect 37875 30209 37887 30243
rect 37829 30203 37887 30209
rect 32953 30107 33011 30113
rect 32953 30073 32965 30107
rect 32999 30073 33011 30107
rect 32953 30067 33011 30073
rect 33597 30107 33655 30113
rect 33597 30073 33609 30107
rect 33643 30104 33655 30107
rect 34514 30104 34520 30116
rect 33643 30076 34520 30104
rect 33643 30073 33655 30076
rect 33597 30067 33655 30073
rect 34514 30064 34520 30076
rect 34572 30064 34578 30116
rect 34241 30039 34299 30045
rect 34241 30005 34253 30039
rect 34287 30036 34299 30039
rect 34606 30036 34612 30048
rect 34287 30008 34612 30036
rect 34287 30005 34299 30008
rect 34241 29999 34299 30005
rect 34606 29996 34612 30008
rect 34664 29996 34670 30048
rect 38010 30036 38016 30048
rect 37971 30008 38016 30036
rect 38010 29996 38016 30008
rect 38068 29996 38074 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 33502 29832 33508 29844
rect 33463 29804 33508 29832
rect 33502 29792 33508 29804
rect 33560 29792 33566 29844
rect 30190 29656 30196 29708
rect 30248 29696 30254 29708
rect 31665 29699 31723 29705
rect 31665 29696 31677 29699
rect 30248 29668 31677 29696
rect 30248 29656 30254 29668
rect 31665 29665 31677 29668
rect 31711 29696 31723 29699
rect 32306 29696 32312 29708
rect 31711 29668 32312 29696
rect 31711 29665 31723 29668
rect 31665 29659 31723 29665
rect 32306 29656 32312 29668
rect 32364 29696 32370 29708
rect 32861 29699 32919 29705
rect 32861 29696 32873 29699
rect 32364 29668 32873 29696
rect 32364 29656 32370 29668
rect 32861 29665 32873 29668
rect 32907 29665 32919 29699
rect 32861 29659 32919 29665
rect 31941 29631 31999 29637
rect 31941 29597 31953 29631
rect 31987 29628 31999 29631
rect 32122 29628 32128 29640
rect 31987 29600 32128 29628
rect 31987 29597 31999 29600
rect 31941 29591 31999 29597
rect 32122 29588 32128 29600
rect 32180 29588 32186 29640
rect 33137 29631 33195 29637
rect 33137 29597 33149 29631
rect 33183 29628 33195 29631
rect 33410 29628 33416 29640
rect 33183 29600 33416 29628
rect 33183 29597 33195 29600
rect 33137 29591 33195 29597
rect 33410 29588 33416 29600
rect 33468 29588 33474 29640
rect 33502 29588 33508 29640
rect 33560 29628 33566 29640
rect 37829 29631 37887 29637
rect 37829 29628 37841 29631
rect 33560 29600 37841 29628
rect 33560 29588 33566 29600
rect 37829 29597 37841 29600
rect 37875 29597 37887 29631
rect 37829 29591 37887 29597
rect 31849 29563 31907 29569
rect 31849 29529 31861 29563
rect 31895 29560 31907 29563
rect 32398 29560 32404 29572
rect 31895 29532 32404 29560
rect 31895 29529 31907 29532
rect 31849 29523 31907 29529
rect 32398 29520 32404 29532
rect 32456 29560 32462 29572
rect 33965 29563 34023 29569
rect 33965 29560 33977 29563
rect 32456 29532 33977 29560
rect 32456 29520 32462 29532
rect 33965 29529 33977 29532
rect 34011 29529 34023 29563
rect 33965 29523 34023 29529
rect 32309 29495 32367 29501
rect 32309 29461 32321 29495
rect 32355 29492 32367 29495
rect 32766 29492 32772 29504
rect 32355 29464 32772 29492
rect 32355 29461 32367 29464
rect 32309 29455 32367 29461
rect 32766 29452 32772 29464
rect 32824 29452 32830 29504
rect 33045 29495 33103 29501
rect 33045 29461 33057 29495
rect 33091 29492 33103 29495
rect 33594 29492 33600 29504
rect 33091 29464 33600 29492
rect 33091 29461 33103 29464
rect 33045 29455 33103 29461
rect 33594 29452 33600 29464
rect 33652 29452 33658 29504
rect 38010 29492 38016 29504
rect 37971 29464 38016 29492
rect 38010 29452 38016 29464
rect 38068 29452 38074 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 31110 29288 31116 29300
rect 31071 29260 31116 29288
rect 31110 29248 31116 29260
rect 31168 29248 31174 29300
rect 31481 29291 31539 29297
rect 31481 29257 31493 29291
rect 31527 29257 31539 29291
rect 31481 29251 31539 29257
rect 32309 29291 32367 29297
rect 32309 29257 32321 29291
rect 32355 29288 32367 29291
rect 33502 29288 33508 29300
rect 32355 29260 33508 29288
rect 32355 29257 32367 29260
rect 32309 29251 32367 29257
rect 31496 29152 31524 29251
rect 33502 29248 33508 29260
rect 33560 29248 33566 29300
rect 32125 29155 32183 29161
rect 32125 29152 32137 29155
rect 31496 29124 32137 29152
rect 32125 29121 32137 29124
rect 32171 29121 32183 29155
rect 32766 29152 32772 29164
rect 32727 29124 32772 29152
rect 32125 29115 32183 29121
rect 32766 29112 32772 29124
rect 32824 29112 32830 29164
rect 30190 29044 30196 29096
rect 30248 29084 30254 29096
rect 30837 29087 30895 29093
rect 30837 29084 30849 29087
rect 30248 29056 30849 29084
rect 30248 29044 30254 29056
rect 30837 29053 30849 29056
rect 30883 29053 30895 29087
rect 30837 29047 30895 29053
rect 31021 29087 31079 29093
rect 31021 29053 31033 29087
rect 31067 29084 31079 29087
rect 32306 29084 32312 29096
rect 31067 29056 32312 29084
rect 31067 29053 31079 29056
rect 31021 29047 31079 29053
rect 32306 29044 32312 29056
rect 32364 29044 32370 29096
rect 34146 29084 34152 29096
rect 32968 29056 34152 29084
rect 32968 29025 32996 29056
rect 34146 29044 34152 29056
rect 34204 29044 34210 29096
rect 32953 29019 33011 29025
rect 32953 28985 32965 29019
rect 32999 28985 33011 29019
rect 33594 29016 33600 29028
rect 33555 28988 33600 29016
rect 32953 28979 33011 28985
rect 33594 28976 33600 28988
rect 33652 28976 33658 29028
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 31389 28679 31447 28685
rect 31389 28645 31401 28679
rect 31435 28676 31447 28679
rect 31435 28648 35894 28676
rect 31435 28645 31447 28648
rect 31389 28639 31447 28645
rect 30190 28608 30196 28620
rect 30151 28580 30196 28608
rect 30190 28568 30196 28580
rect 30248 28568 30254 28620
rect 30285 28611 30343 28617
rect 30285 28577 30297 28611
rect 30331 28608 30343 28611
rect 30650 28608 30656 28620
rect 30331 28580 30656 28608
rect 30331 28577 30343 28580
rect 30285 28571 30343 28577
rect 30650 28568 30656 28580
rect 30708 28608 30714 28620
rect 31849 28611 31907 28617
rect 31849 28608 31861 28611
rect 30708 28580 31861 28608
rect 30708 28568 30714 28580
rect 31849 28577 31861 28580
rect 31895 28577 31907 28611
rect 31849 28571 31907 28577
rect 30374 28540 30380 28552
rect 30335 28512 30380 28540
rect 30374 28500 30380 28512
rect 30432 28500 30438 28552
rect 31205 28543 31263 28549
rect 31205 28540 31217 28543
rect 30760 28512 31217 28540
rect 30760 28413 30788 28512
rect 31205 28509 31217 28512
rect 31251 28509 31263 28543
rect 35866 28540 35894 28648
rect 37829 28543 37887 28549
rect 37829 28540 37841 28543
rect 35866 28512 37841 28540
rect 31205 28503 31263 28509
rect 37829 28509 37841 28512
rect 37875 28509 37887 28543
rect 37829 28503 37887 28509
rect 30745 28407 30803 28413
rect 30745 28373 30757 28407
rect 30791 28373 30803 28407
rect 30745 28367 30803 28373
rect 32306 28364 32312 28416
rect 32364 28404 32370 28416
rect 32401 28407 32459 28413
rect 32401 28404 32413 28407
rect 32364 28376 32413 28404
rect 32364 28364 32370 28376
rect 32401 28373 32413 28376
rect 32447 28373 32459 28407
rect 38010 28404 38016 28416
rect 37971 28376 38016 28404
rect 32401 28367 32459 28373
rect 38010 28364 38016 28376
rect 38068 28364 38074 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 28261 28203 28319 28209
rect 28261 28169 28273 28203
rect 28307 28169 28319 28203
rect 29638 28200 29644 28212
rect 29599 28172 29644 28200
rect 28261 28163 28319 28169
rect 23842 28092 23848 28144
rect 23900 28132 23906 28144
rect 28276 28132 28304 28163
rect 29638 28160 29644 28172
rect 29696 28160 29702 28212
rect 31481 28203 31539 28209
rect 31481 28169 31493 28203
rect 31527 28200 31539 28203
rect 33686 28200 33692 28212
rect 31527 28172 33692 28200
rect 31527 28169 31539 28172
rect 31481 28163 31539 28169
rect 31662 28132 31668 28144
rect 23900 28104 31668 28132
rect 23900 28092 23906 28104
rect 31662 28092 31668 28104
rect 31720 28092 31726 28144
rect 28166 28064 28172 28076
rect 28079 28036 28172 28064
rect 28166 28024 28172 28036
rect 28224 28064 28230 28076
rect 28810 28064 28816 28076
rect 28224 28036 28816 28064
rect 28224 28024 28230 28036
rect 28810 28024 28816 28036
rect 28868 28064 28874 28076
rect 30561 28067 30619 28073
rect 30561 28064 30573 28067
rect 28868 28036 30573 28064
rect 28868 28024 28874 28036
rect 30561 28033 30573 28036
rect 30607 28064 30619 28067
rect 31772 28064 31800 28172
rect 33686 28160 33692 28172
rect 33744 28160 33750 28212
rect 37826 28064 37832 28076
rect 30607 28036 31800 28064
rect 37787 28036 37832 28064
rect 30607 28033 30619 28036
rect 30561 28027 30619 28033
rect 37826 28024 37832 28036
rect 37884 28024 37890 28076
rect 29178 27956 29184 28008
rect 29236 27996 29242 28008
rect 29365 27999 29423 28005
rect 29365 27996 29377 27999
rect 29236 27968 29377 27996
rect 29236 27956 29242 27968
rect 29365 27965 29377 27968
rect 29411 27965 29423 27999
rect 29365 27959 29423 27965
rect 29549 27999 29607 28005
rect 29549 27965 29561 27999
rect 29595 27996 29607 27999
rect 30466 27996 30472 28008
rect 29595 27968 30472 27996
rect 29595 27965 29607 27968
rect 29549 27959 29607 27965
rect 29380 27928 29408 27959
rect 30466 27956 30472 27968
rect 30524 27956 30530 28008
rect 30190 27928 30196 27940
rect 29380 27900 30196 27928
rect 30190 27888 30196 27900
rect 30248 27928 30254 27940
rect 30745 27931 30803 27937
rect 30745 27928 30757 27931
rect 30248 27900 30757 27928
rect 30248 27888 30254 27900
rect 30745 27897 30757 27900
rect 30791 27897 30803 27931
rect 30745 27891 30803 27897
rect 29914 27820 29920 27872
rect 29972 27860 29978 27872
rect 30009 27863 30067 27869
rect 30009 27860 30021 27863
rect 29972 27832 30021 27860
rect 29972 27820 29978 27832
rect 30009 27829 30021 27832
rect 30055 27829 30067 27863
rect 38010 27860 38016 27872
rect 37971 27832 38016 27860
rect 30009 27823 30067 27829
rect 38010 27820 38016 27832
rect 38068 27820 38074 27872
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 28721 27659 28779 27665
rect 28721 27625 28733 27659
rect 28767 27656 28779 27659
rect 28810 27656 28816 27668
rect 28767 27628 28816 27656
rect 28767 27625 28779 27628
rect 28721 27619 28779 27625
rect 28810 27616 28816 27628
rect 28868 27616 28874 27668
rect 30101 27591 30159 27597
rect 30101 27557 30113 27591
rect 30147 27588 30159 27591
rect 37826 27588 37832 27600
rect 30147 27560 37832 27588
rect 30147 27557 30159 27560
rect 30101 27551 30159 27557
rect 37826 27548 37832 27560
rect 37884 27548 37890 27600
rect 30466 27480 30472 27532
rect 30524 27520 30530 27532
rect 30561 27523 30619 27529
rect 30561 27520 30573 27523
rect 30524 27492 30573 27520
rect 30524 27480 30530 27492
rect 30561 27489 30573 27492
rect 30607 27489 30619 27523
rect 30561 27483 30619 27489
rect 29914 27452 29920 27464
rect 29875 27424 29920 27452
rect 29914 27412 29920 27424
rect 29972 27412 29978 27464
rect 37826 27452 37832 27464
rect 37787 27424 37832 27452
rect 37826 27412 37832 27424
rect 37884 27412 37890 27464
rect 38010 27316 38016 27328
rect 37971 27288 38016 27316
rect 38010 27276 38016 27288
rect 38068 27276 38074 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 28718 27072 28724 27124
rect 28776 27112 28782 27124
rect 28905 27115 28963 27121
rect 28905 27112 28917 27115
rect 28776 27084 28917 27112
rect 28776 27072 28782 27084
rect 28905 27081 28917 27084
rect 28951 27081 28963 27115
rect 28905 27075 28963 27081
rect 29273 27115 29331 27121
rect 29273 27081 29285 27115
rect 29319 27081 29331 27115
rect 29273 27075 29331 27081
rect 29917 27115 29975 27121
rect 29917 27081 29929 27115
rect 29963 27112 29975 27115
rect 37826 27112 37832 27124
rect 29963 27084 37832 27112
rect 29963 27081 29975 27084
rect 29917 27075 29975 27081
rect 29178 26976 29184 26988
rect 28644 26948 29184 26976
rect 27982 26868 27988 26920
rect 28040 26908 28046 26920
rect 28644 26917 28672 26948
rect 29178 26936 29184 26948
rect 29236 26936 29242 26988
rect 29288 26976 29316 27075
rect 37826 27072 37832 27084
rect 37884 27072 37890 27124
rect 29733 26979 29791 26985
rect 29733 26976 29745 26979
rect 29288 26948 29745 26976
rect 29733 26945 29745 26948
rect 29779 26945 29791 26979
rect 37826 26976 37832 26988
rect 37787 26948 37832 26976
rect 29733 26939 29791 26945
rect 37826 26936 37832 26948
rect 37884 26936 37890 26988
rect 28629 26911 28687 26917
rect 28629 26908 28641 26911
rect 28040 26880 28641 26908
rect 28040 26868 28046 26880
rect 28629 26877 28641 26880
rect 28675 26877 28687 26911
rect 28629 26871 28687 26877
rect 28813 26911 28871 26917
rect 28813 26877 28825 26911
rect 28859 26908 28871 26911
rect 29086 26908 29092 26920
rect 28859 26880 29092 26908
rect 28859 26877 28871 26880
rect 28813 26871 28871 26877
rect 29086 26868 29092 26880
rect 29144 26908 29150 26920
rect 30377 26911 30435 26917
rect 30377 26908 30389 26911
rect 29144 26880 30389 26908
rect 29144 26868 29150 26880
rect 30377 26877 30389 26880
rect 30423 26877 30435 26911
rect 30377 26871 30435 26877
rect 38010 26772 38016 26784
rect 37971 26744 38016 26772
rect 38010 26732 38016 26744
rect 38068 26732 38074 26784
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 27982 26432 27988 26444
rect 27943 26404 27988 26432
rect 27982 26392 27988 26404
rect 28040 26392 28046 26444
rect 28169 26367 28227 26373
rect 28169 26333 28181 26367
rect 28215 26364 28227 26367
rect 28258 26364 28264 26376
rect 28215 26336 28264 26364
rect 28215 26333 28227 26336
rect 28169 26327 28227 26333
rect 28258 26324 28264 26336
rect 28316 26324 28322 26376
rect 28077 26299 28135 26305
rect 28077 26265 28089 26299
rect 28123 26296 28135 26299
rect 28442 26296 28448 26308
rect 28123 26268 28448 26296
rect 28123 26265 28135 26268
rect 28077 26259 28135 26265
rect 28442 26256 28448 26268
rect 28500 26296 28506 26308
rect 29549 26299 29607 26305
rect 29549 26296 29561 26299
rect 28500 26268 29561 26296
rect 28500 26256 28506 26268
rect 29549 26265 29561 26268
rect 29595 26265 29607 26299
rect 29549 26259 29607 26265
rect 28534 26228 28540 26240
rect 28495 26200 28540 26228
rect 28534 26188 28540 26200
rect 28592 26188 28598 26240
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 27338 26024 27344 26036
rect 27299 25996 27344 26024
rect 27338 25984 27344 25996
rect 27396 25984 27402 26036
rect 28997 26027 29055 26033
rect 28997 25993 29009 26027
rect 29043 26024 29055 26027
rect 37826 26024 37832 26036
rect 29043 25996 37832 26024
rect 29043 25993 29055 25996
rect 28997 25987 29055 25993
rect 37826 25984 37832 25996
rect 37884 25984 37890 26036
rect 27154 25916 27160 25968
rect 27212 25956 27218 25968
rect 27249 25959 27307 25965
rect 27249 25956 27261 25959
rect 27212 25928 27261 25956
rect 27212 25916 27218 25928
rect 27249 25925 27261 25928
rect 27295 25956 27307 25959
rect 29457 25959 29515 25965
rect 29457 25956 29469 25959
rect 27295 25928 29469 25956
rect 27295 25925 27307 25928
rect 27249 25919 27307 25925
rect 29457 25925 29469 25928
rect 29503 25925 29515 25959
rect 29457 25919 29515 25925
rect 27890 25848 27896 25900
rect 27948 25888 27954 25900
rect 28169 25891 28227 25897
rect 28169 25888 28181 25891
rect 27948 25860 28181 25888
rect 27948 25848 27954 25860
rect 28169 25857 28181 25860
rect 28215 25857 28227 25891
rect 28169 25851 28227 25857
rect 28534 25848 28540 25900
rect 28592 25888 28598 25900
rect 28813 25891 28871 25897
rect 28813 25888 28825 25891
rect 28592 25860 28825 25888
rect 28592 25848 28598 25860
rect 28813 25857 28825 25860
rect 28859 25857 28871 25891
rect 37829 25891 37887 25897
rect 37829 25888 37841 25891
rect 28813 25851 28871 25857
rect 35866 25860 37841 25888
rect 27157 25823 27215 25829
rect 27157 25789 27169 25823
rect 27203 25789 27215 25823
rect 27157 25783 27215 25789
rect 27172 25752 27200 25783
rect 27982 25752 27988 25764
rect 27172 25724 27988 25752
rect 27982 25712 27988 25724
rect 28040 25712 28046 25764
rect 28353 25755 28411 25761
rect 28353 25721 28365 25755
rect 28399 25752 28411 25755
rect 35866 25752 35894 25860
rect 37829 25857 37841 25860
rect 37875 25857 37887 25891
rect 37829 25851 37887 25857
rect 38010 25752 38016 25764
rect 28399 25724 35894 25752
rect 37971 25724 38016 25752
rect 28399 25721 28411 25724
rect 28353 25715 28411 25721
rect 38010 25712 38016 25724
rect 38068 25712 38074 25764
rect 27706 25684 27712 25696
rect 27667 25656 27712 25684
rect 27706 25644 27712 25656
rect 27764 25644 27770 25696
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 27890 25480 27896 25492
rect 27851 25452 27896 25480
rect 27890 25440 27896 25452
rect 27948 25440 27954 25492
rect 27341 25347 27399 25353
rect 27341 25313 27353 25347
rect 27387 25344 27399 25347
rect 27982 25344 27988 25356
rect 27387 25316 27988 25344
rect 27387 25313 27399 25316
rect 27341 25307 27399 25313
rect 27982 25304 27988 25316
rect 28040 25304 28046 25356
rect 27522 25276 27528 25288
rect 27483 25248 27528 25276
rect 27522 25236 27528 25248
rect 27580 25236 27586 25288
rect 27706 25236 27712 25288
rect 27764 25276 27770 25288
rect 28353 25279 28411 25285
rect 28353 25276 28365 25279
rect 27764 25248 28365 25276
rect 27764 25236 27770 25248
rect 28353 25245 28365 25248
rect 28399 25245 28411 25279
rect 37829 25279 37887 25285
rect 37829 25276 37841 25279
rect 28353 25239 28411 25245
rect 35866 25248 37841 25276
rect 27433 25143 27491 25149
rect 27433 25109 27445 25143
rect 27479 25140 27491 25143
rect 27798 25140 27804 25152
rect 27479 25112 27804 25140
rect 27479 25109 27491 25112
rect 27433 25103 27491 25109
rect 27798 25100 27804 25112
rect 27856 25100 27862 25152
rect 28537 25143 28595 25149
rect 28537 25109 28549 25143
rect 28583 25140 28595 25143
rect 35866 25140 35894 25248
rect 37829 25245 37841 25248
rect 37875 25245 37887 25279
rect 37829 25239 37887 25245
rect 38010 25140 38016 25152
rect 28583 25112 35894 25140
rect 37971 25112 38016 25140
rect 28583 25109 28595 25112
rect 28537 25103 28595 25109
rect 38010 25100 38016 25112
rect 38068 25100 38074 25152
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 26786 24760 26792 24812
rect 26844 24800 26850 24812
rect 37829 24803 37887 24809
rect 37829 24800 37841 24803
rect 26844 24772 37841 24800
rect 26844 24760 26850 24772
rect 37829 24769 37841 24772
rect 37875 24769 37887 24803
rect 37829 24763 37887 24769
rect 26050 24556 26056 24608
rect 26108 24596 26114 24608
rect 26237 24599 26295 24605
rect 26237 24596 26249 24599
rect 26108 24568 26249 24596
rect 26108 24556 26114 24568
rect 26237 24565 26249 24568
rect 26283 24565 26295 24599
rect 26237 24559 26295 24565
rect 27798 24556 27804 24608
rect 27856 24596 27862 24608
rect 27985 24599 28043 24605
rect 27985 24596 27997 24599
rect 27856 24568 27997 24596
rect 27856 24556 27862 24568
rect 27985 24565 27997 24568
rect 28031 24565 28043 24599
rect 38010 24596 38016 24608
rect 37971 24568 38016 24596
rect 27985 24559 28043 24565
rect 38010 24556 38016 24568
rect 38068 24556 38074 24608
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 26786 24392 26792 24404
rect 26747 24364 26792 24392
rect 26786 24352 26792 24364
rect 26844 24352 26850 24404
rect 26145 24327 26203 24333
rect 26145 24293 26157 24327
rect 26191 24293 26203 24327
rect 26145 24287 26203 24293
rect 24486 24216 24492 24268
rect 24544 24256 24550 24268
rect 25501 24259 25559 24265
rect 25501 24256 25513 24259
rect 24544 24228 25513 24256
rect 24544 24216 24550 24228
rect 25501 24225 25513 24228
rect 25547 24225 25559 24259
rect 25501 24219 25559 24225
rect 25774 24188 25780 24200
rect 25735 24160 25780 24188
rect 25774 24148 25780 24160
rect 25832 24148 25838 24200
rect 26160 24188 26188 24287
rect 26605 24191 26663 24197
rect 26605 24188 26617 24191
rect 26160 24160 26617 24188
rect 26605 24157 26617 24160
rect 26651 24157 26663 24191
rect 37826 24188 37832 24200
rect 37787 24160 37832 24188
rect 26605 24151 26663 24157
rect 37826 24148 37832 24160
rect 37884 24148 37890 24200
rect 25685 24055 25743 24061
rect 25685 24021 25697 24055
rect 25731 24052 25743 24055
rect 26050 24052 26056 24064
rect 25731 24024 26056 24052
rect 25731 24021 25743 24024
rect 25685 24015 25743 24021
rect 26050 24012 26056 24024
rect 26108 24012 26114 24064
rect 38010 24052 38016 24064
rect 37971 24024 38016 24052
rect 38010 24012 38016 24024
rect 38068 24012 38074 24064
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 25225 23851 25283 23857
rect 25225 23817 25237 23851
rect 25271 23848 25283 23851
rect 25314 23848 25320 23860
rect 25271 23820 25320 23848
rect 25271 23817 25283 23820
rect 25225 23811 25283 23817
rect 25314 23808 25320 23820
rect 25372 23808 25378 23860
rect 25593 23851 25651 23857
rect 25593 23817 25605 23851
rect 25639 23817 25651 23851
rect 25593 23811 25651 23817
rect 25608 23712 25636 23811
rect 26053 23715 26111 23721
rect 26053 23712 26065 23715
rect 25608 23684 26065 23712
rect 26053 23681 26065 23684
rect 26099 23681 26111 23715
rect 26053 23675 26111 23681
rect 24486 23604 24492 23656
rect 24544 23644 24550 23656
rect 24949 23647 25007 23653
rect 24949 23644 24961 23647
rect 24544 23616 24961 23644
rect 24544 23604 24550 23616
rect 24949 23613 24961 23616
rect 24995 23613 25007 23647
rect 24949 23607 25007 23613
rect 25133 23647 25191 23653
rect 25133 23613 25145 23647
rect 25179 23644 25191 23647
rect 26234 23644 26240 23656
rect 25179 23616 26240 23644
rect 25179 23613 25191 23616
rect 25133 23607 25191 23613
rect 26234 23604 26240 23616
rect 26292 23604 26298 23656
rect 23014 23536 23020 23588
rect 23072 23576 23078 23588
rect 23569 23579 23627 23585
rect 23569 23576 23581 23579
rect 23072 23548 23581 23576
rect 23072 23536 23078 23548
rect 23569 23545 23581 23548
rect 23615 23576 23627 23579
rect 28166 23576 28172 23588
rect 23615 23548 28172 23576
rect 23615 23545 23627 23548
rect 23569 23539 23627 23545
rect 28166 23536 28172 23548
rect 28224 23536 28230 23588
rect 26237 23511 26295 23517
rect 26237 23477 26249 23511
rect 26283 23508 26295 23511
rect 37826 23508 37832 23520
rect 26283 23480 37832 23508
rect 26283 23477 26295 23480
rect 26237 23471 26295 23477
rect 37826 23468 37832 23480
rect 37884 23468 37890 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 36814 23304 36820 23316
rect 36775 23276 36820 23304
rect 36814 23264 36820 23276
rect 36872 23264 36878 23316
rect 23106 23128 23112 23180
rect 23164 23168 23170 23180
rect 24486 23168 24492 23180
rect 23164 23140 24492 23168
rect 23164 23128 23170 23140
rect 24486 23128 24492 23140
rect 24544 23128 24550 23180
rect 24673 23171 24731 23177
rect 24673 23137 24685 23171
rect 24719 23168 24731 23171
rect 25222 23168 25228 23180
rect 24719 23140 25228 23168
rect 24719 23137 24731 23140
rect 24673 23131 24731 23137
rect 25222 23128 25228 23140
rect 25280 23128 25286 23180
rect 23014 23100 23020 23112
rect 22975 23072 23020 23100
rect 23014 23060 23020 23072
rect 23072 23060 23078 23112
rect 24762 23100 24768 23112
rect 24723 23072 24768 23100
rect 24762 23060 24768 23072
rect 24820 23060 24826 23112
rect 25593 23103 25651 23109
rect 25593 23100 25605 23103
rect 25148 23072 25605 23100
rect 23106 22964 23112 22976
rect 23067 22936 23112 22964
rect 23106 22924 23112 22936
rect 23164 22924 23170 22976
rect 25148 22973 25176 23072
rect 25593 23069 25605 23072
rect 25639 23069 25651 23103
rect 25593 23063 25651 23069
rect 36722 23060 36728 23112
rect 36780 23100 36786 23112
rect 37001 23103 37059 23109
rect 37001 23100 37013 23103
rect 36780 23072 37013 23100
rect 36780 23060 36786 23072
rect 37001 23069 37013 23072
rect 37047 23069 37059 23103
rect 37001 23063 37059 23069
rect 37829 23103 37887 23109
rect 37829 23069 37841 23103
rect 37875 23069 37887 23103
rect 37829 23063 37887 23069
rect 37844 23032 37872 23063
rect 25792 23004 37872 23032
rect 25792 22973 25820 23004
rect 25133 22967 25191 22973
rect 25133 22933 25145 22967
rect 25179 22933 25191 22967
rect 25133 22927 25191 22933
rect 25777 22967 25835 22973
rect 25777 22933 25789 22967
rect 25823 22933 25835 22967
rect 25777 22927 25835 22933
rect 26234 22924 26240 22976
rect 26292 22964 26298 22976
rect 38010 22964 38016 22976
rect 26292 22936 26337 22964
rect 37971 22936 38016 22964
rect 26292 22924 26298 22936
rect 38010 22924 38016 22936
rect 38068 22924 38074 22976
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 23750 22760 23756 22772
rect 23711 22732 23756 22760
rect 23750 22720 23756 22732
rect 23808 22720 23814 22772
rect 24121 22763 24179 22769
rect 24121 22729 24133 22763
rect 24167 22729 24179 22763
rect 36354 22760 36360 22772
rect 36315 22732 36360 22760
rect 24121 22723 24179 22729
rect 24136 22624 24164 22723
rect 36354 22720 36360 22732
rect 36412 22720 36418 22772
rect 36722 22760 36728 22772
rect 36683 22732 36728 22760
rect 36722 22720 36728 22732
rect 36780 22720 36786 22772
rect 24581 22627 24639 22633
rect 24581 22624 24593 22627
rect 24136 22596 24593 22624
rect 24581 22593 24593 22596
rect 24627 22593 24639 22627
rect 37829 22627 37887 22633
rect 37829 22624 37841 22627
rect 24581 22587 24639 22593
rect 26206 22596 37841 22624
rect 22738 22516 22744 22568
rect 22796 22556 22802 22568
rect 23106 22556 23112 22568
rect 22796 22528 23112 22556
rect 22796 22516 22802 22528
rect 23106 22516 23112 22528
rect 23164 22556 23170 22568
rect 23477 22559 23535 22565
rect 23477 22556 23489 22559
rect 23164 22528 23489 22556
rect 23164 22516 23170 22528
rect 23477 22525 23489 22528
rect 23523 22525 23535 22559
rect 23477 22519 23535 22525
rect 23661 22559 23719 22565
rect 23661 22525 23673 22559
rect 23707 22525 23719 22559
rect 23661 22519 23719 22525
rect 23676 22488 23704 22519
rect 24578 22488 24584 22500
rect 23676 22460 24584 22488
rect 24578 22448 24584 22460
rect 24636 22448 24642 22500
rect 24765 22491 24823 22497
rect 24765 22457 24777 22491
rect 24811 22488 24823 22491
rect 26206 22488 26234 22596
rect 37829 22593 37841 22596
rect 37875 22593 37887 22627
rect 37829 22587 37887 22593
rect 36081 22559 36139 22565
rect 36081 22556 36093 22559
rect 24811 22460 26234 22488
rect 35866 22528 36093 22556
rect 24811 22457 24823 22460
rect 24765 22451 24823 22457
rect 25222 22420 25228 22432
rect 25183 22392 25228 22420
rect 25222 22380 25228 22392
rect 25280 22380 25286 22432
rect 25314 22380 25320 22432
rect 25372 22420 25378 22432
rect 35437 22423 35495 22429
rect 35437 22420 35449 22423
rect 25372 22392 35449 22420
rect 25372 22380 25378 22392
rect 35437 22389 35449 22392
rect 35483 22420 35495 22423
rect 35866 22420 35894 22528
rect 36081 22525 36093 22528
rect 36127 22525 36139 22559
rect 36081 22519 36139 22525
rect 36265 22559 36323 22565
rect 36265 22525 36277 22559
rect 36311 22556 36323 22559
rect 36630 22556 36636 22568
rect 36311 22528 36636 22556
rect 36311 22525 36323 22528
rect 36265 22519 36323 22525
rect 36630 22516 36636 22528
rect 36688 22556 36694 22568
rect 37277 22559 37335 22565
rect 37277 22556 37289 22559
rect 36688 22528 37289 22556
rect 36688 22516 36694 22528
rect 37277 22525 37289 22528
rect 37323 22525 37335 22559
rect 37277 22519 37335 22525
rect 38010 22420 38016 22432
rect 35483 22392 35894 22420
rect 37971 22392 38016 22420
rect 35483 22389 35495 22392
rect 35437 22383 35495 22389
rect 38010 22380 38016 22392
rect 38068 22380 38074 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 20254 22176 20260 22228
rect 20312 22216 20318 22228
rect 25314 22216 25320 22228
rect 20312 22188 25320 22216
rect 20312 22176 20318 22188
rect 25314 22176 25320 22188
rect 25372 22176 25378 22228
rect 22370 21972 22376 22024
rect 22428 22012 22434 22024
rect 22465 22015 22523 22021
rect 22465 22012 22477 22015
rect 22428 21984 22477 22012
rect 22428 21972 22434 21984
rect 22465 21981 22477 21984
rect 22511 21981 22523 22015
rect 37826 22012 37832 22024
rect 37787 21984 37832 22012
rect 22465 21975 22523 21981
rect 37826 21972 37832 21984
rect 37884 21972 37890 22024
rect 22278 21876 22284 21888
rect 22239 21848 22284 21876
rect 22278 21836 22284 21848
rect 22336 21836 22342 21888
rect 23290 21836 23296 21888
rect 23348 21876 23354 21888
rect 23477 21879 23535 21885
rect 23477 21876 23489 21879
rect 23348 21848 23489 21876
rect 23348 21836 23354 21848
rect 23477 21845 23489 21848
rect 23523 21845 23535 21879
rect 23477 21839 23535 21845
rect 24489 21879 24547 21885
rect 24489 21845 24501 21879
rect 24535 21876 24547 21879
rect 24578 21876 24584 21888
rect 24535 21848 24584 21876
rect 24535 21845 24547 21848
rect 24489 21839 24547 21845
rect 24578 21836 24584 21848
rect 24636 21836 24642 21888
rect 38010 21876 38016 21888
rect 37971 21848 38016 21876
rect 38010 21836 38016 21848
rect 38068 21836 38074 21888
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 22830 21632 22836 21684
rect 22888 21672 22894 21684
rect 23017 21675 23075 21681
rect 23017 21672 23029 21675
rect 22888 21644 23029 21672
rect 22888 21632 22894 21644
rect 23017 21641 23029 21644
rect 23063 21641 23075 21675
rect 23017 21635 23075 21641
rect 23385 21675 23443 21681
rect 23385 21641 23397 21675
rect 23431 21641 23443 21675
rect 23385 21635 23443 21641
rect 23400 21536 23428 21635
rect 23845 21539 23903 21545
rect 23845 21536 23857 21539
rect 23400 21508 23857 21536
rect 23845 21505 23857 21508
rect 23891 21505 23903 21539
rect 23845 21499 23903 21505
rect 37461 21539 37519 21545
rect 37461 21505 37473 21539
rect 37507 21536 37519 21539
rect 38102 21536 38108 21548
rect 37507 21508 38108 21536
rect 37507 21505 37519 21508
rect 37461 21499 37519 21505
rect 38102 21496 38108 21508
rect 38160 21496 38166 21548
rect 22738 21468 22744 21480
rect 22699 21440 22744 21468
rect 22738 21428 22744 21440
rect 22796 21428 22802 21480
rect 22925 21471 22983 21477
rect 22925 21437 22937 21471
rect 22971 21468 22983 21471
rect 23290 21468 23296 21480
rect 22971 21440 23296 21468
rect 22971 21437 22983 21440
rect 22925 21431 22983 21437
rect 23290 21428 23296 21440
rect 23348 21428 23354 21480
rect 24026 21332 24032 21344
rect 23987 21304 24032 21332
rect 24026 21292 24032 21304
rect 24084 21292 24090 21344
rect 37918 21332 37924 21344
rect 37879 21304 37924 21332
rect 37918 21292 37924 21304
rect 37976 21292 37982 21344
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 22370 21128 22376 21140
rect 22331 21100 22376 21128
rect 22370 21088 22376 21100
rect 22428 21088 22434 21140
rect 23753 21131 23811 21137
rect 23753 21097 23765 21131
rect 23799 21128 23811 21131
rect 23842 21128 23848 21140
rect 23799 21100 23848 21128
rect 23799 21097 23811 21100
rect 23753 21091 23811 21097
rect 23842 21088 23848 21100
rect 23900 21088 23906 21140
rect 24026 21088 24032 21140
rect 24084 21128 24090 21140
rect 37826 21128 37832 21140
rect 24084 21100 37832 21128
rect 24084 21088 24090 21100
rect 37826 21088 37832 21100
rect 37884 21088 37890 21140
rect 22281 21063 22339 21069
rect 22281 21029 22293 21063
rect 22327 21060 22339 21063
rect 22327 21032 23060 21060
rect 22327 21029 22339 21032
rect 22281 21023 22339 21029
rect 12618 20884 12624 20936
rect 12676 20924 12682 20936
rect 23032 20933 23060 21032
rect 21913 20927 21971 20933
rect 21913 20924 21925 20927
rect 12676 20896 21925 20924
rect 12676 20884 12682 20896
rect 21913 20893 21925 20896
rect 21959 20924 21971 20927
rect 22925 20927 22983 20933
rect 22925 20924 22937 20927
rect 21959 20896 22937 20924
rect 21959 20893 21971 20896
rect 21913 20887 21971 20893
rect 22925 20893 22937 20896
rect 22971 20893 22983 20927
rect 22925 20887 22983 20893
rect 23017 20927 23075 20933
rect 23017 20893 23029 20927
rect 23063 20924 23075 20927
rect 37918 20924 37924 20936
rect 23063 20896 37924 20924
rect 23063 20893 23075 20896
rect 23017 20887 23075 20893
rect 22940 20856 22968 20887
rect 37918 20884 37924 20896
rect 37976 20884 37982 20936
rect 23842 20856 23848 20868
rect 22940 20828 23848 20856
rect 23842 20816 23848 20828
rect 23900 20816 23906 20868
rect 23198 20788 23204 20800
rect 23159 20760 23204 20788
rect 23198 20748 23204 20760
rect 23256 20748 23262 20800
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 22186 20584 22192 20596
rect 22147 20556 22192 20584
rect 22186 20544 22192 20556
rect 22244 20544 22250 20596
rect 23753 20587 23811 20593
rect 23753 20553 23765 20587
rect 23799 20584 23811 20587
rect 23842 20584 23848 20596
rect 23799 20556 23848 20584
rect 23799 20553 23811 20556
rect 23753 20547 23811 20553
rect 23842 20544 23848 20556
rect 23900 20544 23906 20596
rect 23198 20448 23204 20460
rect 23159 20420 23204 20448
rect 23198 20408 23204 20420
rect 23256 20408 23262 20460
rect 31018 20408 31024 20460
rect 31076 20448 31082 20460
rect 37829 20451 37887 20457
rect 37829 20448 37841 20451
rect 31076 20420 37841 20448
rect 31076 20408 31082 20420
rect 37829 20417 37841 20420
rect 37875 20417 37887 20451
rect 37829 20411 37887 20417
rect 22002 20340 22008 20392
rect 22060 20380 22066 20392
rect 22281 20383 22339 20389
rect 22281 20380 22293 20383
rect 22060 20352 22293 20380
rect 22060 20340 22066 20352
rect 22281 20349 22293 20352
rect 22327 20349 22339 20383
rect 22281 20343 22339 20349
rect 22373 20383 22431 20389
rect 22373 20349 22385 20383
rect 22419 20380 22431 20383
rect 22738 20380 22744 20392
rect 22419 20352 22744 20380
rect 22419 20349 22431 20352
rect 22373 20343 22431 20349
rect 20438 20272 20444 20324
rect 20496 20312 20502 20324
rect 22388 20312 22416 20343
rect 22738 20340 22744 20352
rect 22796 20340 22802 20392
rect 38010 20312 38016 20324
rect 20496 20284 22416 20312
rect 37971 20284 38016 20312
rect 20496 20272 20502 20284
rect 38010 20272 38016 20284
rect 38068 20272 38074 20324
rect 21818 20244 21824 20256
rect 21779 20216 21824 20244
rect 21818 20204 21824 20216
rect 21876 20204 21882 20256
rect 22922 20204 22928 20256
rect 22980 20244 22986 20256
rect 23017 20247 23075 20253
rect 23017 20244 23029 20247
rect 22980 20216 23029 20244
rect 22980 20204 22986 20216
rect 23017 20213 23029 20216
rect 23063 20213 23075 20247
rect 23017 20207 23075 20213
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 19889 20043 19947 20049
rect 19889 20009 19901 20043
rect 19935 20040 19947 20043
rect 20898 20040 20904 20052
rect 19935 20012 20904 20040
rect 19935 20009 19947 20012
rect 19889 20003 19947 20009
rect 20898 20000 20904 20012
rect 20956 20040 20962 20052
rect 23014 20040 23020 20052
rect 20956 20012 23020 20040
rect 20956 20000 20962 20012
rect 23014 20000 23020 20012
rect 23072 20000 23078 20052
rect 20438 19864 20444 19916
rect 20496 19904 20502 19916
rect 20533 19907 20591 19913
rect 20533 19904 20545 19907
rect 20496 19876 20545 19904
rect 20496 19864 20502 19876
rect 20533 19873 20545 19876
rect 20579 19873 20591 19907
rect 20533 19867 20591 19873
rect 20806 19836 20812 19848
rect 20767 19808 20812 19836
rect 20806 19796 20812 19808
rect 20864 19796 20870 19848
rect 21818 19836 21824 19848
rect 21779 19808 21824 19836
rect 21818 19796 21824 19808
rect 21876 19796 21882 19848
rect 37826 19836 37832 19848
rect 37787 19808 37832 19836
rect 37826 19796 37832 19808
rect 37884 19796 37890 19848
rect 20714 19700 20720 19712
rect 20675 19672 20720 19700
rect 20714 19660 20720 19672
rect 20772 19660 20778 19712
rect 21082 19660 21088 19712
rect 21140 19700 21146 19712
rect 21177 19703 21235 19709
rect 21177 19700 21189 19703
rect 21140 19672 21189 19700
rect 21140 19660 21146 19672
rect 21177 19669 21189 19672
rect 21223 19669 21235 19703
rect 21177 19663 21235 19669
rect 22005 19703 22063 19709
rect 22005 19669 22017 19703
rect 22051 19700 22063 19703
rect 31018 19700 31024 19712
rect 22051 19672 31024 19700
rect 22051 19669 22063 19672
rect 22005 19663 22063 19669
rect 31018 19660 31024 19672
rect 31076 19660 31082 19712
rect 38010 19700 38016 19712
rect 37971 19672 38016 19700
rect 38010 19660 38016 19672
rect 38068 19660 38074 19712
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 21269 19499 21327 19505
rect 21269 19465 21281 19499
rect 21315 19496 21327 19499
rect 37826 19496 37832 19508
rect 21315 19468 37832 19496
rect 21315 19465 21327 19468
rect 21269 19459 21327 19465
rect 37826 19456 37832 19468
rect 37884 19456 37890 19508
rect 19613 19431 19671 19437
rect 19613 19397 19625 19431
rect 19659 19428 19671 19431
rect 20898 19428 20904 19440
rect 19659 19400 20904 19428
rect 19659 19397 19671 19400
rect 19613 19391 19671 19397
rect 20898 19388 20904 19400
rect 20956 19388 20962 19440
rect 21082 19360 21088 19372
rect 21043 19332 21088 19360
rect 21082 19320 21088 19332
rect 21140 19320 21146 19372
rect 34514 19320 34520 19372
rect 34572 19360 34578 19372
rect 37829 19363 37887 19369
rect 37829 19360 37841 19363
rect 34572 19332 37841 19360
rect 34572 19320 34578 19332
rect 37829 19329 37841 19332
rect 37875 19329 37887 19363
rect 37829 19323 37887 19329
rect 20162 19252 20168 19304
rect 20220 19292 20226 19304
rect 20530 19292 20536 19304
rect 20220 19264 20536 19292
rect 20220 19252 20226 19264
rect 20530 19252 20536 19264
rect 20588 19252 20594 19304
rect 17954 19116 17960 19168
rect 18012 19156 18018 19168
rect 19337 19159 19395 19165
rect 19337 19156 19349 19159
rect 18012 19128 19349 19156
rect 18012 19116 18018 19128
rect 19337 19125 19349 19128
rect 19383 19125 19395 19159
rect 38010 19156 38016 19168
rect 37971 19128 38016 19156
rect 19337 19119 19395 19125
rect 38010 19116 38016 19128
rect 38068 19116 38074 19168
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 19334 18776 19340 18828
rect 19392 18816 19398 18828
rect 19797 18819 19855 18825
rect 19797 18816 19809 18819
rect 19392 18788 19809 18816
rect 19392 18776 19398 18788
rect 19797 18785 19809 18788
rect 19843 18816 19855 18819
rect 20438 18816 20444 18828
rect 19843 18788 20444 18816
rect 19843 18785 19855 18788
rect 19797 18779 19855 18785
rect 20438 18776 20444 18788
rect 20496 18776 20502 18828
rect 19981 18751 20039 18757
rect 19981 18717 19993 18751
rect 20027 18748 20039 18751
rect 20070 18748 20076 18760
rect 20027 18720 20076 18748
rect 20027 18717 20039 18720
rect 19981 18711 20039 18717
rect 20070 18708 20076 18720
rect 20128 18708 20134 18760
rect 20901 18751 20959 18757
rect 20901 18748 20913 18751
rect 20456 18720 20913 18748
rect 20073 18615 20131 18621
rect 20073 18581 20085 18615
rect 20119 18612 20131 18615
rect 20162 18612 20168 18624
rect 20119 18584 20168 18612
rect 20119 18581 20131 18584
rect 20073 18575 20131 18581
rect 20162 18572 20168 18584
rect 20220 18572 20226 18624
rect 20456 18621 20484 18720
rect 20901 18717 20913 18720
rect 20947 18717 20959 18751
rect 37826 18748 37832 18760
rect 37787 18720 37832 18748
rect 20901 18711 20959 18717
rect 37826 18708 37832 18720
rect 37884 18708 37890 18760
rect 20441 18615 20499 18621
rect 20441 18581 20453 18615
rect 20487 18581 20499 18615
rect 20441 18575 20499 18581
rect 21085 18615 21143 18621
rect 21085 18581 21097 18615
rect 21131 18612 21143 18615
rect 34514 18612 34520 18624
rect 21131 18584 34520 18612
rect 21131 18581 21143 18584
rect 21085 18575 21143 18581
rect 34514 18572 34520 18584
rect 34572 18572 34578 18624
rect 38010 18612 38016 18624
rect 37971 18584 38016 18612
rect 38010 18572 38016 18584
rect 38068 18572 38074 18624
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 18230 18408 18236 18420
rect 18191 18380 18236 18408
rect 18230 18368 18236 18380
rect 18288 18368 18294 18420
rect 19426 18408 19432 18420
rect 19387 18380 19432 18408
rect 19426 18368 19432 18380
rect 19484 18368 19490 18420
rect 19797 18411 19855 18417
rect 19797 18377 19809 18411
rect 19843 18377 19855 18411
rect 19797 18371 19855 18377
rect 19334 18340 19340 18352
rect 19168 18312 19340 18340
rect 18049 18207 18107 18213
rect 18049 18173 18061 18207
rect 18095 18173 18107 18207
rect 18049 18167 18107 18173
rect 18141 18207 18199 18213
rect 18141 18173 18153 18207
rect 18187 18204 18199 18207
rect 18506 18204 18512 18216
rect 18187 18176 18512 18204
rect 18187 18173 18199 18176
rect 18141 18167 18199 18173
rect 18064 18136 18092 18167
rect 18506 18164 18512 18176
rect 18564 18164 18570 18216
rect 19168 18213 19196 18312
rect 19334 18300 19340 18312
rect 19392 18300 19398 18352
rect 19812 18272 19840 18371
rect 20257 18275 20315 18281
rect 20257 18272 20269 18275
rect 19812 18244 20269 18272
rect 20257 18241 20269 18244
rect 20303 18241 20315 18275
rect 20257 18235 20315 18241
rect 19153 18207 19211 18213
rect 19153 18173 19165 18207
rect 19199 18173 19211 18207
rect 19153 18167 19211 18173
rect 19337 18207 19395 18213
rect 19337 18173 19349 18207
rect 19383 18204 19395 18207
rect 20346 18204 20352 18216
rect 19383 18176 20352 18204
rect 19383 18173 19395 18176
rect 19337 18167 19395 18173
rect 19168 18136 19196 18167
rect 20346 18164 20352 18176
rect 20404 18164 20410 18216
rect 18064 18108 19196 18136
rect 18601 18071 18659 18077
rect 18601 18037 18613 18071
rect 18647 18068 18659 18071
rect 19334 18068 19340 18080
rect 18647 18040 19340 18068
rect 18647 18037 18659 18040
rect 18601 18031 18659 18037
rect 19334 18028 19340 18040
rect 19392 18028 19398 18080
rect 20441 18071 20499 18077
rect 20441 18037 20453 18071
rect 20487 18068 20499 18071
rect 37826 18068 37832 18080
rect 20487 18040 37832 18068
rect 20487 18037 20499 18040
rect 20441 18031 20499 18037
rect 37826 18028 37832 18040
rect 37884 18028 37890 18080
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 18230 17824 18236 17876
rect 18288 17864 18294 17876
rect 18601 17867 18659 17873
rect 18601 17864 18613 17867
rect 18288 17836 18613 17864
rect 18288 17824 18294 17836
rect 18601 17833 18613 17836
rect 18647 17833 18659 17867
rect 18601 17827 18659 17833
rect 19426 17824 19432 17876
rect 19484 17864 19490 17876
rect 19981 17867 20039 17873
rect 19981 17864 19993 17867
rect 19484 17836 19993 17864
rect 19484 17824 19490 17836
rect 19981 17833 19993 17836
rect 20027 17833 20039 17867
rect 19981 17827 20039 17833
rect 19334 17660 19340 17672
rect 19295 17632 19340 17660
rect 19334 17620 19340 17632
rect 19392 17620 19398 17672
rect 37829 17663 37887 17669
rect 37829 17629 37841 17663
rect 37875 17629 37887 17663
rect 37829 17623 37887 17629
rect 37277 17595 37335 17601
rect 37277 17592 37289 17595
rect 19536 17564 37289 17592
rect 19536 17533 19564 17564
rect 37277 17561 37289 17564
rect 37323 17592 37335 17595
rect 37844 17592 37872 17623
rect 37323 17564 37872 17592
rect 37323 17561 37335 17564
rect 37277 17555 37335 17561
rect 19521 17527 19579 17533
rect 19521 17493 19533 17527
rect 19567 17493 19579 17527
rect 38010 17524 38016 17536
rect 37971 17496 38016 17524
rect 19521 17487 19579 17493
rect 38010 17484 38016 17496
rect 38068 17484 38074 17536
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 18138 17184 18144 17196
rect 18099 17156 18144 17184
rect 18138 17144 18144 17156
rect 18196 17144 18202 17196
rect 37829 17187 37887 17193
rect 37829 17184 37841 17187
rect 37292 17156 37841 17184
rect 37292 16989 37320 17156
rect 37829 17153 37841 17156
rect 37875 17153 37887 17187
rect 37829 17147 37887 17153
rect 18325 16983 18383 16989
rect 18325 16949 18337 16983
rect 18371 16980 18383 16983
rect 37277 16983 37335 16989
rect 37277 16980 37289 16983
rect 18371 16952 37289 16980
rect 18371 16949 18383 16952
rect 18325 16943 18383 16949
rect 37277 16949 37289 16952
rect 37323 16949 37335 16983
rect 38010 16980 38016 16992
rect 37971 16952 38016 16980
rect 37277 16943 37335 16949
rect 38010 16940 38016 16952
rect 38068 16940 38074 16992
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 18138 16736 18144 16788
rect 18196 16776 18202 16788
rect 18325 16779 18383 16785
rect 18325 16776 18337 16779
rect 18196 16748 18337 16776
rect 18196 16736 18202 16748
rect 18325 16745 18337 16748
rect 18371 16745 18383 16779
rect 20898 16776 20904 16788
rect 20859 16748 20904 16776
rect 18325 16739 18383 16745
rect 20898 16736 20904 16748
rect 20956 16736 20962 16788
rect 17954 16708 17960 16720
rect 17788 16680 17960 16708
rect 17788 16649 17816 16680
rect 17954 16668 17960 16680
rect 18012 16668 18018 16720
rect 17773 16643 17831 16649
rect 17773 16609 17785 16643
rect 17819 16609 17831 16643
rect 17773 16603 17831 16609
rect 17865 16643 17923 16649
rect 17865 16609 17877 16643
rect 17911 16640 17923 16643
rect 18138 16640 18144 16652
rect 17911 16612 18144 16640
rect 17911 16609 17923 16612
rect 17865 16603 17923 16609
rect 18138 16600 18144 16612
rect 18196 16600 18202 16652
rect 20441 16575 20499 16581
rect 20441 16541 20453 16575
rect 20487 16572 20499 16575
rect 20898 16572 20904 16584
rect 20487 16544 20904 16572
rect 20487 16541 20499 16544
rect 20441 16535 20499 16541
rect 20898 16532 20904 16544
rect 20956 16532 20962 16584
rect 37829 16575 37887 16581
rect 37829 16572 37841 16575
rect 37292 16544 37841 16572
rect 17957 16507 18015 16513
rect 17957 16473 17969 16507
rect 18003 16504 18015 16507
rect 18046 16504 18052 16516
rect 18003 16476 18052 16504
rect 18003 16473 18015 16476
rect 17957 16467 18015 16473
rect 18046 16464 18052 16476
rect 18104 16504 18110 16516
rect 19245 16507 19303 16513
rect 19245 16504 19257 16507
rect 18104 16476 19257 16504
rect 18104 16464 18110 16476
rect 19245 16473 19257 16476
rect 19291 16473 19303 16507
rect 20162 16504 20168 16516
rect 20123 16476 20168 16504
rect 19245 16467 19303 16473
rect 20162 16464 20168 16476
rect 20220 16464 20226 16516
rect 37292 16448 37320 16544
rect 37829 16541 37841 16544
rect 37875 16541 37887 16575
rect 37829 16535 37887 16541
rect 37274 16436 37280 16448
rect 37235 16408 37280 16436
rect 37274 16396 37280 16408
rect 37332 16396 37338 16448
rect 38010 16436 38016 16448
rect 37971 16408 38016 16436
rect 38010 16396 38016 16408
rect 38068 16396 38074 16448
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 17497 16235 17555 16241
rect 17497 16201 17509 16235
rect 17543 16201 17555 16235
rect 17497 16195 17555 16201
rect 17129 16099 17187 16105
rect 17129 16065 17141 16099
rect 17175 16096 17187 16099
rect 17512 16096 17540 16195
rect 37274 16164 37280 16176
rect 26206 16136 37280 16164
rect 17957 16099 18015 16105
rect 17957 16096 17969 16099
rect 17175 16068 17448 16096
rect 17512 16068 17969 16096
rect 17175 16065 17187 16068
rect 17129 16059 17187 16065
rect 16206 15988 16212 16040
rect 16264 16028 16270 16040
rect 16945 16031 17003 16037
rect 16945 16028 16957 16031
rect 16264 16000 16957 16028
rect 16264 15988 16270 16000
rect 16945 15997 16957 16000
rect 16991 15997 17003 16031
rect 16945 15991 17003 15997
rect 17037 16031 17095 16037
rect 17037 15997 17049 16031
rect 17083 16028 17095 16031
rect 17310 16028 17316 16040
rect 17083 16000 17316 16028
rect 17083 15997 17095 16000
rect 17037 15991 17095 15997
rect 16960 15960 16988 15991
rect 17310 15988 17316 16000
rect 17368 15988 17374 16040
rect 17420 16028 17448 16068
rect 17957 16065 17969 16068
rect 18003 16065 18015 16099
rect 17957 16059 18015 16065
rect 17862 16028 17868 16040
rect 17420 16000 17868 16028
rect 17862 15988 17868 16000
rect 17920 15988 17926 16040
rect 17954 15960 17960 15972
rect 16960 15932 17960 15960
rect 17954 15920 17960 15932
rect 18012 15920 18018 15972
rect 18141 15895 18199 15901
rect 18141 15861 18153 15895
rect 18187 15892 18199 15895
rect 26206 15892 26234 16136
rect 37274 16124 37280 16136
rect 37332 16124 37338 16176
rect 37829 16099 37887 16105
rect 37829 16096 37841 16099
rect 37292 16068 37841 16096
rect 37292 15904 37320 16068
rect 37829 16065 37841 16068
rect 37875 16065 37887 16099
rect 37829 16059 37887 16065
rect 37274 15892 37280 15904
rect 18187 15864 26234 15892
rect 37235 15864 37280 15892
rect 18187 15861 18199 15864
rect 18141 15855 18199 15861
rect 37274 15852 37280 15864
rect 37332 15852 37338 15904
rect 38010 15892 38016 15904
rect 37971 15864 38016 15892
rect 38010 15852 38016 15864
rect 38068 15852 38074 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 17862 15688 17868 15700
rect 17823 15660 17868 15688
rect 17862 15648 17868 15660
rect 17920 15648 17926 15700
rect 16761 15623 16819 15629
rect 16761 15589 16773 15623
rect 16807 15589 16819 15623
rect 16761 15583 16819 15589
rect 16206 15552 16212 15564
rect 16167 15524 16212 15552
rect 16206 15512 16212 15524
rect 16264 15512 16270 15564
rect 16390 15484 16396 15496
rect 16351 15456 16396 15484
rect 16390 15444 16396 15456
rect 16448 15444 16454 15496
rect 16776 15484 16804 15583
rect 17221 15487 17279 15493
rect 17221 15484 17233 15487
rect 16776 15456 17233 15484
rect 17221 15453 17233 15456
rect 17267 15453 17279 15487
rect 17221 15447 17279 15453
rect 17420 15388 26234 15416
rect 16114 15308 16120 15360
rect 16172 15348 16178 15360
rect 17420 15357 17448 15388
rect 16301 15351 16359 15357
rect 16301 15348 16313 15351
rect 16172 15320 16313 15348
rect 16172 15308 16178 15320
rect 16301 15317 16313 15320
rect 16347 15317 16359 15351
rect 16301 15311 16359 15317
rect 17405 15351 17463 15357
rect 17405 15317 17417 15351
rect 17451 15317 17463 15351
rect 26206 15348 26234 15388
rect 37274 15348 37280 15360
rect 26206 15320 37280 15348
rect 17405 15311 17463 15317
rect 37274 15308 37280 15320
rect 37332 15308 37338 15360
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 15746 15144 15752 15156
rect 15707 15116 15752 15144
rect 15746 15104 15752 15116
rect 15804 15104 15810 15156
rect 16390 15104 16396 15156
rect 16448 15144 16454 15156
rect 17313 15147 17371 15153
rect 17313 15144 17325 15147
rect 16448 15116 17325 15144
rect 16448 15104 16454 15116
rect 17313 15113 17325 15116
rect 17359 15113 17371 15147
rect 17313 15107 17371 15113
rect 15378 14968 15384 15020
rect 15436 15008 15442 15020
rect 15657 15011 15715 15017
rect 15657 15008 15669 15011
rect 15436 14980 15669 15008
rect 15436 14968 15442 14980
rect 15657 14977 15669 14980
rect 15703 14977 15715 15011
rect 16669 15011 16727 15017
rect 16669 15008 16681 15011
rect 15657 14971 15715 14977
rect 16546 14980 16681 15008
rect 15194 14900 15200 14952
rect 15252 14940 15258 14952
rect 15565 14943 15623 14949
rect 15565 14940 15577 14943
rect 15252 14912 15577 14940
rect 15252 14900 15258 14912
rect 15565 14909 15577 14912
rect 15611 14940 15623 14943
rect 16206 14940 16212 14952
rect 15611 14912 16212 14940
rect 15611 14909 15623 14912
rect 15565 14903 15623 14909
rect 16206 14900 16212 14912
rect 16264 14900 16270 14952
rect 16117 14875 16175 14881
rect 16117 14841 16129 14875
rect 16163 14872 16175 14875
rect 16546 14872 16574 14980
rect 16669 14977 16681 14980
rect 16715 14977 16727 15011
rect 37829 15011 37887 15017
rect 37829 15008 37841 15011
rect 16669 14971 16727 14977
rect 37292 14980 37841 15008
rect 16163 14844 16574 14872
rect 16853 14875 16911 14881
rect 16163 14841 16175 14844
rect 16117 14835 16175 14841
rect 16853 14841 16865 14875
rect 16899 14872 16911 14875
rect 16899 14844 26234 14872
rect 16899 14841 16911 14844
rect 16853 14835 16911 14841
rect 26206 14804 26234 14844
rect 37292 14813 37320 14980
rect 37829 14977 37841 14980
rect 37875 14977 37887 15011
rect 37829 14971 37887 14977
rect 38010 14872 38016 14884
rect 37971 14844 38016 14872
rect 38010 14832 38016 14844
rect 38068 14832 38074 14884
rect 37277 14807 37335 14813
rect 37277 14804 37289 14807
rect 26206 14776 37289 14804
rect 37277 14773 37289 14776
rect 37323 14773 37335 14807
rect 37277 14767 37335 14773
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 15746 14560 15752 14612
rect 15804 14600 15810 14612
rect 16485 14603 16543 14609
rect 16485 14600 16497 14603
rect 15804 14572 16497 14600
rect 15804 14560 15810 14572
rect 16485 14569 16497 14572
rect 16531 14569 16543 14603
rect 16485 14563 16543 14569
rect 15381 14535 15439 14541
rect 15381 14501 15393 14535
rect 15427 14501 15439 14535
rect 15381 14495 15439 14501
rect 14829 14467 14887 14473
rect 14829 14433 14841 14467
rect 14875 14464 14887 14467
rect 15194 14464 15200 14476
rect 14875 14436 15200 14464
rect 14875 14433 14887 14436
rect 14829 14427 14887 14433
rect 15194 14424 15200 14436
rect 15252 14424 15258 14476
rect 15010 14396 15016 14408
rect 14971 14368 15016 14396
rect 15010 14356 15016 14368
rect 15068 14356 15074 14408
rect 15396 14396 15424 14495
rect 15841 14399 15899 14405
rect 15841 14396 15853 14399
rect 15396 14368 15853 14396
rect 15841 14365 15853 14368
rect 15887 14365 15899 14399
rect 37829 14399 37887 14405
rect 37829 14396 37841 14399
rect 15841 14359 15899 14365
rect 37292 14368 37841 14396
rect 16040 14300 16574 14328
rect 14826 14220 14832 14272
rect 14884 14260 14890 14272
rect 16040 14269 16068 14300
rect 14921 14263 14979 14269
rect 14921 14260 14933 14263
rect 14884 14232 14933 14260
rect 14884 14220 14890 14232
rect 14921 14229 14933 14232
rect 14967 14229 14979 14263
rect 14921 14223 14979 14229
rect 16025 14263 16083 14269
rect 16025 14229 16037 14263
rect 16071 14229 16083 14263
rect 16546 14260 16574 14300
rect 37292 14269 37320 14368
rect 37829 14365 37841 14368
rect 37875 14365 37887 14399
rect 37829 14359 37887 14365
rect 37277 14263 37335 14269
rect 37277 14260 37289 14263
rect 16546 14232 37289 14260
rect 16025 14223 16083 14229
rect 37277 14229 37289 14232
rect 37323 14229 37335 14263
rect 38010 14260 38016 14272
rect 37971 14232 38016 14260
rect 37277 14223 37335 14229
rect 38010 14220 38016 14232
rect 38068 14220 38074 14272
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 14918 14056 14924 14068
rect 14879 14028 14924 14056
rect 14918 14016 14924 14028
rect 14976 14016 14982 14068
rect 15010 14016 15016 14068
rect 15068 14056 15074 14068
rect 15473 14059 15531 14065
rect 15473 14056 15485 14059
rect 15068 14028 15485 14056
rect 15068 14016 15074 14028
rect 15473 14025 15485 14028
rect 15519 14025 15531 14059
rect 15473 14019 15531 14025
rect 12345 13923 12403 13929
rect 12345 13920 12357 13923
rect 6886 13892 12357 13920
rect 4706 13812 4712 13864
rect 4764 13852 4770 13864
rect 6886 13852 6914 13892
rect 12345 13889 12357 13892
rect 12391 13889 12403 13923
rect 12345 13883 12403 13889
rect 15470 13880 15476 13932
rect 15528 13920 15534 13932
rect 37277 13923 37335 13929
rect 37277 13920 37289 13923
rect 15528 13892 37289 13920
rect 15528 13880 15534 13892
rect 37277 13889 37289 13892
rect 37323 13920 37335 13923
rect 37829 13923 37887 13929
rect 37829 13920 37841 13923
rect 37323 13892 37841 13920
rect 37323 13889 37335 13892
rect 37277 13883 37335 13889
rect 37829 13889 37841 13892
rect 37875 13889 37887 13923
rect 37829 13883 37887 13889
rect 12066 13852 12072 13864
rect 4764 13824 6914 13852
rect 12027 13824 12072 13852
rect 4764 13812 4770 13824
rect 12066 13812 12072 13824
rect 12124 13812 12130 13864
rect 38010 13716 38016 13728
rect 37971 13688 38016 13716
rect 38010 13676 38016 13688
rect 38068 13676 38074 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 12066 13512 12072 13524
rect 12027 13484 12072 13512
rect 12066 13472 12072 13484
rect 12124 13472 12130 13524
rect 15470 13512 15476 13524
rect 15431 13484 15476 13512
rect 15470 13472 15476 13484
rect 15528 13472 15534 13524
rect 12253 13447 12311 13453
rect 12253 13413 12265 13447
rect 12299 13444 12311 13447
rect 12894 13444 12900 13456
rect 12299 13416 12900 13444
rect 12299 13413 12311 13416
rect 12253 13407 12311 13413
rect 12894 13404 12900 13416
rect 12952 13404 12958 13456
rect 15102 13444 15108 13456
rect 14292 13416 15108 13444
rect 12529 13379 12587 13385
rect 12529 13345 12541 13379
rect 12575 13376 12587 13379
rect 12618 13376 12624 13388
rect 12575 13348 12624 13376
rect 12575 13345 12587 13348
rect 12529 13339 12587 13345
rect 12618 13336 12624 13348
rect 12676 13336 12682 13388
rect 13354 13336 13360 13388
rect 13412 13376 13418 13388
rect 14292 13385 14320 13416
rect 15102 13404 15108 13416
rect 15160 13404 15166 13456
rect 14277 13379 14335 13385
rect 14277 13376 14289 13379
rect 13412 13348 14289 13376
rect 13412 13336 13418 13348
rect 14277 13345 14289 13348
rect 14323 13345 14335 13379
rect 14918 13376 14924 13388
rect 14277 13339 14335 13345
rect 14476 13348 14924 13376
rect 14476 13317 14504 13348
rect 14918 13336 14924 13348
rect 14976 13336 14982 13388
rect 14461 13311 14519 13317
rect 14461 13277 14473 13311
rect 14507 13277 14519 13311
rect 15289 13311 15347 13317
rect 15289 13308 15301 13311
rect 14461 13271 14519 13277
rect 14844 13280 15301 13308
rect 12894 13132 12900 13184
rect 12952 13172 12958 13184
rect 12989 13175 13047 13181
rect 12989 13172 13001 13175
rect 12952 13144 13001 13172
rect 12952 13132 12958 13144
rect 12989 13141 13001 13144
rect 13035 13141 13047 13175
rect 14366 13172 14372 13184
rect 14327 13144 14372 13172
rect 12989 13135 13047 13141
rect 14366 13132 14372 13144
rect 14424 13132 14430 13184
rect 14844 13181 14872 13280
rect 15289 13277 15301 13280
rect 15335 13277 15347 13311
rect 37829 13311 37887 13317
rect 37829 13308 37841 13311
rect 15289 13271 15347 13277
rect 37292 13280 37841 13308
rect 37292 13184 37320 13280
rect 37829 13277 37841 13280
rect 37875 13277 37887 13311
rect 37829 13271 37887 13277
rect 14829 13175 14887 13181
rect 14829 13141 14841 13175
rect 14875 13141 14887 13175
rect 37274 13172 37280 13184
rect 37235 13144 37280 13172
rect 14829 13135 14887 13141
rect 37274 13132 37280 13144
rect 37332 13132 37338 13184
rect 38010 13172 38016 13184
rect 37971 13144 38016 13172
rect 38010 13132 38016 13144
rect 38068 13132 38074 13184
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 12618 12968 12624 12980
rect 12579 12940 12624 12968
rect 12618 12928 12624 12940
rect 12676 12928 12682 12980
rect 13538 12968 13544 12980
rect 13499 12940 13544 12968
rect 13538 12928 13544 12940
rect 13596 12928 13602 12980
rect 13909 12971 13967 12977
rect 13909 12937 13921 12971
rect 13955 12937 13967 12971
rect 13909 12931 13967 12937
rect 13556 12832 13584 12928
rect 13924 12832 13952 12931
rect 14369 12835 14427 12841
rect 14369 12832 14381 12835
rect 13556 12804 13860 12832
rect 13924 12804 14381 12832
rect 13354 12764 13360 12776
rect 13315 12736 13360 12764
rect 13354 12724 13360 12736
rect 13412 12724 13418 12776
rect 13449 12767 13507 12773
rect 13449 12733 13461 12767
rect 13495 12764 13507 12767
rect 13630 12764 13636 12776
rect 13495 12736 13636 12764
rect 13495 12733 13507 12736
rect 13449 12727 13507 12733
rect 13630 12724 13636 12736
rect 13688 12724 13694 12776
rect 13832 12764 13860 12804
rect 14369 12801 14381 12804
rect 14415 12801 14427 12835
rect 14369 12795 14427 12801
rect 15013 12767 15071 12773
rect 15013 12764 15025 12767
rect 13832 12736 15025 12764
rect 15013 12733 15025 12736
rect 15059 12733 15071 12767
rect 15013 12727 15071 12733
rect 14553 12699 14611 12705
rect 14553 12665 14565 12699
rect 14599 12696 14611 12699
rect 14599 12668 16574 12696
rect 14599 12665 14611 12668
rect 14553 12659 14611 12665
rect 16546 12628 16574 12668
rect 37274 12628 37280 12640
rect 16546 12600 37280 12628
rect 37274 12588 37280 12600
rect 37332 12588 37338 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 13354 12356 13360 12368
rect 12820 12328 13360 12356
rect 12820 12300 12848 12328
rect 13354 12316 13360 12328
rect 13412 12316 13418 12368
rect 12802 12288 12808 12300
rect 12715 12260 12808 12288
rect 12802 12248 12808 12260
rect 12860 12248 12866 12300
rect 14737 12291 14795 12297
rect 14737 12288 14749 12291
rect 13004 12260 14749 12288
rect 13004 12232 13032 12260
rect 14737 12257 14749 12260
rect 14783 12257 14795 12291
rect 14737 12251 14795 12257
rect 12986 12220 12992 12232
rect 12947 12192 12992 12220
rect 12986 12180 12992 12192
rect 13044 12180 13050 12232
rect 14093 12223 14151 12229
rect 14093 12220 14105 12223
rect 13372 12192 14105 12220
rect 12897 12155 12955 12161
rect 12897 12121 12909 12155
rect 12943 12152 12955 12155
rect 13170 12152 13176 12164
rect 12943 12124 13176 12152
rect 12943 12121 12955 12124
rect 12897 12115 12955 12121
rect 13170 12112 13176 12124
rect 13228 12112 13234 12164
rect 13372 12093 13400 12192
rect 14093 12189 14105 12192
rect 14139 12189 14151 12223
rect 37829 12223 37887 12229
rect 37829 12220 37841 12223
rect 14093 12183 14151 12189
rect 37292 12192 37841 12220
rect 14292 12124 16574 12152
rect 14292 12093 14320 12124
rect 13357 12087 13415 12093
rect 13357 12053 13369 12087
rect 13403 12053 13415 12087
rect 13357 12047 13415 12053
rect 14277 12087 14335 12093
rect 14277 12053 14289 12087
rect 14323 12053 14335 12087
rect 16546 12084 16574 12124
rect 37292 12093 37320 12192
rect 37829 12189 37841 12192
rect 37875 12189 37887 12223
rect 37829 12183 37887 12189
rect 37277 12087 37335 12093
rect 37277 12084 37289 12087
rect 16546 12056 37289 12084
rect 14277 12047 14335 12053
rect 37277 12053 37289 12056
rect 37323 12053 37335 12087
rect 38010 12084 38016 12096
rect 37971 12056 38016 12084
rect 37277 12047 37335 12053
rect 38010 12044 38016 12056
rect 38068 12044 38074 12096
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 12158 11880 12164 11892
rect 12119 11852 12164 11880
rect 12158 11840 12164 11852
rect 12216 11880 12222 11892
rect 12989 11883 13047 11889
rect 12989 11880 13001 11883
rect 12216 11852 13001 11880
rect 12216 11840 12222 11852
rect 12989 11849 13001 11852
rect 13035 11849 13047 11883
rect 12989 11843 13047 11849
rect 13357 11883 13415 11889
rect 13357 11849 13369 11883
rect 13403 11849 13415 11883
rect 13357 11843 13415 11849
rect 13372 11744 13400 11843
rect 13817 11747 13875 11753
rect 13817 11744 13829 11747
rect 13372 11716 13829 11744
rect 13817 11713 13829 11716
rect 13863 11713 13875 11747
rect 37829 11747 37887 11753
rect 37829 11744 37841 11747
rect 13817 11707 13875 11713
rect 37292 11716 37841 11744
rect 12802 11676 12808 11688
rect 12763 11648 12808 11676
rect 12802 11636 12808 11648
rect 12860 11636 12866 11688
rect 12897 11679 12955 11685
rect 12897 11645 12909 11679
rect 12943 11676 12955 11679
rect 13078 11676 13084 11688
rect 12943 11648 13084 11676
rect 12943 11645 12955 11648
rect 12897 11639 12955 11645
rect 13078 11636 13084 11648
rect 13136 11636 13142 11688
rect 37292 11549 37320 11716
rect 37829 11713 37841 11716
rect 37875 11713 37887 11747
rect 37829 11707 37887 11713
rect 14001 11543 14059 11549
rect 14001 11509 14013 11543
rect 14047 11540 14059 11543
rect 37277 11543 37335 11549
rect 37277 11540 37289 11543
rect 14047 11512 37289 11540
rect 14047 11509 14059 11512
rect 14001 11503 14059 11509
rect 37277 11509 37289 11512
rect 37323 11509 37335 11543
rect 38010 11540 38016 11552
rect 37971 11512 38016 11540
rect 37277 11503 37335 11509
rect 38010 11500 38016 11512
rect 38068 11500 38074 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 11974 11336 11980 11348
rect 11935 11308 11980 11336
rect 11974 11296 11980 11308
rect 12032 11296 12038 11348
rect 12802 11228 12808 11280
rect 12860 11228 12866 11280
rect 13173 11271 13231 11277
rect 13173 11237 13185 11271
rect 13219 11237 13231 11271
rect 13173 11231 13231 11237
rect 14277 11271 14335 11277
rect 14277 11237 14289 11271
rect 14323 11268 14335 11271
rect 38010 11268 38016 11280
rect 14323 11240 16574 11268
rect 37971 11240 38016 11268
rect 14323 11237 14335 11240
rect 14277 11231 14335 11237
rect 12621 11203 12679 11209
rect 12621 11169 12633 11203
rect 12667 11200 12679 11203
rect 12820 11200 12848 11228
rect 12667 11172 12848 11200
rect 12667 11169 12679 11172
rect 12621 11163 12679 11169
rect 11974 11092 11980 11144
rect 12032 11132 12038 11144
rect 12805 11135 12863 11141
rect 12805 11132 12817 11135
rect 12032 11104 12817 11132
rect 12032 11092 12038 11104
rect 12805 11101 12817 11104
rect 12851 11101 12863 11135
rect 13188 11132 13216 11231
rect 14093 11135 14151 11141
rect 14093 11132 14105 11135
rect 13188 11104 14105 11132
rect 12805 11095 12863 11101
rect 14093 11101 14105 11104
rect 14139 11101 14151 11135
rect 16546 11132 16574 11240
rect 38010 11228 38016 11240
rect 38068 11228 38074 11280
rect 37277 11135 37335 11141
rect 37277 11132 37289 11135
rect 16546 11104 37289 11132
rect 14093 11095 14151 11101
rect 37277 11101 37289 11104
rect 37323 11132 37335 11135
rect 37829 11135 37887 11141
rect 37829 11132 37841 11135
rect 37323 11104 37841 11132
rect 37323 11101 37335 11104
rect 37277 11095 37335 11101
rect 37829 11101 37841 11104
rect 37875 11101 37887 11135
rect 37829 11095 37887 11101
rect 2682 11024 2688 11076
rect 2740 11064 2746 11076
rect 11330 11064 11336 11076
rect 2740 11036 11336 11064
rect 2740 11024 2746 11036
rect 11330 11024 11336 11036
rect 11388 11024 11394 11076
rect 12713 11067 12771 11073
rect 12713 11033 12725 11067
rect 12759 11064 12771 11067
rect 13262 11064 13268 11076
rect 12759 11036 13268 11064
rect 12759 11033 12771 11036
rect 12713 11027 12771 11033
rect 13262 11024 13268 11036
rect 13320 11024 13326 11076
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 10410 10792 10416 10804
rect 10371 10764 10416 10792
rect 10410 10752 10416 10764
rect 10468 10752 10474 10804
rect 11330 10752 11336 10804
rect 11388 10792 11394 10804
rect 11885 10795 11943 10801
rect 11885 10792 11897 10795
rect 11388 10764 11897 10792
rect 11388 10752 11394 10764
rect 11885 10761 11897 10764
rect 11931 10761 11943 10795
rect 20162 10792 20168 10804
rect 11885 10755 11943 10761
rect 16546 10764 20168 10792
rect 9861 10727 9919 10733
rect 9861 10693 9873 10727
rect 9907 10724 9919 10727
rect 10134 10724 10140 10736
rect 9907 10696 10140 10724
rect 9907 10693 9919 10696
rect 9861 10687 9919 10693
rect 10134 10684 10140 10696
rect 10192 10724 10198 10736
rect 16546 10724 16574 10764
rect 20162 10752 20168 10764
rect 20220 10752 20226 10804
rect 37918 10724 37924 10736
rect 10192 10696 16574 10724
rect 26206 10696 37924 10724
rect 10192 10684 10198 10696
rect 10502 10616 10508 10668
rect 10560 10656 10566 10668
rect 11793 10659 11851 10665
rect 11793 10656 11805 10659
rect 10560 10628 11805 10656
rect 10560 10616 10566 10628
rect 11793 10625 11805 10628
rect 11839 10625 11851 10659
rect 11793 10619 11851 10625
rect 12618 10616 12624 10668
rect 12676 10656 12682 10668
rect 12713 10659 12771 10665
rect 12713 10656 12725 10659
rect 12676 10628 12725 10656
rect 12676 10616 12682 10628
rect 12713 10625 12725 10628
rect 12759 10625 12771 10659
rect 12894 10656 12900 10668
rect 12807 10628 12900 10656
rect 12713 10619 12771 10625
rect 12894 10616 12900 10628
rect 12952 10616 12958 10668
rect 13081 10659 13139 10665
rect 13081 10625 13093 10659
rect 13127 10656 13139 10659
rect 13725 10659 13783 10665
rect 13725 10656 13737 10659
rect 13127 10628 13737 10656
rect 13127 10625 13139 10628
rect 13081 10619 13139 10625
rect 13725 10625 13737 10628
rect 13771 10625 13783 10659
rect 13725 10619 13783 10625
rect 10965 10591 11023 10597
rect 10965 10557 10977 10591
rect 11011 10588 11023 10591
rect 11701 10591 11759 10597
rect 11701 10588 11713 10591
rect 11011 10560 11713 10588
rect 11011 10557 11023 10560
rect 10965 10551 11023 10557
rect 11701 10557 11713 10560
rect 11747 10588 11759 10591
rect 12636 10588 12664 10616
rect 11747 10560 12664 10588
rect 12912 10588 12940 10616
rect 12912 10560 14320 10588
rect 11747 10557 11759 10560
rect 11701 10551 11759 10557
rect 14292 10529 14320 10560
rect 14277 10523 14335 10529
rect 14277 10489 14289 10523
rect 14323 10520 14335 10523
rect 14323 10492 16574 10520
rect 14323 10489 14335 10492
rect 14277 10483 14335 10489
rect 12253 10455 12311 10461
rect 12253 10421 12265 10455
rect 12299 10452 12311 10455
rect 12434 10452 12440 10464
rect 12299 10424 12440 10452
rect 12299 10421 12311 10424
rect 12253 10415 12311 10421
rect 12434 10412 12440 10424
rect 12492 10412 12498 10464
rect 13446 10412 13452 10464
rect 13504 10452 13510 10464
rect 13541 10455 13599 10461
rect 13541 10452 13553 10455
rect 13504 10424 13553 10452
rect 13504 10412 13510 10424
rect 13541 10421 13553 10424
rect 13587 10421 13599 10455
rect 13541 10415 13599 10421
rect 13722 10412 13728 10464
rect 13780 10452 13786 10464
rect 14737 10455 14795 10461
rect 14737 10452 14749 10455
rect 13780 10424 14749 10452
rect 13780 10412 13786 10424
rect 14737 10421 14749 10424
rect 14783 10421 14795 10455
rect 16546 10452 16574 10492
rect 26206 10452 26234 10696
rect 37918 10684 37924 10696
rect 37976 10684 37982 10736
rect 37829 10659 37887 10665
rect 37829 10656 37841 10659
rect 37292 10628 37841 10656
rect 37292 10464 37320 10628
rect 37829 10625 37841 10628
rect 37875 10625 37887 10659
rect 37829 10619 37887 10625
rect 37274 10452 37280 10464
rect 16546 10424 26234 10452
rect 37235 10424 37280 10452
rect 14737 10415 14795 10421
rect 37274 10412 37280 10424
rect 37332 10412 37338 10464
rect 38010 10452 38016 10464
rect 37971 10424 38016 10452
rect 38010 10412 38016 10424
rect 38068 10412 38074 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 10781 10183 10839 10189
rect 10781 10149 10793 10183
rect 10827 10180 10839 10183
rect 10827 10152 11284 10180
rect 10827 10149 10839 10152
rect 10781 10143 10839 10149
rect 9585 10115 9643 10121
rect 9585 10081 9597 10115
rect 9631 10112 9643 10115
rect 10134 10112 10140 10124
rect 9631 10084 10140 10112
rect 9631 10081 9643 10084
rect 9585 10075 9643 10081
rect 10134 10072 10140 10084
rect 10192 10072 10198 10124
rect 11256 10121 11284 10152
rect 11241 10115 11299 10121
rect 11241 10081 11253 10115
rect 11287 10081 11299 10115
rect 11241 10075 11299 10081
rect 12618 10072 12624 10124
rect 12676 10112 12682 10124
rect 13081 10115 13139 10121
rect 13081 10112 13093 10115
rect 12676 10084 13093 10112
rect 12676 10072 12682 10084
rect 13081 10081 13093 10084
rect 13127 10112 13139 10115
rect 13722 10112 13728 10124
rect 13127 10084 13728 10112
rect 13127 10081 13139 10084
rect 13081 10075 13139 10081
rect 13722 10072 13728 10084
rect 13780 10112 13786 10124
rect 14093 10115 14151 10121
rect 14093 10112 14105 10115
rect 13780 10084 14105 10112
rect 13780 10072 13786 10084
rect 14093 10081 14105 10084
rect 14139 10081 14151 10115
rect 14093 10075 14151 10081
rect 10410 10044 10416 10056
rect 10371 10016 10416 10044
rect 10410 10004 10416 10016
rect 10468 10004 10474 10056
rect 11517 10047 11575 10053
rect 11517 10013 11529 10047
rect 11563 10044 11575 10047
rect 37274 10044 37280 10056
rect 11563 10016 37280 10044
rect 11563 10013 11575 10016
rect 11517 10007 11575 10013
rect 37274 10004 37280 10016
rect 37332 10004 37338 10056
rect 3418 9936 3424 9988
rect 3476 9976 3482 9988
rect 11974 9976 11980 9988
rect 3476 9948 11980 9976
rect 3476 9936 3482 9948
rect 11974 9936 11980 9948
rect 12032 9976 12038 9988
rect 12897 9979 12955 9985
rect 12897 9976 12909 9979
rect 12032 9948 12909 9976
rect 12032 9936 12038 9948
rect 12897 9945 12909 9948
rect 12943 9945 12955 9979
rect 12897 9939 12955 9945
rect 10318 9908 10324 9920
rect 10279 9880 10324 9908
rect 10318 9868 10324 9880
rect 10376 9868 10382 9920
rect 12526 9908 12532 9920
rect 12487 9880 12532 9908
rect 12526 9868 12532 9880
rect 12584 9868 12590 9920
rect 12986 9868 12992 9920
rect 13044 9908 13050 9920
rect 13044 9880 13089 9908
rect 13044 9868 13050 9880
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 9309 9639 9367 9645
rect 9309 9605 9321 9639
rect 9355 9636 9367 9639
rect 10042 9636 10048 9648
rect 9355 9608 10048 9636
rect 9355 9605 9367 9608
rect 9309 9599 9367 9605
rect 10042 9596 10048 9608
rect 10100 9596 10106 9648
rect 10134 9596 10140 9648
rect 10192 9596 10198 9648
rect 11974 9636 11980 9648
rect 11935 9608 11980 9636
rect 11974 9596 11980 9608
rect 12032 9596 12038 9648
rect 10152 9568 10180 9596
rect 9140 9540 10180 9568
rect 8202 9460 8208 9512
rect 8260 9500 8266 9512
rect 9140 9509 9168 9540
rect 12434 9528 12440 9580
rect 12492 9568 12498 9580
rect 12529 9571 12587 9577
rect 12529 9568 12541 9571
rect 12492 9540 12541 9568
rect 12492 9528 12498 9540
rect 12529 9537 12541 9540
rect 12575 9537 12587 9571
rect 37829 9571 37887 9577
rect 37829 9568 37841 9571
rect 12529 9531 12587 9537
rect 37292 9540 37841 9568
rect 9125 9503 9183 9509
rect 9125 9500 9137 9503
rect 8260 9472 9137 9500
rect 8260 9460 8266 9472
rect 9125 9469 9137 9472
rect 9171 9469 9183 9503
rect 9125 9463 9183 9469
rect 9217 9503 9275 9509
rect 9217 9469 9229 9503
rect 9263 9500 9275 9503
rect 9490 9500 9496 9512
rect 9263 9472 9496 9500
rect 9263 9469 9275 9472
rect 9217 9463 9275 9469
rect 9490 9460 9496 9472
rect 9548 9460 9554 9512
rect 10137 9503 10195 9509
rect 10137 9469 10149 9503
rect 10183 9469 10195 9503
rect 10137 9463 10195 9469
rect 10413 9503 10471 9509
rect 10413 9469 10425 9503
rect 10459 9469 10471 9503
rect 12802 9500 12808 9512
rect 12763 9472 12808 9500
rect 10413 9463 10471 9469
rect 9677 9435 9735 9441
rect 9677 9401 9689 9435
rect 9723 9432 9735 9435
rect 10152 9432 10180 9463
rect 9723 9404 10180 9432
rect 10428 9432 10456 9463
rect 12802 9460 12808 9472
rect 12860 9460 12866 9512
rect 37292 9441 37320 9540
rect 37829 9537 37841 9540
rect 37875 9537 37887 9571
rect 37829 9531 37887 9537
rect 37277 9435 37335 9441
rect 37277 9432 37289 9435
rect 10428 9404 37289 9432
rect 9723 9401 9735 9404
rect 9677 9395 9735 9401
rect 37277 9401 37289 9404
rect 37323 9401 37335 9435
rect 38010 9432 38016 9444
rect 37971 9404 38016 9432
rect 37277 9395 37335 9401
rect 38010 9392 38016 9404
rect 38068 9392 38074 9444
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 9585 9163 9643 9169
rect 9585 9129 9597 9163
rect 9631 9160 9643 9163
rect 10042 9160 10048 9172
rect 9631 9132 10048 9160
rect 9631 9129 9643 9132
rect 9585 9123 9643 9129
rect 10042 9120 10048 9132
rect 10100 9120 10106 9172
rect 12526 8984 12532 9036
rect 12584 9024 12590 9036
rect 12621 9027 12679 9033
rect 12621 9024 12633 9027
rect 12584 8996 12633 9024
rect 12584 8984 12590 8996
rect 12621 8993 12633 8996
rect 12667 8993 12679 9027
rect 12621 8987 12679 8993
rect 9582 8916 9588 8968
rect 9640 8956 9646 8968
rect 10045 8959 10103 8965
rect 10045 8956 10057 8959
rect 9640 8928 10057 8956
rect 9640 8916 9646 8928
rect 10045 8925 10057 8928
rect 10091 8925 10103 8959
rect 10045 8919 10103 8925
rect 10321 8959 10379 8965
rect 10321 8925 10333 8959
rect 10367 8925 10379 8959
rect 12342 8956 12348 8968
rect 12303 8928 12348 8956
rect 10321 8919 10379 8925
rect 10336 8888 10364 8919
rect 12342 8916 12348 8928
rect 12400 8916 12406 8968
rect 37829 8959 37887 8965
rect 37829 8925 37841 8959
rect 37875 8925 37887 8959
rect 37829 8919 37887 8925
rect 37277 8891 37335 8897
rect 37277 8888 37289 8891
rect 10336 8860 37289 8888
rect 37277 8857 37289 8860
rect 37323 8888 37335 8891
rect 37844 8888 37872 8919
rect 37323 8860 37872 8888
rect 37323 8857 37335 8860
rect 37277 8851 37335 8857
rect 38010 8820 38016 8832
rect 37971 8792 38016 8820
rect 38010 8780 38016 8792
rect 38068 8780 38074 8832
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 9214 8616 9220 8628
rect 9175 8588 9220 8616
rect 9214 8576 9220 8588
rect 9272 8576 9278 8628
rect 9582 8616 9588 8628
rect 9543 8588 9588 8616
rect 9582 8576 9588 8588
rect 9640 8576 9646 8628
rect 9232 8548 9260 8576
rect 10045 8551 10103 8557
rect 10045 8548 10057 8551
rect 9232 8520 10057 8548
rect 10045 8517 10057 8520
rect 10091 8517 10103 8551
rect 10045 8511 10103 8517
rect 37829 8483 37887 8489
rect 37829 8449 37841 8483
rect 37875 8449 37887 8483
rect 37829 8443 37887 8449
rect 8202 8372 8208 8424
rect 8260 8412 8266 8424
rect 8389 8415 8447 8421
rect 8389 8412 8401 8415
rect 8260 8384 8401 8412
rect 8260 8372 8266 8384
rect 8389 8381 8401 8384
rect 8435 8412 8447 8415
rect 8941 8415 8999 8421
rect 8941 8412 8953 8415
rect 8435 8384 8953 8412
rect 8435 8381 8447 8384
rect 8389 8375 8447 8381
rect 8941 8381 8953 8384
rect 8987 8381 8999 8415
rect 9122 8412 9128 8424
rect 9083 8384 9128 8412
rect 8941 8375 8999 8381
rect 9122 8372 9128 8384
rect 9180 8372 9186 8424
rect 9766 8372 9772 8424
rect 9824 8412 9830 8424
rect 37277 8415 37335 8421
rect 37277 8412 37289 8415
rect 9824 8384 37289 8412
rect 9824 8372 9830 8384
rect 37277 8381 37289 8384
rect 37323 8412 37335 8415
rect 37844 8412 37872 8443
rect 37323 8384 37872 8412
rect 37323 8381 37335 8384
rect 37277 8375 37335 8381
rect 9950 8304 9956 8356
rect 10008 8344 10014 8356
rect 10597 8347 10655 8353
rect 10597 8344 10609 8347
rect 10008 8316 10609 8344
rect 10008 8304 10014 8316
rect 10597 8313 10609 8316
rect 10643 8313 10655 8347
rect 38010 8344 38016 8356
rect 37971 8316 38016 8344
rect 10597 8307 10655 8313
rect 38010 8304 38016 8316
rect 38068 8304 38074 8356
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 8938 8072 8944 8084
rect 8899 8044 8944 8072
rect 8938 8032 8944 8044
rect 8996 8032 9002 8084
rect 8389 8007 8447 8013
rect 8389 7973 8401 8007
rect 8435 8004 8447 8007
rect 8435 7976 9536 8004
rect 8435 7973 8447 7976
rect 8389 7967 8447 7973
rect 7837 7939 7895 7945
rect 7837 7905 7849 7939
rect 7883 7936 7895 7939
rect 8202 7936 8208 7948
rect 7883 7908 8208 7936
rect 7883 7905 7895 7908
rect 7837 7899 7895 7905
rect 8202 7896 8208 7908
rect 8260 7896 8266 7948
rect 9508 7945 9536 7976
rect 9493 7939 9551 7945
rect 9493 7905 9505 7939
rect 9539 7905 9551 7939
rect 9766 7936 9772 7948
rect 9727 7908 9772 7936
rect 9493 7899 9551 7905
rect 9766 7896 9772 7908
rect 9824 7896 9830 7948
rect 8021 7871 8079 7877
rect 8021 7837 8033 7871
rect 8067 7868 8079 7871
rect 8938 7868 8944 7880
rect 8067 7840 8944 7868
rect 8067 7837 8079 7840
rect 8021 7831 8079 7837
rect 8938 7828 8944 7840
rect 8996 7828 9002 7880
rect 37829 7871 37887 7877
rect 37829 7868 37841 7871
rect 37292 7840 37841 7868
rect 37292 7744 37320 7840
rect 37829 7837 37841 7840
rect 37875 7837 37887 7871
rect 37829 7831 37887 7837
rect 7926 7732 7932 7744
rect 7887 7704 7932 7732
rect 7926 7692 7932 7704
rect 7984 7692 7990 7744
rect 37274 7732 37280 7744
rect 37235 7704 37280 7732
rect 37274 7692 37280 7704
rect 37332 7692 37338 7744
rect 38010 7732 38016 7744
rect 37971 7704 38016 7732
rect 38010 7692 38016 7704
rect 38068 7692 38074 7744
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 8018 7488 8024 7540
rect 8076 7528 8082 7540
rect 8205 7531 8263 7537
rect 8205 7528 8217 7531
rect 8076 7500 8217 7528
rect 8076 7488 8082 7500
rect 8205 7497 8217 7500
rect 8251 7528 8263 7531
rect 10413 7531 10471 7537
rect 10413 7528 10425 7531
rect 8251 7500 10425 7528
rect 8251 7497 8263 7500
rect 8205 7491 8263 7497
rect 10413 7497 10425 7500
rect 10459 7497 10471 7531
rect 10413 7491 10471 7497
rect 8202 7392 8208 7404
rect 7944 7364 8208 7392
rect 7377 7327 7435 7333
rect 7377 7293 7389 7327
rect 7423 7324 7435 7327
rect 7834 7324 7840 7336
rect 7423 7296 7840 7324
rect 7423 7293 7435 7296
rect 7377 7287 7435 7293
rect 7834 7284 7840 7296
rect 7892 7324 7898 7336
rect 7944 7333 7972 7364
rect 8202 7352 8208 7364
rect 8260 7352 8266 7404
rect 7929 7327 7987 7333
rect 7929 7324 7941 7327
rect 7892 7296 7941 7324
rect 7892 7284 7898 7296
rect 7929 7293 7941 7296
rect 7975 7293 7987 7327
rect 8110 7324 8116 7336
rect 8071 7296 8116 7324
rect 7929 7287 7987 7293
rect 8110 7284 8116 7296
rect 8168 7284 8174 7336
rect 9125 7327 9183 7333
rect 9125 7293 9137 7327
rect 9171 7293 9183 7327
rect 9125 7287 9183 7293
rect 9401 7327 9459 7333
rect 9401 7293 9413 7327
rect 9447 7324 9459 7327
rect 37274 7324 37280 7336
rect 9447 7296 37280 7324
rect 9447 7293 9459 7296
rect 9401 7287 9459 7293
rect 8573 7259 8631 7265
rect 8573 7225 8585 7259
rect 8619 7256 8631 7259
rect 9140 7256 9168 7287
rect 37274 7284 37280 7296
rect 37332 7284 37338 7336
rect 8619 7228 9168 7256
rect 8619 7225 8631 7228
rect 8573 7219 8631 7225
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 6546 6848 6552 6860
rect 6507 6820 6552 6848
rect 6546 6808 6552 6820
rect 6604 6848 6610 6860
rect 7193 6851 7251 6857
rect 6604 6820 6914 6848
rect 6604 6808 6610 6820
rect 6886 6780 6914 6820
rect 7193 6817 7205 6851
rect 7239 6848 7251 6851
rect 7834 6848 7840 6860
rect 7239 6820 7840 6848
rect 7239 6817 7251 6820
rect 7193 6811 7251 6817
rect 7834 6808 7840 6820
rect 7892 6808 7898 6860
rect 9217 6851 9275 6857
rect 9217 6817 9229 6851
rect 9263 6848 9275 6851
rect 9263 6820 16574 6848
rect 9263 6817 9275 6820
rect 9217 6811 9275 6817
rect 8021 6783 8079 6789
rect 8021 6780 8033 6783
rect 6886 6752 8033 6780
rect 8021 6749 8033 6752
rect 8067 6749 8079 6783
rect 8938 6780 8944 6792
rect 8899 6752 8944 6780
rect 8021 6743 8079 6749
rect 8938 6740 8944 6752
rect 8996 6740 9002 6792
rect 10226 6780 10232 6792
rect 10187 6752 10232 6780
rect 10226 6740 10232 6752
rect 10284 6740 10290 6792
rect 10505 6783 10563 6789
rect 10505 6749 10517 6783
rect 10551 6749 10563 6783
rect 16546 6780 16574 6820
rect 37277 6783 37335 6789
rect 37277 6780 37289 6783
rect 16546 6752 37289 6780
rect 10505 6743 10563 6749
rect 37277 6749 37289 6752
rect 37323 6780 37335 6783
rect 37829 6783 37887 6789
rect 37829 6780 37841 6783
rect 37323 6752 37841 6780
rect 37323 6749 37335 6752
rect 37277 6743 37335 6749
rect 37829 6749 37841 6752
rect 37875 6749 37887 6783
rect 37829 6743 37887 6749
rect 5166 6672 5172 6724
rect 5224 6712 5230 6724
rect 7929 6715 7987 6721
rect 7929 6712 7941 6715
rect 5224 6684 7941 6712
rect 5224 6672 5230 6684
rect 7929 6681 7941 6684
rect 7975 6681 7987 6715
rect 10520 6712 10548 6743
rect 37182 6712 37188 6724
rect 10520 6684 37188 6712
rect 7929 6675 7987 6681
rect 37182 6672 37188 6684
rect 37240 6672 37246 6724
rect 8386 6644 8392 6656
rect 8347 6616 8392 6644
rect 8386 6604 8392 6616
rect 8444 6604 8450 6656
rect 38010 6644 38016 6656
rect 37971 6616 38016 6644
rect 38010 6604 38016 6616
rect 38068 6604 38074 6656
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 7098 6440 7104 6452
rect 7059 6412 7104 6440
rect 7098 6400 7104 6412
rect 7156 6440 7162 6452
rect 8021 6443 8079 6449
rect 8021 6440 8033 6443
rect 7156 6412 8033 6440
rect 7156 6400 7162 6412
rect 8021 6409 8033 6412
rect 8067 6409 8079 6443
rect 8021 6403 8079 6409
rect 8389 6443 8447 6449
rect 8389 6409 8401 6443
rect 8435 6440 8447 6443
rect 8938 6440 8944 6452
rect 8435 6412 8944 6440
rect 8435 6409 8447 6412
rect 8389 6403 8447 6409
rect 8938 6400 8944 6412
rect 8996 6400 9002 6452
rect 9950 6400 9956 6452
rect 10008 6440 10014 6452
rect 10137 6443 10195 6449
rect 10137 6440 10149 6443
rect 10008 6412 10149 6440
rect 10008 6400 10014 6412
rect 10137 6409 10149 6412
rect 10183 6409 10195 6443
rect 10137 6403 10195 6409
rect 37182 6400 37188 6452
rect 37240 6440 37246 6452
rect 37277 6443 37335 6449
rect 37277 6440 37289 6443
rect 37240 6412 37289 6440
rect 37240 6400 37246 6412
rect 37277 6409 37289 6412
rect 37323 6409 37335 6443
rect 37277 6403 37335 6409
rect 7006 6264 7012 6316
rect 7064 6304 7070 6316
rect 7929 6307 7987 6313
rect 7929 6304 7941 6307
rect 7064 6276 7941 6304
rect 7064 6264 7070 6276
rect 7929 6273 7941 6276
rect 7975 6273 7987 6307
rect 7929 6267 7987 6273
rect 8386 6264 8392 6316
rect 8444 6304 8450 6316
rect 8849 6307 8907 6313
rect 8849 6304 8861 6307
rect 8444 6276 8861 6304
rect 8444 6264 8450 6276
rect 8849 6273 8861 6276
rect 8895 6273 8907 6307
rect 37292 6304 37320 6403
rect 37829 6307 37887 6313
rect 37829 6304 37841 6307
rect 37292 6276 37841 6304
rect 8849 6267 8907 6273
rect 37829 6273 37841 6276
rect 37875 6273 37887 6307
rect 37829 6267 37887 6273
rect 7742 6236 7748 6248
rect 7703 6208 7748 6236
rect 7742 6196 7748 6208
rect 7800 6196 7806 6248
rect 9125 6239 9183 6245
rect 9125 6205 9137 6239
rect 9171 6236 9183 6239
rect 37274 6236 37280 6248
rect 9171 6208 37280 6236
rect 9171 6205 9183 6208
rect 9125 6199 9183 6205
rect 37274 6196 37280 6208
rect 37332 6196 37338 6248
rect 38010 6100 38016 6112
rect 37971 6072 38016 6100
rect 38010 6060 38016 6072
rect 38068 6060 38074 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 6362 5856 6368 5908
rect 6420 5896 6426 5908
rect 8297 5899 8355 5905
rect 6420 5868 6914 5896
rect 6420 5856 6426 5868
rect 6886 5692 6914 5868
rect 8297 5865 8309 5899
rect 8343 5896 8355 5899
rect 10226 5896 10232 5908
rect 8343 5868 10232 5896
rect 8343 5865 8355 5868
rect 8297 5859 8355 5865
rect 10226 5856 10232 5868
rect 10284 5856 10290 5908
rect 37274 5896 37280 5908
rect 37235 5868 37280 5896
rect 37274 5856 37280 5868
rect 37332 5856 37338 5908
rect 7742 5760 7748 5772
rect 7703 5732 7748 5760
rect 7742 5720 7748 5732
rect 7800 5720 7806 5772
rect 7101 5695 7159 5701
rect 7101 5692 7113 5695
rect 6886 5664 7113 5692
rect 7101 5661 7113 5664
rect 7147 5692 7159 5695
rect 7929 5695 7987 5701
rect 7929 5692 7941 5695
rect 7147 5664 7941 5692
rect 7147 5661 7159 5664
rect 7101 5655 7159 5661
rect 7929 5661 7941 5664
rect 7975 5661 7987 5695
rect 8938 5692 8944 5704
rect 8899 5664 8944 5692
rect 7929 5655 7987 5661
rect 8938 5652 8944 5664
rect 8996 5652 9002 5704
rect 9214 5692 9220 5704
rect 9175 5664 9220 5692
rect 9214 5652 9220 5664
rect 9272 5652 9278 5704
rect 37292 5692 37320 5856
rect 37829 5695 37887 5701
rect 37829 5692 37841 5695
rect 37292 5664 37841 5692
rect 37829 5661 37841 5664
rect 37875 5661 37887 5695
rect 37829 5655 37887 5661
rect 7834 5556 7840 5568
rect 7795 5528 7840 5556
rect 7834 5516 7840 5528
rect 7892 5516 7898 5568
rect 38010 5556 38016 5568
rect 37971 5528 38016 5556
rect 38010 5516 38016 5528
rect 38068 5516 38074 5568
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 4890 5312 4896 5364
rect 4948 5352 4954 5364
rect 8297 5355 8355 5361
rect 4948 5324 6914 5352
rect 4948 5312 4954 5324
rect 6886 5284 6914 5324
rect 8297 5321 8309 5355
rect 8343 5352 8355 5355
rect 8938 5352 8944 5364
rect 8343 5324 8944 5352
rect 8343 5321 8355 5324
rect 8297 5315 8355 5321
rect 8938 5312 8944 5324
rect 8996 5312 9002 5364
rect 9401 5355 9459 5361
rect 9401 5321 9413 5355
rect 9447 5352 9459 5355
rect 9950 5352 9956 5364
rect 9447 5324 9956 5352
rect 9447 5321 9459 5324
rect 9401 5315 9459 5321
rect 7101 5287 7159 5293
rect 7101 5284 7113 5287
rect 6886 5256 7113 5284
rect 7101 5253 7113 5256
rect 7147 5284 7159 5287
rect 7929 5287 7987 5293
rect 7929 5284 7941 5287
rect 7147 5256 7941 5284
rect 7147 5253 7159 5256
rect 7101 5247 7159 5253
rect 7929 5253 7941 5256
rect 7975 5253 7987 5287
rect 7929 5247 7987 5253
rect 8849 5287 8907 5293
rect 8849 5253 8861 5287
rect 8895 5284 8907 5287
rect 9416 5284 9444 5315
rect 9950 5312 9956 5324
rect 10008 5312 10014 5364
rect 8895 5256 9444 5284
rect 8895 5253 8907 5256
rect 8849 5247 8907 5253
rect 5534 5176 5540 5228
rect 5592 5216 5598 5228
rect 7837 5219 7895 5225
rect 7837 5216 7849 5219
rect 5592 5188 7849 5216
rect 5592 5176 5598 5188
rect 7837 5185 7849 5188
rect 7883 5185 7895 5219
rect 7837 5179 7895 5185
rect 7742 5148 7748 5160
rect 7655 5120 7748 5148
rect 7742 5108 7748 5120
rect 7800 5148 7806 5160
rect 8864 5148 8892 5247
rect 9214 5176 9220 5228
rect 9272 5216 9278 5228
rect 37277 5219 37335 5225
rect 37277 5216 37289 5219
rect 9272 5188 37289 5216
rect 9272 5176 9278 5188
rect 37277 5185 37289 5188
rect 37323 5216 37335 5219
rect 37829 5219 37887 5225
rect 37829 5216 37841 5219
rect 37323 5188 37841 5216
rect 37323 5185 37335 5188
rect 37277 5179 37335 5185
rect 37829 5185 37841 5188
rect 37875 5185 37887 5219
rect 37829 5179 37887 5185
rect 7800 5120 8892 5148
rect 7800 5108 7806 5120
rect 38010 5012 38016 5024
rect 37971 4984 38016 5012
rect 38010 4972 38016 4984
rect 38068 4972 38074 5024
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 36722 4428 36728 4480
rect 36780 4468 36786 4480
rect 36817 4471 36875 4477
rect 36817 4468 36829 4471
rect 36780 4440 36829 4468
rect 36780 4428 36786 4440
rect 36817 4437 36829 4440
rect 36863 4437 36875 4471
rect 36817 4431 36875 4437
rect 37553 4471 37611 4477
rect 37553 4437 37565 4471
rect 37599 4468 37611 4471
rect 37642 4468 37648 4480
rect 37599 4440 37648 4468
rect 37599 4437 37611 4440
rect 37553 4431 37611 4437
rect 37642 4428 37648 4440
rect 37700 4428 37706 4480
rect 38010 4468 38016 4480
rect 37971 4440 38016 4468
rect 38010 4428 38016 4440
rect 38068 4428 38074 4480
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 38010 4196 38016 4208
rect 37971 4168 38016 4196
rect 38010 4156 38016 4168
rect 38068 4156 38074 4208
rect 37829 4131 37887 4137
rect 37829 4097 37841 4131
rect 37875 4128 37887 4131
rect 37918 4128 37924 4140
rect 37875 4100 37924 4128
rect 37875 4097 37887 4100
rect 37829 4091 37887 4097
rect 37918 4088 37924 4100
rect 37976 4088 37982 4140
rect 12342 3952 12348 4004
rect 12400 3992 12406 4004
rect 37277 3995 37335 4001
rect 37277 3992 37289 3995
rect 12400 3964 37289 3992
rect 12400 3952 12406 3964
rect 37277 3961 37289 3964
rect 37323 3992 37335 3995
rect 37826 3992 37832 4004
rect 37323 3964 37832 3992
rect 37323 3961 37335 3964
rect 37277 3955 37335 3961
rect 37826 3952 37832 3964
rect 37884 3952 37890 4004
rect 34698 3924 34704 3936
rect 34659 3896 34704 3924
rect 34698 3884 34704 3896
rect 34756 3884 34762 3936
rect 36170 3924 36176 3936
rect 36131 3896 36176 3924
rect 36170 3884 36176 3896
rect 36228 3884 36234 3936
rect 36446 3884 36452 3936
rect 36504 3924 36510 3936
rect 36633 3927 36691 3933
rect 36633 3924 36645 3927
rect 36504 3896 36645 3924
rect 36504 3884 36510 3896
rect 36633 3893 36645 3896
rect 36679 3893 36691 3927
rect 36633 3887 36691 3893
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 34790 3612 34796 3664
rect 34848 3612 34854 3664
rect 34808 3584 34836 3612
rect 35069 3587 35127 3593
rect 35069 3584 35081 3587
rect 34808 3556 35081 3584
rect 35069 3553 35081 3556
rect 35115 3553 35127 3587
rect 36538 3584 36544 3596
rect 36499 3556 36544 3584
rect 35069 3547 35127 3553
rect 36538 3544 36544 3556
rect 36596 3544 36602 3596
rect 34698 3476 34704 3528
rect 34756 3516 34762 3528
rect 34793 3519 34851 3525
rect 34793 3516 34805 3519
rect 34756 3488 34805 3516
rect 34756 3476 34762 3488
rect 34793 3485 34805 3488
rect 34839 3485 34851 3519
rect 34793 3479 34851 3485
rect 36170 3476 36176 3528
rect 36228 3516 36234 3528
rect 36265 3519 36323 3525
rect 36265 3516 36277 3519
rect 36228 3488 36277 3516
rect 36228 3476 36234 3488
rect 36265 3485 36277 3488
rect 36311 3485 36323 3519
rect 37826 3516 37832 3528
rect 37787 3488 37832 3516
rect 36265 3479 36323 3485
rect 37826 3476 37832 3488
rect 37884 3476 37890 3528
rect 5258 3380 5264 3392
rect 5219 3352 5264 3380
rect 5258 3340 5264 3352
rect 5316 3340 5322 3392
rect 30282 3380 30288 3392
rect 30243 3352 30288 3380
rect 30282 3340 30288 3352
rect 30340 3340 30346 3392
rect 31754 3340 31760 3392
rect 31812 3380 31818 3392
rect 31941 3383 31999 3389
rect 31941 3380 31953 3383
rect 31812 3352 31953 3380
rect 31812 3340 31818 3352
rect 31941 3349 31953 3352
rect 31987 3349 31999 3383
rect 31941 3343 31999 3349
rect 33042 3340 33048 3392
rect 33100 3380 33106 3392
rect 33229 3383 33287 3389
rect 33229 3380 33241 3383
rect 33100 3352 33241 3380
rect 33100 3340 33106 3352
rect 33229 3349 33241 3352
rect 33275 3349 33287 3383
rect 38010 3380 38016 3392
rect 37971 3352 38016 3380
rect 33229 3343 33287 3349
rect 38010 3340 38016 3352
rect 38068 3340 38074 3392
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 4801 3179 4859 3185
rect 4801 3145 4813 3179
rect 4847 3176 4859 3179
rect 5534 3176 5540 3188
rect 4847 3148 5540 3176
rect 4847 3145 4859 3148
rect 4801 3139 4859 3145
rect 5534 3136 5540 3148
rect 5592 3136 5598 3188
rect 9122 3136 9128 3188
rect 9180 3176 9186 3188
rect 9217 3179 9275 3185
rect 9217 3176 9229 3179
rect 9180 3148 9229 3176
rect 9180 3136 9186 3148
rect 9217 3145 9229 3148
rect 9263 3145 9275 3179
rect 14366 3176 14372 3188
rect 14327 3148 14372 3176
rect 9217 3139 9275 3145
rect 14366 3136 14372 3148
rect 14424 3136 14430 3188
rect 22002 3176 22008 3188
rect 21963 3148 22008 3176
rect 22002 3136 22008 3148
rect 22060 3136 22066 3188
rect 22922 3136 22928 3188
rect 22980 3176 22986 3188
rect 23017 3179 23075 3185
rect 23017 3176 23029 3179
rect 22980 3148 23029 3176
rect 22980 3136 22986 3148
rect 23017 3145 23029 3148
rect 23063 3145 23075 3179
rect 23017 3139 23075 3145
rect 26050 3136 26056 3188
rect 26108 3176 26114 3188
rect 26145 3179 26203 3185
rect 26145 3176 26157 3179
rect 26108 3148 26157 3176
rect 26108 3136 26114 3148
rect 26145 3145 26157 3148
rect 26191 3145 26203 3179
rect 29086 3176 29092 3188
rect 29047 3148 29092 3176
rect 26145 3139 26203 3145
rect 29086 3136 29092 3148
rect 29144 3136 29150 3188
rect 36446 3176 36452 3188
rect 35866 3148 36452 3176
rect 12802 3068 12808 3120
rect 12860 3108 12866 3120
rect 35866 3108 35894 3148
rect 36446 3136 36452 3148
rect 36504 3136 36510 3188
rect 37734 3136 37740 3188
rect 37792 3176 37798 3188
rect 37921 3179 37979 3185
rect 37921 3176 37933 3179
rect 37792 3148 37933 3176
rect 37792 3136 37798 3148
rect 37921 3145 37933 3148
rect 37967 3145 37979 3179
rect 37921 3139 37979 3145
rect 12860 3080 35894 3108
rect 12860 3068 12866 3080
rect 4157 3043 4215 3049
rect 4157 3009 4169 3043
rect 4203 3040 4215 3043
rect 4614 3040 4620 3052
rect 4203 3012 4620 3040
rect 4203 3009 4215 3012
rect 4157 3003 4215 3009
rect 4614 3000 4620 3012
rect 4672 3000 4678 3052
rect 8573 3043 8631 3049
rect 8573 3009 8585 3043
rect 8619 3040 8631 3043
rect 8938 3040 8944 3052
rect 8619 3012 8944 3040
rect 8619 3009 8631 3012
rect 8573 3003 8631 3009
rect 8938 3000 8944 3012
rect 8996 3040 9002 3052
rect 9033 3043 9091 3049
rect 9033 3040 9045 3043
rect 8996 3012 9045 3040
rect 8996 3000 9002 3012
rect 9033 3009 9045 3012
rect 9079 3009 9091 3043
rect 9033 3003 9091 3009
rect 13725 3043 13783 3049
rect 13725 3009 13737 3043
rect 13771 3040 13783 3043
rect 14090 3040 14096 3052
rect 13771 3012 14096 3040
rect 13771 3009 13783 3012
rect 13725 3003 13783 3009
rect 14090 3000 14096 3012
rect 14148 3040 14154 3052
rect 14185 3043 14243 3049
rect 14185 3040 14197 3043
rect 14148 3012 14197 3040
rect 14148 3000 14154 3012
rect 14185 3009 14197 3012
rect 14231 3009 14243 3043
rect 14185 3003 14243 3009
rect 21450 3000 21456 3052
rect 21508 3040 21514 3052
rect 21821 3043 21879 3049
rect 21821 3040 21833 3043
rect 21508 3012 21833 3040
rect 21508 3000 21514 3012
rect 21821 3009 21833 3012
rect 21867 3040 21879 3043
rect 22465 3043 22523 3049
rect 22465 3040 22477 3043
rect 21867 3012 22477 3040
rect 21867 3009 21879 3012
rect 21821 3003 21879 3009
rect 22465 3009 22477 3012
rect 22511 3009 22523 3043
rect 22465 3003 22523 3009
rect 25501 3043 25559 3049
rect 25501 3009 25513 3043
rect 25547 3040 25559 3043
rect 25866 3040 25872 3052
rect 25547 3012 25872 3040
rect 25547 3009 25559 3012
rect 25501 3003 25559 3009
rect 25866 3000 25872 3012
rect 25924 3040 25930 3052
rect 25961 3043 26019 3049
rect 25961 3040 25973 3043
rect 25924 3012 25973 3040
rect 25924 3000 25930 3012
rect 25961 3009 25973 3012
rect 26007 3009 26019 3043
rect 25961 3003 26019 3009
rect 28810 3000 28816 3052
rect 28868 3040 28874 3052
rect 28905 3043 28963 3049
rect 28905 3040 28917 3043
rect 28868 3012 28917 3040
rect 28868 3000 28874 3012
rect 28905 3009 28917 3012
rect 28951 3040 28963 3043
rect 29549 3043 29607 3049
rect 29549 3040 29561 3043
rect 28951 3012 29561 3040
rect 28951 3009 28963 3012
rect 28905 3003 28963 3009
rect 29549 3009 29561 3012
rect 29595 3009 29607 3043
rect 30650 3040 30656 3052
rect 30611 3012 30656 3040
rect 29549 3003 29607 3009
rect 30650 3000 30656 3012
rect 30708 3000 30714 3052
rect 32398 3040 32404 3052
rect 32359 3012 32404 3040
rect 32398 3000 32404 3012
rect 32456 3000 32462 3052
rect 32582 3000 32588 3052
rect 32640 3040 32646 3052
rect 33689 3043 33747 3049
rect 33689 3040 33701 3043
rect 32640 3012 33701 3040
rect 32640 3000 32646 3012
rect 33689 3009 33701 3012
rect 33735 3009 33747 3043
rect 33689 3003 33747 3009
rect 34054 3000 34060 3052
rect 34112 3040 34118 3052
rect 34977 3043 35035 3049
rect 34977 3040 34989 3043
rect 34112 3012 34989 3040
rect 34112 3000 34118 3012
rect 34977 3009 34989 3012
rect 35023 3009 35035 3043
rect 36446 3040 36452 3052
rect 36407 3012 36452 3040
rect 34977 3003 35035 3009
rect 36446 3000 36452 3012
rect 36504 3000 36510 3052
rect 37642 3000 37648 3052
rect 37700 3040 37706 3052
rect 37829 3043 37887 3049
rect 37829 3040 37841 3043
rect 37700 3012 37841 3040
rect 37700 3000 37706 3012
rect 37829 3009 37841 3012
rect 37875 3009 37887 3043
rect 37829 3003 37887 3009
rect 30282 2932 30288 2984
rect 30340 2972 30346 2984
rect 30377 2975 30435 2981
rect 30377 2972 30389 2975
rect 30340 2944 30389 2972
rect 30340 2932 30346 2944
rect 30377 2941 30389 2944
rect 30423 2941 30435 2975
rect 30377 2935 30435 2941
rect 31754 2932 31760 2984
rect 31812 2972 31818 2984
rect 32125 2975 32183 2981
rect 32125 2972 32137 2975
rect 31812 2944 32137 2972
rect 31812 2932 31818 2944
rect 32125 2941 32137 2944
rect 32171 2941 32183 2975
rect 32125 2935 32183 2941
rect 32490 2932 32496 2984
rect 32548 2972 32554 2984
rect 33042 2972 33048 2984
rect 32548 2944 33048 2972
rect 32548 2932 32554 2944
rect 33042 2932 33048 2944
rect 33100 2972 33106 2984
rect 33413 2975 33471 2981
rect 33413 2972 33425 2975
rect 33100 2944 33425 2972
rect 33100 2932 33106 2944
rect 33413 2941 33425 2944
rect 33459 2941 33471 2975
rect 33413 2935 33471 2941
rect 33962 2932 33968 2984
rect 34020 2972 34026 2984
rect 34701 2975 34759 2981
rect 34701 2972 34713 2975
rect 34020 2944 34713 2972
rect 34020 2932 34026 2944
rect 34701 2941 34713 2944
rect 34747 2941 34759 2975
rect 34701 2935 34759 2941
rect 3050 2796 3056 2848
rect 3108 2836 3114 2848
rect 3329 2839 3387 2845
rect 3329 2836 3341 2839
rect 3108 2808 3341 2836
rect 3108 2796 3114 2808
rect 3329 2805 3341 2808
rect 3375 2805 3387 2839
rect 3329 2799 3387 2805
rect 5813 2839 5871 2845
rect 5813 2805 5825 2839
rect 5859 2836 5871 2839
rect 5994 2836 6000 2848
rect 5859 2808 6000 2836
rect 5859 2805 5871 2808
rect 5813 2799 5871 2805
rect 5994 2796 6000 2808
rect 6052 2796 6058 2848
rect 6730 2836 6736 2848
rect 6691 2808 6736 2836
rect 6730 2796 6736 2808
rect 6788 2796 6794 2848
rect 7466 2836 7472 2848
rect 7427 2808 7472 2836
rect 7466 2796 7472 2808
rect 7524 2796 7530 2848
rect 9674 2796 9680 2848
rect 9732 2836 9738 2848
rect 9769 2839 9827 2845
rect 9769 2836 9781 2839
rect 9732 2808 9781 2836
rect 9732 2796 9738 2808
rect 9769 2805 9781 2808
rect 9815 2805 9827 2839
rect 10410 2836 10416 2848
rect 10371 2808 10416 2836
rect 9769 2799 9827 2805
rect 10410 2796 10416 2808
rect 10468 2796 10474 2848
rect 10962 2836 10968 2848
rect 10923 2808 10968 2836
rect 10962 2796 10968 2808
rect 11020 2796 11026 2848
rect 11882 2836 11888 2848
rect 11843 2808 11888 2836
rect 11882 2796 11888 2808
rect 11940 2796 11946 2848
rect 12618 2836 12624 2848
rect 12579 2808 12624 2836
rect 12618 2796 12624 2808
rect 12676 2796 12682 2848
rect 14918 2836 14924 2848
rect 14879 2808 14924 2836
rect 14918 2796 14924 2808
rect 14976 2796 14982 2848
rect 15562 2836 15568 2848
rect 15523 2808 15568 2836
rect 15562 2796 15568 2808
rect 15620 2796 15626 2848
rect 16117 2839 16175 2845
rect 16117 2805 16129 2839
rect 16163 2836 16175 2839
rect 16298 2836 16304 2848
rect 16163 2808 16304 2836
rect 16163 2805 16175 2808
rect 16117 2799 16175 2805
rect 16298 2796 16304 2808
rect 16356 2796 16362 2848
rect 17034 2836 17040 2848
rect 16995 2808 17040 2836
rect 17034 2796 17040 2808
rect 17092 2796 17098 2848
rect 17770 2836 17776 2848
rect 17731 2808 17776 2836
rect 17770 2796 17776 2808
rect 17828 2796 17834 2848
rect 18598 2836 18604 2848
rect 18559 2808 18604 2836
rect 18598 2796 18604 2808
rect 18656 2796 18662 2848
rect 19242 2836 19248 2848
rect 19203 2808 19248 2836
rect 19242 2796 19248 2808
rect 19300 2796 19306 2848
rect 19978 2836 19984 2848
rect 19939 2808 19984 2836
rect 19978 2796 19984 2808
rect 20036 2796 20042 2848
rect 20717 2839 20775 2845
rect 20717 2805 20729 2839
rect 20763 2836 20775 2839
rect 20806 2836 20812 2848
rect 20763 2808 20812 2836
rect 20763 2805 20775 2808
rect 20717 2799 20775 2805
rect 20806 2796 20812 2808
rect 20864 2796 20870 2848
rect 24210 2836 24216 2848
rect 24171 2808 24216 2836
rect 24210 2796 24216 2808
rect 24268 2796 24274 2848
rect 24394 2796 24400 2848
rect 24452 2836 24458 2848
rect 24857 2839 24915 2845
rect 24857 2836 24869 2839
rect 24452 2808 24869 2836
rect 24452 2796 24458 2808
rect 24857 2805 24869 2808
rect 24903 2836 24915 2839
rect 25038 2836 25044 2848
rect 24903 2808 25044 2836
rect 24903 2805 24915 2808
rect 24857 2799 24915 2805
rect 25038 2796 25044 2808
rect 25096 2796 25102 2848
rect 26970 2836 26976 2848
rect 26931 2808 26976 2836
rect 26970 2796 26976 2808
rect 27028 2796 27034 2848
rect 27614 2836 27620 2848
rect 27575 2808 27620 2836
rect 27614 2796 27620 2808
rect 27672 2796 27678 2848
rect 33226 2796 33232 2848
rect 33284 2836 33290 2848
rect 34606 2836 34612 2848
rect 33284 2808 34612 2836
rect 33284 2796 33290 2808
rect 34606 2796 34612 2808
rect 34664 2796 34670 2848
rect 36630 2836 36636 2848
rect 36591 2808 36636 2836
rect 36630 2796 36636 2808
rect 36688 2796 36694 2848
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 5166 2632 5172 2644
rect 5127 2604 5172 2632
rect 5166 2592 5172 2604
rect 5224 2592 5230 2644
rect 5813 2635 5871 2641
rect 5813 2601 5825 2635
rect 5859 2632 5871 2635
rect 7834 2632 7840 2644
rect 5859 2604 7840 2632
rect 5859 2601 5871 2604
rect 5813 2595 5871 2601
rect 7834 2592 7840 2604
rect 7892 2592 7898 2644
rect 7926 2592 7932 2644
rect 7984 2632 7990 2644
rect 8205 2635 8263 2641
rect 8205 2632 8217 2635
rect 7984 2604 8217 2632
rect 7984 2592 7990 2604
rect 8205 2601 8217 2604
rect 8251 2601 8263 2635
rect 9490 2632 9496 2644
rect 9451 2604 9496 2632
rect 8205 2595 8263 2601
rect 9490 2592 9496 2604
rect 9548 2592 9554 2644
rect 10318 2632 10324 2644
rect 10279 2604 10324 2632
rect 10318 2592 10324 2604
rect 10376 2592 10382 2644
rect 12897 2635 12955 2641
rect 12897 2601 12909 2635
rect 12943 2632 12955 2635
rect 13170 2632 13176 2644
rect 12943 2604 13176 2632
rect 12943 2601 12955 2604
rect 12897 2595 12955 2601
rect 13170 2592 13176 2604
rect 13228 2592 13234 2644
rect 13541 2635 13599 2641
rect 13541 2601 13553 2635
rect 13587 2632 13599 2635
rect 13630 2632 13636 2644
rect 13587 2604 13636 2632
rect 13587 2601 13599 2604
rect 13541 2595 13599 2601
rect 13630 2592 13636 2604
rect 13688 2592 13694 2644
rect 14826 2632 14832 2644
rect 14787 2604 14832 2632
rect 14826 2592 14832 2604
rect 14884 2592 14890 2644
rect 15378 2592 15384 2644
rect 15436 2632 15442 2644
rect 15473 2635 15531 2641
rect 15473 2632 15485 2635
rect 15436 2604 15485 2632
rect 15436 2592 15442 2604
rect 15473 2601 15485 2604
rect 15519 2601 15531 2635
rect 16114 2632 16120 2644
rect 16075 2604 16120 2632
rect 15473 2595 15531 2601
rect 16114 2592 16120 2604
rect 16172 2592 16178 2644
rect 17310 2632 17316 2644
rect 17271 2604 17316 2632
rect 17310 2592 17316 2604
rect 17368 2592 17374 2644
rect 18049 2635 18107 2641
rect 18049 2601 18061 2635
rect 18095 2632 18107 2635
rect 18138 2632 18144 2644
rect 18095 2604 18144 2632
rect 18095 2601 18107 2604
rect 18049 2595 18107 2601
rect 18138 2592 18144 2604
rect 18196 2592 18202 2644
rect 18506 2632 18512 2644
rect 18467 2604 18512 2632
rect 18506 2592 18512 2604
rect 18564 2592 18570 2644
rect 20070 2632 20076 2644
rect 20031 2604 20076 2632
rect 20070 2592 20076 2604
rect 20128 2592 20134 2644
rect 20714 2592 20720 2644
rect 20772 2632 20778 2644
rect 20809 2635 20867 2641
rect 20809 2632 20821 2635
rect 20772 2604 20821 2632
rect 20772 2592 20778 2604
rect 20809 2601 20821 2604
rect 20855 2601 20867 2635
rect 20809 2595 20867 2601
rect 23201 2635 23259 2641
rect 23201 2601 23213 2635
rect 23247 2632 23259 2635
rect 23290 2632 23296 2644
rect 23247 2604 23296 2632
rect 23247 2601 23259 2604
rect 23201 2595 23259 2601
rect 23290 2592 23296 2604
rect 23348 2592 23354 2644
rect 24578 2632 24584 2644
rect 24539 2604 24584 2632
rect 24578 2592 24584 2604
rect 24636 2592 24642 2644
rect 25222 2632 25228 2644
rect 25183 2604 25228 2632
rect 25222 2592 25228 2604
rect 25280 2592 25286 2644
rect 25869 2635 25927 2641
rect 25869 2601 25881 2635
rect 25915 2632 25927 2635
rect 26234 2632 26240 2644
rect 25915 2604 26240 2632
rect 25915 2601 25927 2604
rect 25869 2595 25927 2601
rect 26234 2592 26240 2604
rect 26292 2592 26298 2644
rect 27154 2632 27160 2644
rect 27115 2604 27160 2632
rect 27154 2592 27160 2604
rect 27212 2592 27218 2644
rect 27798 2632 27804 2644
rect 27759 2604 27804 2632
rect 27798 2592 27804 2604
rect 27856 2592 27862 2644
rect 28442 2632 28448 2644
rect 28403 2604 28448 2632
rect 28442 2592 28448 2604
rect 28500 2592 28506 2644
rect 36538 2632 36544 2644
rect 36499 2604 36544 2632
rect 36538 2592 36544 2604
rect 36596 2592 36602 2644
rect 3237 2567 3295 2573
rect 3237 2533 3249 2567
rect 3283 2564 3295 2567
rect 3283 2536 4936 2564
rect 3283 2533 3295 2536
rect 3237 2527 3295 2533
rect 4908 2496 4936 2536
rect 5074 2524 5080 2576
rect 5132 2564 5138 2576
rect 6914 2564 6920 2576
rect 5132 2536 6920 2564
rect 5132 2524 5138 2536
rect 6914 2524 6920 2536
rect 6972 2524 6978 2576
rect 7006 2524 7012 2576
rect 7064 2564 7070 2576
rect 7745 2567 7803 2573
rect 7064 2536 7109 2564
rect 7064 2524 7070 2536
rect 7745 2533 7757 2567
rect 7791 2564 7803 2567
rect 8110 2564 8116 2576
rect 7791 2536 8116 2564
rect 7791 2533 7803 2536
rect 7745 2527 7803 2533
rect 8110 2524 8116 2536
rect 8168 2524 8174 2576
rect 12161 2567 12219 2573
rect 12161 2533 12173 2567
rect 12207 2564 12219 2567
rect 13078 2564 13084 2576
rect 12207 2536 13084 2564
rect 12207 2533 12219 2536
rect 12161 2527 12219 2533
rect 13078 2524 13084 2536
rect 13136 2524 13142 2576
rect 19521 2567 19579 2573
rect 19521 2533 19533 2567
rect 19567 2564 19579 2567
rect 20346 2564 20352 2576
rect 19567 2536 20352 2564
rect 19567 2533 19579 2536
rect 19521 2527 19579 2533
rect 20346 2524 20352 2536
rect 20404 2524 20410 2576
rect 33597 2567 33655 2573
rect 33597 2533 33609 2567
rect 33643 2564 33655 2567
rect 35434 2564 35440 2576
rect 33643 2536 35440 2564
rect 33643 2533 33655 2536
rect 33597 2527 33655 2533
rect 35434 2524 35440 2536
rect 35492 2564 35498 2576
rect 35492 2536 37320 2564
rect 35492 2524 35498 2536
rect 12986 2496 12992 2508
rect 4908 2468 12992 2496
rect 12986 2456 12992 2468
rect 13044 2456 13050 2508
rect 30193 2499 30251 2505
rect 30193 2465 30205 2499
rect 30239 2496 30251 2499
rect 30558 2496 30564 2508
rect 30239 2468 30564 2496
rect 30239 2465 30251 2468
rect 30193 2459 30251 2465
rect 30558 2456 30564 2468
rect 30616 2456 30622 2508
rect 32306 2456 32312 2508
rect 32364 2496 32370 2508
rect 32401 2499 32459 2505
rect 32401 2496 32413 2499
rect 32364 2468 32413 2496
rect 32364 2456 32370 2468
rect 32401 2465 32413 2468
rect 32447 2465 32459 2499
rect 32401 2459 32459 2465
rect 33686 2456 33692 2508
rect 33744 2496 33750 2508
rect 37292 2505 37320 2536
rect 34977 2499 35035 2505
rect 34977 2496 34989 2499
rect 33744 2468 34989 2496
rect 33744 2456 33750 2468
rect 34977 2465 34989 2468
rect 35023 2465 35035 2499
rect 35989 2499 36047 2505
rect 35989 2496 36001 2499
rect 34977 2459 35035 2465
rect 35866 2468 36001 2496
rect 1949 2431 2007 2437
rect 1949 2397 1961 2431
rect 1995 2428 2007 2431
rect 2314 2428 2320 2440
rect 1995 2400 2320 2428
rect 1995 2397 2007 2400
rect 1949 2391 2007 2397
rect 2314 2388 2320 2400
rect 2372 2428 2378 2440
rect 2409 2431 2467 2437
rect 2409 2428 2421 2431
rect 2372 2400 2421 2428
rect 2372 2388 2378 2400
rect 2409 2397 2421 2400
rect 2455 2397 2467 2431
rect 3050 2428 3056 2440
rect 3011 2400 3056 2428
rect 2409 2391 2467 2397
rect 3050 2388 3056 2400
rect 3108 2388 3114 2440
rect 4157 2431 4215 2437
rect 4157 2397 4169 2431
rect 4203 2428 4215 2431
rect 4890 2428 4896 2440
rect 4203 2400 4896 2428
rect 4203 2397 4215 2400
rect 4157 2391 4215 2397
rect 4890 2388 4896 2400
rect 4948 2388 4954 2440
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2428 5043 2431
rect 5258 2428 5264 2440
rect 5031 2400 5264 2428
rect 5031 2397 5043 2400
rect 4985 2391 5043 2397
rect 5258 2388 5264 2400
rect 5316 2388 5322 2440
rect 5629 2431 5687 2437
rect 5629 2397 5641 2431
rect 5675 2428 5687 2431
rect 5994 2428 6000 2440
rect 5675 2400 6000 2428
rect 5675 2397 5687 2400
rect 5629 2391 5687 2397
rect 5994 2388 6000 2400
rect 6052 2388 6058 2440
rect 6730 2388 6736 2440
rect 6788 2428 6794 2440
rect 6825 2431 6883 2437
rect 6825 2428 6837 2431
rect 6788 2400 6837 2428
rect 6788 2388 6794 2400
rect 6825 2397 6837 2400
rect 6871 2397 6883 2431
rect 6825 2391 6883 2397
rect 7466 2388 7472 2440
rect 7524 2428 7530 2440
rect 7561 2431 7619 2437
rect 7561 2428 7573 2431
rect 7524 2400 7573 2428
rect 7524 2388 7530 2400
rect 7561 2397 7573 2400
rect 7607 2397 7619 2431
rect 7561 2391 7619 2397
rect 8294 2388 8300 2440
rect 8352 2428 8358 2440
rect 8389 2431 8447 2437
rect 8389 2428 8401 2431
rect 8352 2400 8401 2428
rect 8352 2388 8358 2400
rect 8389 2397 8401 2400
rect 8435 2428 8447 2431
rect 8941 2431 8999 2437
rect 8941 2428 8953 2431
rect 8435 2400 8953 2428
rect 8435 2397 8447 2400
rect 8389 2391 8447 2397
rect 8941 2397 8953 2400
rect 8987 2397 8999 2431
rect 9674 2428 9680 2440
rect 9635 2400 9680 2428
rect 8941 2391 8999 2397
rect 9674 2388 9680 2400
rect 9732 2388 9738 2440
rect 10137 2431 10195 2437
rect 10137 2397 10149 2431
rect 10183 2428 10195 2431
rect 10410 2428 10416 2440
rect 10183 2400 10416 2428
rect 10183 2397 10195 2400
rect 10137 2391 10195 2397
rect 10410 2388 10416 2400
rect 10468 2388 10474 2440
rect 10781 2431 10839 2437
rect 10781 2397 10793 2431
rect 10827 2428 10839 2431
rect 10962 2428 10968 2440
rect 10827 2400 10968 2428
rect 10827 2397 10839 2400
rect 10781 2391 10839 2397
rect 10962 2388 10968 2400
rect 11020 2388 11026 2440
rect 11882 2388 11888 2440
rect 11940 2428 11946 2440
rect 11977 2431 12035 2437
rect 11977 2428 11989 2431
rect 11940 2400 11989 2428
rect 11940 2388 11946 2400
rect 11977 2397 11989 2400
rect 12023 2397 12035 2431
rect 11977 2391 12035 2397
rect 12618 2388 12624 2440
rect 12676 2428 12682 2440
rect 12713 2431 12771 2437
rect 12713 2428 12725 2431
rect 12676 2400 12725 2428
rect 12676 2388 12682 2400
rect 12713 2397 12725 2400
rect 12759 2397 12771 2431
rect 13354 2428 13360 2440
rect 13315 2400 13360 2428
rect 12713 2391 12771 2397
rect 13354 2388 13360 2400
rect 13412 2428 13418 2440
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 13412 2400 14105 2428
rect 13412 2388 13418 2400
rect 14093 2397 14105 2400
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 14645 2431 14703 2437
rect 14645 2397 14657 2431
rect 14691 2428 14703 2431
rect 14826 2428 14832 2440
rect 14691 2400 14832 2428
rect 14691 2397 14703 2400
rect 14645 2391 14703 2397
rect 14826 2388 14832 2400
rect 14884 2388 14890 2440
rect 15289 2431 15347 2437
rect 15289 2397 15301 2431
rect 15335 2428 15347 2431
rect 15562 2428 15568 2440
rect 15335 2400 15568 2428
rect 15335 2397 15347 2400
rect 15289 2391 15347 2397
rect 15562 2388 15568 2400
rect 15620 2388 15626 2440
rect 15933 2431 15991 2437
rect 15933 2397 15945 2431
rect 15979 2428 15991 2431
rect 16298 2428 16304 2440
rect 15979 2400 16304 2428
rect 15979 2397 15991 2400
rect 15933 2391 15991 2397
rect 16298 2388 16304 2400
rect 16356 2388 16362 2440
rect 17034 2388 17040 2440
rect 17092 2428 17098 2440
rect 17129 2431 17187 2437
rect 17129 2428 17141 2431
rect 17092 2400 17141 2428
rect 17092 2388 17098 2400
rect 17129 2397 17141 2400
rect 17175 2397 17187 2431
rect 17129 2391 17187 2397
rect 17770 2388 17776 2440
rect 17828 2428 17834 2440
rect 17865 2431 17923 2437
rect 17865 2428 17877 2431
rect 17828 2400 17877 2428
rect 17828 2388 17834 2400
rect 17865 2397 17877 2400
rect 17911 2397 17923 2431
rect 17865 2391 17923 2397
rect 18506 2388 18512 2440
rect 18564 2428 18570 2440
rect 18693 2431 18751 2437
rect 18693 2428 18705 2431
rect 18564 2400 18705 2428
rect 18564 2388 18570 2400
rect 18693 2397 18705 2400
rect 18739 2397 18751 2431
rect 19334 2428 19340 2440
rect 19295 2400 19340 2428
rect 18693 2391 18751 2397
rect 19334 2388 19340 2400
rect 19392 2388 19398 2440
rect 19978 2388 19984 2440
rect 20036 2428 20042 2440
rect 20257 2431 20315 2437
rect 20257 2428 20269 2431
rect 20036 2400 20269 2428
rect 20036 2388 20042 2400
rect 20257 2397 20269 2400
rect 20303 2397 20315 2431
rect 20257 2391 20315 2397
rect 20714 2388 20720 2440
rect 20772 2428 20778 2440
rect 20993 2431 21051 2437
rect 20993 2428 21005 2431
rect 20772 2400 21005 2428
rect 20772 2388 20778 2400
rect 20993 2397 21005 2400
rect 21039 2397 21051 2431
rect 20993 2391 21051 2397
rect 22557 2431 22615 2437
rect 22557 2397 22569 2431
rect 22603 2428 22615 2431
rect 22922 2428 22928 2440
rect 22603 2400 22928 2428
rect 22603 2397 22615 2400
rect 22557 2391 22615 2397
rect 22922 2388 22928 2400
rect 22980 2388 22986 2440
rect 23014 2388 23020 2440
rect 23072 2428 23078 2440
rect 23661 2431 23719 2437
rect 23661 2428 23673 2431
rect 23072 2400 23673 2428
rect 23072 2388 23078 2400
rect 23661 2397 23673 2400
rect 23707 2397 23719 2431
rect 23661 2391 23719 2397
rect 23750 2388 23756 2440
rect 23808 2428 23814 2440
rect 24210 2428 24216 2440
rect 23808 2400 24216 2428
rect 23808 2388 23814 2400
rect 24210 2388 24216 2400
rect 24268 2428 24274 2440
rect 24397 2431 24455 2437
rect 24397 2428 24409 2431
rect 24268 2400 24409 2428
rect 24268 2388 24274 2400
rect 24397 2397 24409 2400
rect 24443 2397 24455 2431
rect 25038 2428 25044 2440
rect 24999 2400 25044 2428
rect 24397 2391 24455 2397
rect 25038 2388 25044 2400
rect 25096 2388 25102 2440
rect 25130 2388 25136 2440
rect 25188 2428 25194 2440
rect 25685 2431 25743 2437
rect 25685 2428 25697 2431
rect 25188 2400 25697 2428
rect 25188 2388 25194 2400
rect 25685 2397 25697 2400
rect 25731 2428 25743 2431
rect 26329 2431 26387 2437
rect 26329 2428 26341 2431
rect 25731 2400 26341 2428
rect 25731 2397 25743 2400
rect 25685 2391 25743 2397
rect 26329 2397 26341 2400
rect 26375 2397 26387 2431
rect 26329 2391 26387 2397
rect 26602 2388 26608 2440
rect 26660 2428 26666 2440
rect 26970 2428 26976 2440
rect 26660 2400 26976 2428
rect 26660 2388 26666 2400
rect 26970 2388 26976 2400
rect 27028 2388 27034 2440
rect 27614 2428 27620 2440
rect 27575 2400 27620 2428
rect 27614 2388 27620 2400
rect 27672 2388 27678 2440
rect 28074 2388 28080 2440
rect 28132 2428 28138 2440
rect 28261 2431 28319 2437
rect 28261 2428 28273 2431
rect 28132 2400 28273 2428
rect 28132 2388 28138 2400
rect 28261 2397 28273 2400
rect 28307 2428 28319 2431
rect 28905 2431 28963 2437
rect 28905 2428 28917 2431
rect 28307 2400 28917 2428
rect 28307 2397 28319 2400
rect 28261 2391 28319 2397
rect 28905 2397 28917 2400
rect 28951 2397 28963 2431
rect 28905 2391 28963 2397
rect 29546 2388 29552 2440
rect 29604 2428 29610 2440
rect 30469 2431 30527 2437
rect 30469 2428 30481 2431
rect 29604 2400 30481 2428
rect 29604 2388 29610 2400
rect 30469 2397 30481 2400
rect 30515 2428 30527 2431
rect 30929 2431 30987 2437
rect 30929 2428 30941 2431
rect 30515 2400 30941 2428
rect 30515 2397 30527 2400
rect 30469 2391 30527 2397
rect 30929 2397 30941 2400
rect 30975 2397 30987 2431
rect 32125 2431 32183 2437
rect 32125 2428 32137 2431
rect 30929 2391 30987 2397
rect 31496 2400 32137 2428
rect 10502 2360 10508 2372
rect 2608 2332 10508 2360
rect 2608 2301 2636 2332
rect 10502 2320 10508 2332
rect 10560 2320 10566 2372
rect 13446 2360 13452 2372
rect 10612 2332 13452 2360
rect 2593 2295 2651 2301
rect 2593 2261 2605 2295
rect 2639 2261 2651 2295
rect 2593 2255 2651 2261
rect 3786 2252 3792 2304
rect 3844 2292 3850 2304
rect 3973 2295 4031 2301
rect 3973 2292 3985 2295
rect 3844 2264 3985 2292
rect 3844 2252 3850 2264
rect 3973 2261 3985 2264
rect 4019 2261 4031 2295
rect 3973 2255 4031 2261
rect 6914 2252 6920 2304
rect 6972 2292 6978 2304
rect 10612 2292 10640 2332
rect 13446 2320 13452 2332
rect 13504 2320 13510 2372
rect 6972 2264 10640 2292
rect 10965 2295 11023 2301
rect 6972 2252 6978 2264
rect 10965 2261 10977 2295
rect 11011 2292 11023 2295
rect 13262 2292 13268 2304
rect 11011 2264 13268 2292
rect 11011 2261 11023 2264
rect 10965 2255 11023 2261
rect 13262 2252 13268 2264
rect 13320 2252 13326 2304
rect 22186 2252 22192 2304
rect 22244 2292 22250 2304
rect 22373 2295 22431 2301
rect 22373 2292 22385 2295
rect 22244 2264 22385 2292
rect 22244 2252 22250 2264
rect 22373 2261 22385 2264
rect 22419 2261 22431 2295
rect 22373 2255 22431 2261
rect 31018 2252 31024 2304
rect 31076 2292 31082 2304
rect 31496 2301 31524 2400
rect 32125 2397 32137 2400
rect 32171 2397 32183 2431
rect 32125 2391 32183 2397
rect 34606 2388 34612 2440
rect 34664 2428 34670 2440
rect 34701 2431 34759 2437
rect 34701 2428 34713 2431
rect 34664 2400 34713 2428
rect 34664 2388 34670 2400
rect 34701 2397 34713 2400
rect 34747 2428 34759 2431
rect 35866 2428 35894 2468
rect 35989 2465 36001 2468
rect 36035 2465 36047 2499
rect 35989 2459 36047 2465
rect 37277 2499 37335 2505
rect 37277 2465 37289 2499
rect 37323 2465 37335 2499
rect 37277 2459 37335 2465
rect 36722 2428 36728 2440
rect 34747 2400 35894 2428
rect 36683 2400 36728 2428
rect 34747 2397 34759 2400
rect 34701 2391 34759 2397
rect 36722 2388 36728 2400
rect 36780 2388 36786 2440
rect 37553 2431 37611 2437
rect 37553 2397 37565 2431
rect 37599 2397 37611 2431
rect 37553 2391 37611 2397
rect 35526 2320 35532 2372
rect 35584 2360 35590 2372
rect 37568 2360 37596 2391
rect 35584 2332 37596 2360
rect 35584 2320 35590 2332
rect 31481 2295 31539 2301
rect 31481 2292 31493 2295
rect 31076 2264 31493 2292
rect 31076 2252 31082 2264
rect 31481 2261 31493 2264
rect 31527 2261 31539 2295
rect 31481 2255 31539 2261
rect 33962 2252 33968 2304
rect 34020 2292 34026 2304
rect 34057 2295 34115 2301
rect 34057 2292 34069 2295
rect 34020 2264 34069 2292
rect 34020 2252 34026 2264
rect 34057 2261 34069 2264
rect 34103 2261 34115 2295
rect 34057 2255 34115 2261
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 36176 37408 36228 37460
rect 2320 37272 2372 37324
rect 5264 37272 5316 37324
rect 7472 37272 7524 37324
rect 10416 37340 10468 37392
rect 11888 37272 11940 37324
rect 2688 37247 2740 37256
rect 2688 37213 2697 37247
rect 2697 37213 2731 37247
rect 2731 37213 2740 37247
rect 2688 37204 2740 37213
rect 4988 37204 5040 37256
rect 6552 37204 6604 37256
rect 8024 37204 8076 37256
rect 10416 37247 10468 37256
rect 10416 37213 10425 37247
rect 10425 37213 10459 37247
rect 10459 37213 10468 37247
rect 10416 37204 10468 37213
rect 12164 37204 12216 37256
rect 13360 37247 13412 37256
rect 13360 37213 13369 37247
rect 13369 37213 13403 37247
rect 13403 37213 13412 37247
rect 13360 37204 13412 37213
rect 14832 37204 14884 37256
rect 15568 37204 15620 37256
rect 16304 37204 16356 37256
rect 17040 37204 17092 37256
rect 17776 37204 17828 37256
rect 18512 37204 18564 37256
rect 19248 37204 19300 37256
rect 19984 37204 20036 37256
rect 20720 37204 20772 37256
rect 22284 37247 22336 37256
rect 22284 37213 22293 37247
rect 22293 37213 22327 37247
rect 22327 37213 22336 37247
rect 22284 37204 22336 37213
rect 22928 37204 22980 37256
rect 25136 37272 25188 37324
rect 24584 37247 24636 37256
rect 24584 37213 24593 37247
rect 24593 37213 24627 37247
rect 24627 37213 24636 37247
rect 24584 37204 24636 37213
rect 24860 37204 24912 37256
rect 34704 37272 34756 37324
rect 26608 37204 26660 37256
rect 26976 37247 27028 37256
rect 26976 37213 26985 37247
rect 26985 37213 27019 37247
rect 27019 37213 27028 37247
rect 26976 37204 27028 37213
rect 27344 37204 27396 37256
rect 27620 37204 27672 37256
rect 28080 37204 28132 37256
rect 29368 37204 29420 37256
rect 30012 37204 30064 37256
rect 30472 37204 30524 37256
rect 31760 37204 31812 37256
rect 32220 37204 32272 37256
rect 32496 37204 32548 37256
rect 33232 37204 33284 37256
rect 34520 37204 34572 37256
rect 35900 37204 35952 37256
rect 36452 37204 36504 37256
rect 3792 37068 3844 37120
rect 13544 37111 13596 37120
rect 13544 37077 13553 37111
rect 13553 37077 13587 37111
rect 13587 37077 13596 37111
rect 13544 37068 13596 37077
rect 15016 37068 15068 37120
rect 15752 37068 15804 37120
rect 16396 37068 16448 37120
rect 17868 37068 17920 37120
rect 18052 37111 18104 37120
rect 18052 37077 18061 37111
rect 18061 37077 18095 37111
rect 18095 37077 18104 37111
rect 18052 37068 18104 37077
rect 18236 37068 18288 37120
rect 19432 37068 19484 37120
rect 20536 37068 20588 37120
rect 20812 37068 20864 37120
rect 22192 37068 22244 37120
rect 22836 37068 22888 37120
rect 23756 37068 23808 37120
rect 24768 37068 24820 37120
rect 25320 37068 25372 37120
rect 27344 37068 27396 37120
rect 27528 37068 27580 37120
rect 28264 37111 28316 37120
rect 28264 37077 28273 37111
rect 28273 37077 28307 37111
rect 28307 37077 28316 37111
rect 28264 37068 28316 37077
rect 28724 37068 28776 37120
rect 29644 37068 29696 37120
rect 30380 37068 30432 37120
rect 32128 37111 32180 37120
rect 32128 37077 32137 37111
rect 32137 37077 32171 37111
rect 32171 37077 32180 37111
rect 32128 37068 32180 37077
rect 32588 37068 32640 37120
rect 33416 37111 33468 37120
rect 33416 37077 33425 37111
rect 33425 37077 33459 37111
rect 33459 37077 33468 37111
rect 33416 37068 33468 37077
rect 33784 37068 33836 37120
rect 34796 37068 34848 37120
rect 35532 37068 35584 37120
rect 38016 37111 38068 37120
rect 38016 37077 38025 37111
rect 38025 37077 38059 37111
rect 38059 37077 38068 37111
rect 38016 37068 38068 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 14832 36864 14884 36916
rect 15568 36907 15620 36916
rect 15568 36873 15577 36907
rect 15577 36873 15611 36907
rect 15611 36873 15620 36907
rect 15568 36864 15620 36873
rect 16304 36864 16356 36916
rect 17040 36907 17092 36916
rect 17040 36873 17049 36907
rect 17049 36873 17083 36907
rect 17083 36873 17092 36907
rect 17040 36864 17092 36873
rect 17776 36907 17828 36916
rect 17776 36873 17785 36907
rect 17785 36873 17819 36907
rect 17819 36873 17828 36907
rect 17776 36864 17828 36873
rect 18512 36864 18564 36916
rect 19248 36907 19300 36916
rect 19248 36873 19257 36907
rect 19257 36873 19291 36907
rect 19291 36873 19300 36907
rect 19248 36864 19300 36873
rect 19984 36907 20036 36916
rect 19984 36873 19993 36907
rect 19993 36873 20027 36907
rect 20027 36873 20036 36907
rect 19984 36864 20036 36873
rect 20720 36907 20772 36916
rect 20720 36873 20729 36907
rect 20729 36873 20763 36907
rect 20763 36873 20772 36907
rect 20720 36864 20772 36873
rect 23664 36864 23716 36916
rect 24584 36864 24636 36916
rect 24860 36907 24912 36916
rect 24860 36873 24869 36907
rect 24869 36873 24903 36907
rect 24903 36873 24912 36907
rect 24860 36864 24912 36873
rect 25872 36864 25924 36916
rect 26976 36907 27028 36916
rect 26976 36873 26985 36907
rect 26985 36873 27019 36907
rect 27019 36873 27028 36907
rect 26976 36864 27028 36873
rect 27620 36907 27672 36916
rect 27620 36873 27629 36907
rect 27629 36873 27663 36907
rect 27663 36873 27672 36907
rect 27620 36864 27672 36873
rect 29552 36864 29604 36916
rect 30012 36907 30064 36916
rect 30012 36873 30021 36907
rect 30021 36873 30055 36907
rect 30055 36873 30064 36907
rect 30012 36864 30064 36873
rect 31024 36864 31076 36916
rect 32220 36907 32272 36916
rect 32220 36873 32229 36907
rect 32229 36873 32263 36907
rect 32263 36873 32272 36907
rect 32220 36864 32272 36873
rect 32496 36864 32548 36916
rect 34520 36907 34572 36916
rect 34520 36873 34529 36907
rect 34529 36873 34563 36907
rect 34563 36873 34572 36907
rect 34520 36864 34572 36873
rect 36268 36907 36320 36916
rect 36268 36873 36277 36907
rect 36277 36873 36311 36907
rect 36311 36873 36320 36907
rect 36268 36864 36320 36873
rect 36912 36864 36964 36916
rect 3056 36728 3108 36780
rect 4620 36771 4672 36780
rect 4620 36737 4629 36771
rect 4629 36737 4663 36771
rect 4663 36737 4672 36771
rect 4620 36728 4672 36737
rect 6736 36728 6788 36780
rect 8208 36728 8260 36780
rect 9680 36728 9732 36780
rect 11152 36728 11204 36780
rect 12624 36728 12676 36780
rect 14096 36728 14148 36780
rect 21456 36728 21508 36780
rect 3424 36703 3476 36712
rect 3424 36669 3433 36703
rect 3433 36669 3467 36703
rect 3467 36669 3476 36703
rect 3424 36660 3476 36669
rect 4896 36703 4948 36712
rect 4896 36669 4905 36703
rect 4905 36669 4939 36703
rect 4939 36669 4948 36703
rect 4896 36660 4948 36669
rect 7104 36703 7156 36712
rect 7104 36669 7113 36703
rect 7113 36669 7147 36703
rect 7147 36669 7156 36703
rect 7104 36660 7156 36669
rect 8852 36660 8904 36712
rect 10048 36703 10100 36712
rect 10048 36669 10057 36703
rect 10057 36669 10091 36703
rect 10091 36669 10100 36703
rect 10048 36660 10100 36669
rect 11980 36660 12032 36712
rect 36176 36728 36228 36780
rect 36544 36728 36596 36780
rect 35348 36660 35400 36712
rect 37648 36660 37700 36712
rect 36360 36592 36412 36644
rect 37188 36592 37240 36644
rect 12992 36567 13044 36576
rect 12992 36533 13001 36567
rect 13001 36533 13035 36567
rect 13035 36533 13044 36567
rect 12992 36524 13044 36533
rect 14832 36524 14884 36576
rect 22192 36524 22244 36576
rect 25780 36524 25832 36576
rect 29368 36567 29420 36576
rect 29368 36533 29377 36567
rect 29377 36533 29411 36567
rect 29411 36533 29420 36567
rect 29368 36524 29420 36533
rect 31116 36567 31168 36576
rect 31116 36533 31125 36567
rect 31125 36533 31159 36567
rect 31159 36533 31168 36567
rect 31116 36524 31168 36533
rect 37464 36524 37516 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 4620 36320 4672 36372
rect 4712 36320 4764 36372
rect 4988 36363 5040 36372
rect 4988 36329 4997 36363
rect 4997 36329 5031 36363
rect 5031 36329 5040 36363
rect 4988 36320 5040 36329
rect 6736 36320 6788 36372
rect 8208 36363 8260 36372
rect 8208 36329 8217 36363
rect 8217 36329 8251 36363
rect 8251 36329 8260 36363
rect 8208 36320 8260 36329
rect 9680 36320 9732 36372
rect 11152 36320 11204 36372
rect 11888 36363 11940 36372
rect 11888 36329 11897 36363
rect 11897 36329 11931 36363
rect 11931 36329 11940 36363
rect 11888 36320 11940 36329
rect 12624 36363 12676 36372
rect 12624 36329 12633 36363
rect 12633 36329 12667 36363
rect 12667 36329 12676 36363
rect 12624 36320 12676 36329
rect 35348 36363 35400 36372
rect 35348 36329 35357 36363
rect 35357 36329 35391 36363
rect 35391 36329 35400 36363
rect 35348 36320 35400 36329
rect 6000 36184 6052 36236
rect 8944 36184 8996 36236
rect 38108 36227 38160 36236
rect 38108 36193 38117 36227
rect 38117 36193 38151 36227
rect 38151 36193 38160 36227
rect 38108 36184 38160 36193
rect 6368 36159 6420 36168
rect 6368 36125 6377 36159
rect 6377 36125 6411 36159
rect 6411 36125 6420 36159
rect 6368 36116 6420 36125
rect 9220 36116 9272 36168
rect 36176 36116 36228 36168
rect 37832 36159 37884 36168
rect 37832 36125 37841 36159
rect 37841 36125 37875 36159
rect 37875 36125 37884 36159
rect 37832 36116 37884 36125
rect 36452 36091 36504 36100
rect 36452 36057 36461 36091
rect 36461 36057 36495 36091
rect 36495 36057 36504 36091
rect 36452 36048 36504 36057
rect 35992 36023 36044 36032
rect 35992 35989 36001 36023
rect 36001 35989 36035 36023
rect 36035 35989 36044 36023
rect 35992 35980 36044 35989
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 8944 35819 8996 35828
rect 8944 35785 8953 35819
rect 8953 35785 8987 35819
rect 8987 35785 8996 35819
rect 8944 35776 8996 35785
rect 28816 35776 28868 35828
rect 29368 35776 29420 35828
rect 35808 35776 35860 35828
rect 36176 35819 36228 35828
rect 36176 35785 36185 35819
rect 36185 35785 36219 35819
rect 36219 35785 36228 35819
rect 36176 35776 36228 35785
rect 36728 35640 36780 35692
rect 37648 35572 37700 35624
rect 37096 35504 37148 35556
rect 35900 35436 35952 35488
rect 36452 35436 36504 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 36820 35071 36872 35080
rect 36820 35037 36829 35071
rect 36829 35037 36863 35071
rect 36863 35037 36872 35071
rect 36820 35028 36872 35037
rect 37740 35071 37792 35080
rect 37740 35037 37749 35071
rect 37749 35037 37783 35071
rect 37783 35037 37792 35071
rect 37740 35028 37792 35037
rect 37924 35071 37976 35080
rect 37924 35037 37933 35071
rect 37933 35037 37967 35071
rect 37967 35037 37976 35071
rect 37924 35028 37976 35037
rect 35440 34892 35492 34944
rect 38016 34960 38068 35012
rect 35900 34892 35952 34944
rect 37004 34935 37056 34944
rect 37004 34901 37013 34935
rect 37013 34901 37047 34935
rect 37047 34901 37056 34935
rect 37004 34892 37056 34901
rect 37556 34935 37608 34944
rect 37556 34901 37565 34935
rect 37565 34901 37599 34935
rect 37599 34901 37608 34935
rect 37556 34892 37608 34901
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 35440 34731 35492 34740
rect 35440 34697 35449 34731
rect 35449 34697 35483 34731
rect 35483 34697 35492 34731
rect 35440 34688 35492 34697
rect 36544 34688 36596 34740
rect 37832 34688 37884 34740
rect 37556 34620 37608 34672
rect 35992 34552 36044 34604
rect 37648 34552 37700 34604
rect 38016 34620 38068 34672
rect 37924 34595 37976 34604
rect 37924 34561 37933 34595
rect 37933 34561 37967 34595
rect 37967 34561 37976 34595
rect 37924 34552 37976 34561
rect 38200 34552 38252 34604
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 37740 34144 37792 34196
rect 35900 34008 35952 34060
rect 38016 34008 38068 34060
rect 36268 33983 36320 33992
rect 36268 33949 36277 33983
rect 36277 33949 36311 33983
rect 36311 33949 36320 33983
rect 36268 33940 36320 33949
rect 37464 33983 37516 33992
rect 37464 33949 37473 33983
rect 37473 33949 37507 33983
rect 37507 33949 37516 33983
rect 37464 33940 37516 33949
rect 36452 33804 36504 33856
rect 36544 33804 36596 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 36728 33643 36780 33652
rect 36728 33609 36737 33643
rect 36737 33609 36771 33643
rect 36771 33609 36780 33643
rect 36728 33600 36780 33609
rect 37464 33600 37516 33652
rect 38200 33600 38252 33652
rect 36544 33507 36596 33516
rect 36544 33473 36553 33507
rect 36553 33473 36587 33507
rect 36587 33473 36596 33507
rect 36544 33464 36596 33473
rect 38016 33464 38068 33516
rect 37648 33439 37700 33448
rect 37648 33405 37657 33439
rect 37657 33405 37691 33439
rect 37691 33405 37700 33439
rect 37648 33396 37700 33405
rect 34520 33260 34572 33312
rect 35992 33303 36044 33312
rect 35992 33269 36001 33303
rect 36001 33269 36035 33303
rect 36035 33269 36044 33303
rect 35992 33260 36044 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 37280 33099 37332 33108
rect 37280 33065 37289 33099
rect 37289 33065 37323 33099
rect 37323 33065 37332 33099
rect 37280 33056 37332 33065
rect 34520 32920 34572 32972
rect 35532 32895 35584 32904
rect 35532 32861 35541 32895
rect 35541 32861 35575 32895
rect 35575 32861 35584 32895
rect 35532 32852 35584 32861
rect 37832 32895 37884 32904
rect 37832 32861 37841 32895
rect 37841 32861 37875 32895
rect 37875 32861 37884 32895
rect 37832 32852 37884 32861
rect 35440 32827 35492 32836
rect 35440 32793 35449 32827
rect 35449 32793 35483 32827
rect 35483 32793 35492 32827
rect 35440 32784 35492 32793
rect 35992 32784 36044 32836
rect 38016 32759 38068 32768
rect 38016 32725 38025 32759
rect 38025 32725 38059 32759
rect 38059 32725 38068 32759
rect 38016 32716 38068 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 34796 32555 34848 32564
rect 34796 32521 34805 32555
rect 34805 32521 34839 32555
rect 34839 32521 34848 32555
rect 34796 32512 34848 32521
rect 37832 32512 37884 32564
rect 37832 32419 37884 32428
rect 37832 32385 37841 32419
rect 37841 32385 37875 32419
rect 37875 32385 37884 32419
rect 37832 32376 37884 32385
rect 34520 32351 34572 32360
rect 31668 32172 31720 32224
rect 34520 32317 34529 32351
rect 34529 32317 34563 32351
rect 34563 32317 34572 32351
rect 34520 32308 34572 32317
rect 34704 32351 34756 32360
rect 34704 32317 34713 32351
rect 34713 32317 34747 32351
rect 34747 32317 34756 32351
rect 34704 32308 34756 32317
rect 37648 32240 37700 32292
rect 38016 32215 38068 32224
rect 38016 32181 38025 32215
rect 38025 32181 38059 32215
rect 38059 32181 38068 32215
rect 38016 32172 38068 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 34704 31968 34756 32020
rect 37740 31968 37792 32020
rect 38108 32011 38160 32020
rect 38108 31977 38117 32011
rect 38117 31977 38151 32011
rect 38151 31977 38160 32011
rect 38108 31968 38160 31977
rect 33600 31875 33652 31884
rect 33600 31841 33609 31875
rect 33609 31841 33643 31875
rect 33643 31841 33652 31875
rect 33600 31832 33652 31841
rect 37832 31900 37884 31952
rect 33784 31739 33836 31748
rect 33784 31705 33793 31739
rect 33793 31705 33827 31739
rect 33827 31705 33836 31739
rect 33784 31696 33836 31705
rect 33968 31628 34020 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 34612 31288 34664 31340
rect 33600 31152 33652 31204
rect 35900 31152 35952 31204
rect 38016 31195 38068 31204
rect 38016 31161 38025 31195
rect 38025 31161 38059 31195
rect 38059 31161 38068 31195
rect 38016 31152 38068 31161
rect 33968 31084 34020 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 34520 30676 34572 30728
rect 32496 30540 32548 30592
rect 38016 30583 38068 30592
rect 38016 30549 38025 30583
rect 38025 30549 38059 30583
rect 38059 30549 38068 30583
rect 38016 30540 38068 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 32588 30311 32640 30320
rect 32588 30277 32597 30311
rect 32597 30277 32631 30311
rect 32631 30277 32640 30311
rect 32588 30268 32640 30277
rect 32312 30175 32364 30184
rect 32312 30141 32321 30175
rect 32321 30141 32355 30175
rect 32355 30141 32364 30175
rect 32312 30132 32364 30141
rect 32496 30175 32548 30184
rect 32496 30141 32505 30175
rect 32505 30141 32539 30175
rect 32539 30141 32548 30175
rect 32496 30132 32548 30141
rect 33508 30200 33560 30252
rect 34152 30200 34204 30252
rect 34520 30064 34572 30116
rect 34612 29996 34664 30048
rect 38016 30039 38068 30048
rect 38016 30005 38025 30039
rect 38025 30005 38059 30039
rect 38059 30005 38068 30039
rect 38016 29996 38068 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 33508 29835 33560 29844
rect 33508 29801 33517 29835
rect 33517 29801 33551 29835
rect 33551 29801 33560 29835
rect 33508 29792 33560 29801
rect 30196 29656 30248 29708
rect 32312 29656 32364 29708
rect 32128 29588 32180 29640
rect 33416 29588 33468 29640
rect 33508 29588 33560 29640
rect 32404 29520 32456 29572
rect 32772 29452 32824 29504
rect 33600 29452 33652 29504
rect 38016 29495 38068 29504
rect 38016 29461 38025 29495
rect 38025 29461 38059 29495
rect 38059 29461 38068 29495
rect 38016 29452 38068 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 31116 29291 31168 29300
rect 31116 29257 31125 29291
rect 31125 29257 31159 29291
rect 31159 29257 31168 29291
rect 31116 29248 31168 29257
rect 33508 29248 33560 29300
rect 32772 29155 32824 29164
rect 32772 29121 32781 29155
rect 32781 29121 32815 29155
rect 32815 29121 32824 29155
rect 32772 29112 32824 29121
rect 30196 29044 30248 29096
rect 32312 29044 32364 29096
rect 34152 29044 34204 29096
rect 33600 29019 33652 29028
rect 33600 28985 33609 29019
rect 33609 28985 33643 29019
rect 33643 28985 33652 29019
rect 33600 28976 33652 28985
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 30196 28611 30248 28620
rect 30196 28577 30205 28611
rect 30205 28577 30239 28611
rect 30239 28577 30248 28611
rect 30196 28568 30248 28577
rect 30656 28568 30708 28620
rect 30380 28543 30432 28552
rect 30380 28509 30389 28543
rect 30389 28509 30423 28543
rect 30423 28509 30432 28543
rect 30380 28500 30432 28509
rect 32312 28364 32364 28416
rect 38016 28407 38068 28416
rect 38016 28373 38025 28407
rect 38025 28373 38059 28407
rect 38059 28373 38068 28407
rect 38016 28364 38068 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 29644 28203 29696 28212
rect 23848 28092 23900 28144
rect 29644 28169 29653 28203
rect 29653 28169 29687 28203
rect 29687 28169 29696 28203
rect 29644 28160 29696 28169
rect 31668 28092 31720 28144
rect 28172 28067 28224 28076
rect 28172 28033 28181 28067
rect 28181 28033 28215 28067
rect 28215 28033 28224 28067
rect 28172 28024 28224 28033
rect 28816 28024 28868 28076
rect 33692 28160 33744 28212
rect 37832 28067 37884 28076
rect 37832 28033 37841 28067
rect 37841 28033 37875 28067
rect 37875 28033 37884 28067
rect 37832 28024 37884 28033
rect 29184 27956 29236 28008
rect 30472 27956 30524 28008
rect 30196 27888 30248 27940
rect 29920 27820 29972 27872
rect 38016 27863 38068 27872
rect 38016 27829 38025 27863
rect 38025 27829 38059 27863
rect 38059 27829 38068 27863
rect 38016 27820 38068 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 28816 27616 28868 27668
rect 37832 27548 37884 27600
rect 30472 27480 30524 27532
rect 29920 27455 29972 27464
rect 29920 27421 29929 27455
rect 29929 27421 29963 27455
rect 29963 27421 29972 27455
rect 29920 27412 29972 27421
rect 37832 27455 37884 27464
rect 37832 27421 37841 27455
rect 37841 27421 37875 27455
rect 37875 27421 37884 27455
rect 37832 27412 37884 27421
rect 38016 27319 38068 27328
rect 38016 27285 38025 27319
rect 38025 27285 38059 27319
rect 38059 27285 38068 27319
rect 38016 27276 38068 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 28724 27072 28776 27124
rect 27988 26868 28040 26920
rect 29184 26936 29236 26988
rect 37832 27072 37884 27124
rect 37832 26979 37884 26988
rect 37832 26945 37841 26979
rect 37841 26945 37875 26979
rect 37875 26945 37884 26979
rect 37832 26936 37884 26945
rect 29092 26868 29144 26920
rect 38016 26775 38068 26784
rect 38016 26741 38025 26775
rect 38025 26741 38059 26775
rect 38059 26741 38068 26775
rect 38016 26732 38068 26741
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 27988 26435 28040 26444
rect 27988 26401 27997 26435
rect 27997 26401 28031 26435
rect 28031 26401 28040 26435
rect 27988 26392 28040 26401
rect 28264 26324 28316 26376
rect 28448 26256 28500 26308
rect 28540 26231 28592 26240
rect 28540 26197 28549 26231
rect 28549 26197 28583 26231
rect 28583 26197 28592 26231
rect 28540 26188 28592 26197
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 27344 26027 27396 26036
rect 27344 25993 27353 26027
rect 27353 25993 27387 26027
rect 27387 25993 27396 26027
rect 27344 25984 27396 25993
rect 37832 25984 37884 26036
rect 27160 25916 27212 25968
rect 27896 25848 27948 25900
rect 28540 25848 28592 25900
rect 27988 25712 28040 25764
rect 38016 25755 38068 25764
rect 38016 25721 38025 25755
rect 38025 25721 38059 25755
rect 38059 25721 38068 25755
rect 38016 25712 38068 25721
rect 27712 25687 27764 25696
rect 27712 25653 27721 25687
rect 27721 25653 27755 25687
rect 27755 25653 27764 25687
rect 27712 25644 27764 25653
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 27896 25483 27948 25492
rect 27896 25449 27905 25483
rect 27905 25449 27939 25483
rect 27939 25449 27948 25483
rect 27896 25440 27948 25449
rect 27988 25304 28040 25356
rect 27528 25279 27580 25288
rect 27528 25245 27537 25279
rect 27537 25245 27571 25279
rect 27571 25245 27580 25279
rect 27528 25236 27580 25245
rect 27712 25236 27764 25288
rect 27804 25100 27856 25152
rect 38016 25143 38068 25152
rect 38016 25109 38025 25143
rect 38025 25109 38059 25143
rect 38059 25109 38068 25143
rect 38016 25100 38068 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 26792 24760 26844 24812
rect 26056 24556 26108 24608
rect 27804 24556 27856 24608
rect 38016 24599 38068 24608
rect 38016 24565 38025 24599
rect 38025 24565 38059 24599
rect 38059 24565 38068 24599
rect 38016 24556 38068 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 26792 24395 26844 24404
rect 26792 24361 26801 24395
rect 26801 24361 26835 24395
rect 26835 24361 26844 24395
rect 26792 24352 26844 24361
rect 24492 24216 24544 24268
rect 25780 24191 25832 24200
rect 25780 24157 25789 24191
rect 25789 24157 25823 24191
rect 25823 24157 25832 24191
rect 25780 24148 25832 24157
rect 37832 24191 37884 24200
rect 37832 24157 37841 24191
rect 37841 24157 37875 24191
rect 37875 24157 37884 24191
rect 37832 24148 37884 24157
rect 26056 24012 26108 24064
rect 38016 24055 38068 24064
rect 38016 24021 38025 24055
rect 38025 24021 38059 24055
rect 38059 24021 38068 24055
rect 38016 24012 38068 24021
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 25320 23808 25372 23860
rect 24492 23604 24544 23656
rect 26240 23604 26292 23656
rect 23020 23536 23072 23588
rect 28172 23536 28224 23588
rect 37832 23468 37884 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 36820 23307 36872 23316
rect 36820 23273 36829 23307
rect 36829 23273 36863 23307
rect 36863 23273 36872 23307
rect 36820 23264 36872 23273
rect 23112 23128 23164 23180
rect 24492 23171 24544 23180
rect 24492 23137 24501 23171
rect 24501 23137 24535 23171
rect 24535 23137 24544 23171
rect 24492 23128 24544 23137
rect 25228 23128 25280 23180
rect 23020 23103 23072 23112
rect 23020 23069 23029 23103
rect 23029 23069 23063 23103
rect 23063 23069 23072 23103
rect 23020 23060 23072 23069
rect 24768 23103 24820 23112
rect 24768 23069 24777 23103
rect 24777 23069 24811 23103
rect 24811 23069 24820 23103
rect 24768 23060 24820 23069
rect 23112 22967 23164 22976
rect 23112 22933 23121 22967
rect 23121 22933 23155 22967
rect 23155 22933 23164 22967
rect 23112 22924 23164 22933
rect 36728 23060 36780 23112
rect 26240 22967 26292 22976
rect 26240 22933 26249 22967
rect 26249 22933 26283 22967
rect 26283 22933 26292 22967
rect 38016 22967 38068 22976
rect 26240 22924 26292 22933
rect 38016 22933 38025 22967
rect 38025 22933 38059 22967
rect 38059 22933 38068 22967
rect 38016 22924 38068 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 23756 22763 23808 22772
rect 23756 22729 23765 22763
rect 23765 22729 23799 22763
rect 23799 22729 23808 22763
rect 23756 22720 23808 22729
rect 36360 22763 36412 22772
rect 36360 22729 36369 22763
rect 36369 22729 36403 22763
rect 36403 22729 36412 22763
rect 36360 22720 36412 22729
rect 36728 22763 36780 22772
rect 36728 22729 36737 22763
rect 36737 22729 36771 22763
rect 36771 22729 36780 22763
rect 36728 22720 36780 22729
rect 22744 22516 22796 22568
rect 23112 22516 23164 22568
rect 24584 22448 24636 22500
rect 25228 22423 25280 22432
rect 25228 22389 25237 22423
rect 25237 22389 25271 22423
rect 25271 22389 25280 22423
rect 25228 22380 25280 22389
rect 25320 22380 25372 22432
rect 36636 22516 36688 22568
rect 38016 22423 38068 22432
rect 38016 22389 38025 22423
rect 38025 22389 38059 22423
rect 38059 22389 38068 22423
rect 38016 22380 38068 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 20260 22176 20312 22228
rect 25320 22176 25372 22228
rect 22376 21972 22428 22024
rect 37832 22015 37884 22024
rect 37832 21981 37841 22015
rect 37841 21981 37875 22015
rect 37875 21981 37884 22015
rect 37832 21972 37884 21981
rect 22284 21879 22336 21888
rect 22284 21845 22293 21879
rect 22293 21845 22327 21879
rect 22327 21845 22336 21879
rect 22284 21836 22336 21845
rect 23296 21836 23348 21888
rect 24584 21836 24636 21888
rect 38016 21879 38068 21888
rect 38016 21845 38025 21879
rect 38025 21845 38059 21879
rect 38059 21845 38068 21879
rect 38016 21836 38068 21845
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 22836 21632 22888 21684
rect 38108 21539 38160 21548
rect 38108 21505 38117 21539
rect 38117 21505 38151 21539
rect 38151 21505 38160 21539
rect 38108 21496 38160 21505
rect 22744 21471 22796 21480
rect 22744 21437 22753 21471
rect 22753 21437 22787 21471
rect 22787 21437 22796 21471
rect 22744 21428 22796 21437
rect 23296 21428 23348 21480
rect 24032 21335 24084 21344
rect 24032 21301 24041 21335
rect 24041 21301 24075 21335
rect 24075 21301 24084 21335
rect 24032 21292 24084 21301
rect 37924 21335 37976 21344
rect 37924 21301 37933 21335
rect 37933 21301 37967 21335
rect 37967 21301 37976 21335
rect 37924 21292 37976 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 22376 21131 22428 21140
rect 22376 21097 22385 21131
rect 22385 21097 22419 21131
rect 22419 21097 22428 21131
rect 22376 21088 22428 21097
rect 23848 21088 23900 21140
rect 24032 21088 24084 21140
rect 37832 21088 37884 21140
rect 12624 20884 12676 20936
rect 37924 20884 37976 20936
rect 23848 20816 23900 20868
rect 23204 20791 23256 20800
rect 23204 20757 23213 20791
rect 23213 20757 23247 20791
rect 23247 20757 23256 20791
rect 23204 20748 23256 20757
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 22192 20587 22244 20596
rect 22192 20553 22201 20587
rect 22201 20553 22235 20587
rect 22235 20553 22244 20587
rect 22192 20544 22244 20553
rect 23848 20544 23900 20596
rect 23204 20451 23256 20460
rect 23204 20417 23213 20451
rect 23213 20417 23247 20451
rect 23247 20417 23256 20451
rect 23204 20408 23256 20417
rect 31024 20408 31076 20460
rect 22008 20340 22060 20392
rect 20444 20272 20496 20324
rect 22744 20340 22796 20392
rect 38016 20315 38068 20324
rect 38016 20281 38025 20315
rect 38025 20281 38059 20315
rect 38059 20281 38068 20315
rect 38016 20272 38068 20281
rect 21824 20247 21876 20256
rect 21824 20213 21833 20247
rect 21833 20213 21867 20247
rect 21867 20213 21876 20247
rect 21824 20204 21876 20213
rect 22928 20204 22980 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 20904 20000 20956 20052
rect 23020 20000 23072 20052
rect 20444 19864 20496 19916
rect 20812 19839 20864 19848
rect 20812 19805 20821 19839
rect 20821 19805 20855 19839
rect 20855 19805 20864 19839
rect 20812 19796 20864 19805
rect 21824 19839 21876 19848
rect 21824 19805 21833 19839
rect 21833 19805 21867 19839
rect 21867 19805 21876 19839
rect 21824 19796 21876 19805
rect 37832 19839 37884 19848
rect 37832 19805 37841 19839
rect 37841 19805 37875 19839
rect 37875 19805 37884 19839
rect 37832 19796 37884 19805
rect 20720 19703 20772 19712
rect 20720 19669 20729 19703
rect 20729 19669 20763 19703
rect 20763 19669 20772 19703
rect 20720 19660 20772 19669
rect 21088 19660 21140 19712
rect 31024 19660 31076 19712
rect 38016 19703 38068 19712
rect 38016 19669 38025 19703
rect 38025 19669 38059 19703
rect 38059 19669 38068 19703
rect 38016 19660 38068 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 37832 19456 37884 19508
rect 20904 19388 20956 19440
rect 21088 19363 21140 19372
rect 21088 19329 21097 19363
rect 21097 19329 21131 19363
rect 21131 19329 21140 19363
rect 21088 19320 21140 19329
rect 34520 19320 34572 19372
rect 20168 19252 20220 19304
rect 20536 19295 20588 19304
rect 20536 19261 20545 19295
rect 20545 19261 20579 19295
rect 20579 19261 20588 19295
rect 20536 19252 20588 19261
rect 17960 19116 18012 19168
rect 38016 19159 38068 19168
rect 38016 19125 38025 19159
rect 38025 19125 38059 19159
rect 38059 19125 38068 19159
rect 38016 19116 38068 19125
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 19340 18776 19392 18828
rect 20444 18776 20496 18828
rect 20076 18708 20128 18760
rect 20168 18572 20220 18624
rect 37832 18751 37884 18760
rect 37832 18717 37841 18751
rect 37841 18717 37875 18751
rect 37875 18717 37884 18751
rect 37832 18708 37884 18717
rect 34520 18572 34572 18624
rect 38016 18615 38068 18624
rect 38016 18581 38025 18615
rect 38025 18581 38059 18615
rect 38059 18581 38068 18615
rect 38016 18572 38068 18581
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 18236 18411 18288 18420
rect 18236 18377 18245 18411
rect 18245 18377 18279 18411
rect 18279 18377 18288 18411
rect 18236 18368 18288 18377
rect 19432 18411 19484 18420
rect 19432 18377 19441 18411
rect 19441 18377 19475 18411
rect 19475 18377 19484 18411
rect 19432 18368 19484 18377
rect 18512 18164 18564 18216
rect 19340 18300 19392 18352
rect 20352 18164 20404 18216
rect 19340 18028 19392 18080
rect 37832 18028 37884 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 18236 17824 18288 17876
rect 19432 17824 19484 17876
rect 19340 17663 19392 17672
rect 19340 17629 19349 17663
rect 19349 17629 19383 17663
rect 19383 17629 19392 17663
rect 19340 17620 19392 17629
rect 38016 17527 38068 17536
rect 38016 17493 38025 17527
rect 38025 17493 38059 17527
rect 38059 17493 38068 17527
rect 38016 17484 38068 17493
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 18144 17187 18196 17196
rect 18144 17153 18153 17187
rect 18153 17153 18187 17187
rect 18187 17153 18196 17187
rect 18144 17144 18196 17153
rect 38016 16983 38068 16992
rect 38016 16949 38025 16983
rect 38025 16949 38059 16983
rect 38059 16949 38068 16983
rect 38016 16940 38068 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 18144 16736 18196 16788
rect 20904 16779 20956 16788
rect 20904 16745 20913 16779
rect 20913 16745 20947 16779
rect 20947 16745 20956 16779
rect 20904 16736 20956 16745
rect 17960 16668 18012 16720
rect 18144 16600 18196 16652
rect 20904 16532 20956 16584
rect 18052 16464 18104 16516
rect 20168 16507 20220 16516
rect 20168 16473 20177 16507
rect 20177 16473 20211 16507
rect 20211 16473 20220 16507
rect 20168 16464 20220 16473
rect 37280 16439 37332 16448
rect 37280 16405 37289 16439
rect 37289 16405 37323 16439
rect 37323 16405 37332 16439
rect 37280 16396 37332 16405
rect 38016 16439 38068 16448
rect 38016 16405 38025 16439
rect 38025 16405 38059 16439
rect 38059 16405 38068 16439
rect 38016 16396 38068 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 16212 15988 16264 16040
rect 17316 15988 17368 16040
rect 17868 15988 17920 16040
rect 17960 15920 18012 15972
rect 37280 16124 37332 16176
rect 37280 15895 37332 15904
rect 37280 15861 37289 15895
rect 37289 15861 37323 15895
rect 37323 15861 37332 15895
rect 37280 15852 37332 15861
rect 38016 15895 38068 15904
rect 38016 15861 38025 15895
rect 38025 15861 38059 15895
rect 38059 15861 38068 15895
rect 38016 15852 38068 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 17868 15691 17920 15700
rect 17868 15657 17877 15691
rect 17877 15657 17911 15691
rect 17911 15657 17920 15691
rect 17868 15648 17920 15657
rect 16212 15555 16264 15564
rect 16212 15521 16221 15555
rect 16221 15521 16255 15555
rect 16255 15521 16264 15555
rect 16212 15512 16264 15521
rect 16396 15487 16448 15496
rect 16396 15453 16405 15487
rect 16405 15453 16439 15487
rect 16439 15453 16448 15487
rect 16396 15444 16448 15453
rect 16120 15308 16172 15360
rect 37280 15308 37332 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 15752 15147 15804 15156
rect 15752 15113 15761 15147
rect 15761 15113 15795 15147
rect 15795 15113 15804 15147
rect 15752 15104 15804 15113
rect 16396 15104 16448 15156
rect 15384 14968 15436 15020
rect 15200 14900 15252 14952
rect 16212 14900 16264 14952
rect 38016 14875 38068 14884
rect 38016 14841 38025 14875
rect 38025 14841 38059 14875
rect 38059 14841 38068 14875
rect 38016 14832 38068 14841
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 15752 14560 15804 14612
rect 15200 14424 15252 14476
rect 15016 14399 15068 14408
rect 15016 14365 15025 14399
rect 15025 14365 15059 14399
rect 15059 14365 15068 14399
rect 15016 14356 15068 14365
rect 14832 14220 14884 14272
rect 38016 14263 38068 14272
rect 38016 14229 38025 14263
rect 38025 14229 38059 14263
rect 38059 14229 38068 14263
rect 38016 14220 38068 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 14924 14059 14976 14068
rect 14924 14025 14933 14059
rect 14933 14025 14967 14059
rect 14967 14025 14976 14059
rect 14924 14016 14976 14025
rect 15016 14016 15068 14068
rect 4712 13812 4764 13864
rect 15476 13880 15528 13932
rect 12072 13855 12124 13864
rect 12072 13821 12081 13855
rect 12081 13821 12115 13855
rect 12115 13821 12124 13855
rect 12072 13812 12124 13821
rect 38016 13719 38068 13728
rect 38016 13685 38025 13719
rect 38025 13685 38059 13719
rect 38059 13685 38068 13719
rect 38016 13676 38068 13685
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 12072 13515 12124 13524
rect 12072 13481 12081 13515
rect 12081 13481 12115 13515
rect 12115 13481 12124 13515
rect 12072 13472 12124 13481
rect 15476 13515 15528 13524
rect 15476 13481 15485 13515
rect 15485 13481 15519 13515
rect 15519 13481 15528 13515
rect 15476 13472 15528 13481
rect 12900 13404 12952 13456
rect 12624 13336 12676 13388
rect 13360 13336 13412 13388
rect 15108 13404 15160 13456
rect 14924 13336 14976 13388
rect 12900 13132 12952 13184
rect 14372 13175 14424 13184
rect 14372 13141 14381 13175
rect 14381 13141 14415 13175
rect 14415 13141 14424 13175
rect 14372 13132 14424 13141
rect 37280 13175 37332 13184
rect 37280 13141 37289 13175
rect 37289 13141 37323 13175
rect 37323 13141 37332 13175
rect 37280 13132 37332 13141
rect 38016 13175 38068 13184
rect 38016 13141 38025 13175
rect 38025 13141 38059 13175
rect 38059 13141 38068 13175
rect 38016 13132 38068 13141
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 12624 12971 12676 12980
rect 12624 12937 12633 12971
rect 12633 12937 12667 12971
rect 12667 12937 12676 12971
rect 12624 12928 12676 12937
rect 13544 12971 13596 12980
rect 13544 12937 13553 12971
rect 13553 12937 13587 12971
rect 13587 12937 13596 12971
rect 13544 12928 13596 12937
rect 13360 12767 13412 12776
rect 13360 12733 13369 12767
rect 13369 12733 13403 12767
rect 13403 12733 13412 12767
rect 13360 12724 13412 12733
rect 13636 12724 13688 12776
rect 37280 12588 37332 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 13360 12316 13412 12368
rect 12808 12291 12860 12300
rect 12808 12257 12817 12291
rect 12817 12257 12851 12291
rect 12851 12257 12860 12291
rect 12808 12248 12860 12257
rect 12992 12223 13044 12232
rect 12992 12189 13001 12223
rect 13001 12189 13035 12223
rect 13035 12189 13044 12223
rect 12992 12180 13044 12189
rect 13176 12112 13228 12164
rect 38016 12087 38068 12096
rect 38016 12053 38025 12087
rect 38025 12053 38059 12087
rect 38059 12053 38068 12087
rect 38016 12044 38068 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 12164 11883 12216 11892
rect 12164 11849 12173 11883
rect 12173 11849 12207 11883
rect 12207 11849 12216 11883
rect 12164 11840 12216 11849
rect 12808 11679 12860 11688
rect 12808 11645 12817 11679
rect 12817 11645 12851 11679
rect 12851 11645 12860 11679
rect 12808 11636 12860 11645
rect 13084 11636 13136 11688
rect 38016 11543 38068 11552
rect 38016 11509 38025 11543
rect 38025 11509 38059 11543
rect 38059 11509 38068 11543
rect 38016 11500 38068 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 11980 11339 12032 11348
rect 11980 11305 11989 11339
rect 11989 11305 12023 11339
rect 12023 11305 12032 11339
rect 11980 11296 12032 11305
rect 12808 11228 12860 11280
rect 38016 11271 38068 11280
rect 11980 11092 12032 11144
rect 38016 11237 38025 11271
rect 38025 11237 38059 11271
rect 38059 11237 38068 11271
rect 38016 11228 38068 11237
rect 2688 11024 2740 11076
rect 11336 11067 11388 11076
rect 11336 11033 11345 11067
rect 11345 11033 11379 11067
rect 11379 11033 11388 11067
rect 11336 11024 11388 11033
rect 13268 11024 13320 11076
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 10416 10795 10468 10804
rect 10416 10761 10425 10795
rect 10425 10761 10459 10795
rect 10459 10761 10468 10795
rect 10416 10752 10468 10761
rect 11336 10752 11388 10804
rect 10140 10684 10192 10736
rect 20168 10752 20220 10804
rect 10508 10616 10560 10668
rect 12624 10616 12676 10668
rect 12900 10659 12952 10668
rect 12900 10625 12909 10659
rect 12909 10625 12943 10659
rect 12943 10625 12952 10659
rect 12900 10616 12952 10625
rect 12440 10412 12492 10464
rect 13452 10412 13504 10464
rect 13728 10412 13780 10464
rect 37924 10684 37976 10736
rect 37280 10455 37332 10464
rect 37280 10421 37289 10455
rect 37289 10421 37323 10455
rect 37323 10421 37332 10455
rect 37280 10412 37332 10421
rect 38016 10455 38068 10464
rect 38016 10421 38025 10455
rect 38025 10421 38059 10455
rect 38059 10421 38068 10455
rect 38016 10412 38068 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 10140 10115 10192 10124
rect 10140 10081 10149 10115
rect 10149 10081 10183 10115
rect 10183 10081 10192 10115
rect 10140 10072 10192 10081
rect 12624 10072 12676 10124
rect 13728 10072 13780 10124
rect 10416 10047 10468 10056
rect 10416 10013 10425 10047
rect 10425 10013 10459 10047
rect 10459 10013 10468 10047
rect 10416 10004 10468 10013
rect 37280 10004 37332 10056
rect 3424 9936 3476 9988
rect 11980 9936 12032 9988
rect 10324 9911 10376 9920
rect 10324 9877 10333 9911
rect 10333 9877 10367 9911
rect 10367 9877 10376 9911
rect 10324 9868 10376 9877
rect 12532 9911 12584 9920
rect 12532 9877 12541 9911
rect 12541 9877 12575 9911
rect 12575 9877 12584 9911
rect 12532 9868 12584 9877
rect 12992 9911 13044 9920
rect 12992 9877 13001 9911
rect 13001 9877 13035 9911
rect 13035 9877 13044 9911
rect 12992 9868 13044 9877
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 10048 9596 10100 9648
rect 10140 9596 10192 9648
rect 11980 9639 12032 9648
rect 11980 9605 11989 9639
rect 11989 9605 12023 9639
rect 12023 9605 12032 9639
rect 11980 9596 12032 9605
rect 8208 9460 8260 9512
rect 12440 9528 12492 9580
rect 9496 9460 9548 9512
rect 12808 9503 12860 9512
rect 12808 9469 12817 9503
rect 12817 9469 12851 9503
rect 12851 9469 12860 9503
rect 12808 9460 12860 9469
rect 38016 9435 38068 9444
rect 38016 9401 38025 9435
rect 38025 9401 38059 9435
rect 38059 9401 38068 9435
rect 38016 9392 38068 9401
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 10048 9120 10100 9172
rect 12532 8984 12584 9036
rect 9588 8916 9640 8968
rect 12348 8959 12400 8968
rect 12348 8925 12357 8959
rect 12357 8925 12391 8959
rect 12391 8925 12400 8959
rect 12348 8916 12400 8925
rect 38016 8823 38068 8832
rect 38016 8789 38025 8823
rect 38025 8789 38059 8823
rect 38059 8789 38068 8823
rect 38016 8780 38068 8789
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 9220 8619 9272 8628
rect 9220 8585 9229 8619
rect 9229 8585 9263 8619
rect 9263 8585 9272 8619
rect 9220 8576 9272 8585
rect 9588 8619 9640 8628
rect 9588 8585 9597 8619
rect 9597 8585 9631 8619
rect 9631 8585 9640 8619
rect 9588 8576 9640 8585
rect 8208 8372 8260 8424
rect 9128 8415 9180 8424
rect 9128 8381 9137 8415
rect 9137 8381 9171 8415
rect 9171 8381 9180 8415
rect 9128 8372 9180 8381
rect 9772 8372 9824 8424
rect 9956 8304 10008 8356
rect 38016 8347 38068 8356
rect 38016 8313 38025 8347
rect 38025 8313 38059 8347
rect 38059 8313 38068 8347
rect 38016 8304 38068 8313
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 8944 8075 8996 8084
rect 8944 8041 8953 8075
rect 8953 8041 8987 8075
rect 8987 8041 8996 8075
rect 8944 8032 8996 8041
rect 8208 7896 8260 7948
rect 9772 7939 9824 7948
rect 9772 7905 9781 7939
rect 9781 7905 9815 7939
rect 9815 7905 9824 7939
rect 9772 7896 9824 7905
rect 8944 7828 8996 7880
rect 7932 7735 7984 7744
rect 7932 7701 7941 7735
rect 7941 7701 7975 7735
rect 7975 7701 7984 7735
rect 7932 7692 7984 7701
rect 37280 7735 37332 7744
rect 37280 7701 37289 7735
rect 37289 7701 37323 7735
rect 37323 7701 37332 7735
rect 37280 7692 37332 7701
rect 38016 7735 38068 7744
rect 38016 7701 38025 7735
rect 38025 7701 38059 7735
rect 38059 7701 38068 7735
rect 38016 7692 38068 7701
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 8024 7488 8076 7540
rect 7840 7284 7892 7336
rect 8208 7352 8260 7404
rect 8116 7327 8168 7336
rect 8116 7293 8125 7327
rect 8125 7293 8159 7327
rect 8159 7293 8168 7327
rect 8116 7284 8168 7293
rect 37280 7284 37332 7336
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 6552 6851 6604 6860
rect 6552 6817 6561 6851
rect 6561 6817 6595 6851
rect 6595 6817 6604 6851
rect 6552 6808 6604 6817
rect 7840 6851 7892 6860
rect 7840 6817 7849 6851
rect 7849 6817 7883 6851
rect 7883 6817 7892 6851
rect 7840 6808 7892 6817
rect 8944 6783 8996 6792
rect 8944 6749 8953 6783
rect 8953 6749 8987 6783
rect 8987 6749 8996 6783
rect 8944 6740 8996 6749
rect 10232 6783 10284 6792
rect 10232 6749 10241 6783
rect 10241 6749 10275 6783
rect 10275 6749 10284 6783
rect 10232 6740 10284 6749
rect 5172 6672 5224 6724
rect 37188 6672 37240 6724
rect 8392 6647 8444 6656
rect 8392 6613 8401 6647
rect 8401 6613 8435 6647
rect 8435 6613 8444 6647
rect 8392 6604 8444 6613
rect 38016 6647 38068 6656
rect 38016 6613 38025 6647
rect 38025 6613 38059 6647
rect 38059 6613 38068 6647
rect 38016 6604 38068 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 7104 6443 7156 6452
rect 7104 6409 7113 6443
rect 7113 6409 7147 6443
rect 7147 6409 7156 6443
rect 7104 6400 7156 6409
rect 8944 6400 8996 6452
rect 9956 6400 10008 6452
rect 37188 6400 37240 6452
rect 7012 6264 7064 6316
rect 8392 6264 8444 6316
rect 7748 6239 7800 6248
rect 7748 6205 7757 6239
rect 7757 6205 7791 6239
rect 7791 6205 7800 6239
rect 7748 6196 7800 6205
rect 37280 6196 37332 6248
rect 38016 6103 38068 6112
rect 38016 6069 38025 6103
rect 38025 6069 38059 6103
rect 38059 6069 38068 6103
rect 38016 6060 38068 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 6368 5856 6420 5908
rect 10232 5856 10284 5908
rect 37280 5899 37332 5908
rect 37280 5865 37289 5899
rect 37289 5865 37323 5899
rect 37323 5865 37332 5899
rect 37280 5856 37332 5865
rect 7748 5763 7800 5772
rect 7748 5729 7757 5763
rect 7757 5729 7791 5763
rect 7791 5729 7800 5763
rect 7748 5720 7800 5729
rect 8944 5695 8996 5704
rect 8944 5661 8953 5695
rect 8953 5661 8987 5695
rect 8987 5661 8996 5695
rect 8944 5652 8996 5661
rect 9220 5695 9272 5704
rect 9220 5661 9229 5695
rect 9229 5661 9263 5695
rect 9263 5661 9272 5695
rect 9220 5652 9272 5661
rect 7840 5559 7892 5568
rect 7840 5525 7849 5559
rect 7849 5525 7883 5559
rect 7883 5525 7892 5559
rect 7840 5516 7892 5525
rect 38016 5559 38068 5568
rect 38016 5525 38025 5559
rect 38025 5525 38059 5559
rect 38059 5525 38068 5559
rect 38016 5516 38068 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 4896 5312 4948 5364
rect 8944 5312 8996 5364
rect 9956 5312 10008 5364
rect 5540 5176 5592 5228
rect 7748 5151 7800 5160
rect 7748 5117 7757 5151
rect 7757 5117 7791 5151
rect 7791 5117 7800 5151
rect 9220 5176 9272 5228
rect 7748 5108 7800 5117
rect 38016 5015 38068 5024
rect 38016 4981 38025 5015
rect 38025 4981 38059 5015
rect 38059 4981 38068 5015
rect 38016 4972 38068 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 36728 4428 36780 4480
rect 37648 4428 37700 4480
rect 38016 4471 38068 4480
rect 38016 4437 38025 4471
rect 38025 4437 38059 4471
rect 38059 4437 38068 4471
rect 38016 4428 38068 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 38016 4199 38068 4208
rect 38016 4165 38025 4199
rect 38025 4165 38059 4199
rect 38059 4165 38068 4199
rect 38016 4156 38068 4165
rect 37924 4088 37976 4140
rect 12348 3952 12400 4004
rect 37832 3952 37884 4004
rect 34704 3927 34756 3936
rect 34704 3893 34713 3927
rect 34713 3893 34747 3927
rect 34747 3893 34756 3927
rect 34704 3884 34756 3893
rect 36176 3927 36228 3936
rect 36176 3893 36185 3927
rect 36185 3893 36219 3927
rect 36219 3893 36228 3927
rect 36176 3884 36228 3893
rect 36452 3884 36504 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 34796 3612 34848 3664
rect 36544 3587 36596 3596
rect 36544 3553 36553 3587
rect 36553 3553 36587 3587
rect 36587 3553 36596 3587
rect 36544 3544 36596 3553
rect 34704 3476 34756 3528
rect 36176 3476 36228 3528
rect 37832 3519 37884 3528
rect 37832 3485 37841 3519
rect 37841 3485 37875 3519
rect 37875 3485 37884 3519
rect 37832 3476 37884 3485
rect 5264 3383 5316 3392
rect 5264 3349 5273 3383
rect 5273 3349 5307 3383
rect 5307 3349 5316 3383
rect 5264 3340 5316 3349
rect 30288 3383 30340 3392
rect 30288 3349 30297 3383
rect 30297 3349 30331 3383
rect 30331 3349 30340 3383
rect 30288 3340 30340 3349
rect 31760 3340 31812 3392
rect 33048 3340 33100 3392
rect 38016 3383 38068 3392
rect 38016 3349 38025 3383
rect 38025 3349 38059 3383
rect 38059 3349 38068 3383
rect 38016 3340 38068 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 5540 3136 5592 3188
rect 9128 3136 9180 3188
rect 14372 3179 14424 3188
rect 14372 3145 14381 3179
rect 14381 3145 14415 3179
rect 14415 3145 14424 3179
rect 14372 3136 14424 3145
rect 22008 3179 22060 3188
rect 22008 3145 22017 3179
rect 22017 3145 22051 3179
rect 22051 3145 22060 3179
rect 22008 3136 22060 3145
rect 22928 3136 22980 3188
rect 26056 3136 26108 3188
rect 29092 3179 29144 3188
rect 29092 3145 29101 3179
rect 29101 3145 29135 3179
rect 29135 3145 29144 3179
rect 29092 3136 29144 3145
rect 12808 3068 12860 3120
rect 36452 3136 36504 3188
rect 37740 3136 37792 3188
rect 4620 3043 4672 3052
rect 4620 3009 4629 3043
rect 4629 3009 4663 3043
rect 4663 3009 4672 3043
rect 4620 3000 4672 3009
rect 8944 3000 8996 3052
rect 14096 3000 14148 3052
rect 21456 3000 21508 3052
rect 25872 3000 25924 3052
rect 28816 3000 28868 3052
rect 30656 3043 30708 3052
rect 30656 3009 30665 3043
rect 30665 3009 30699 3043
rect 30699 3009 30708 3043
rect 30656 3000 30708 3009
rect 32404 3043 32456 3052
rect 32404 3009 32413 3043
rect 32413 3009 32447 3043
rect 32447 3009 32456 3043
rect 32404 3000 32456 3009
rect 32588 3000 32640 3052
rect 34060 3000 34112 3052
rect 36452 3043 36504 3052
rect 36452 3009 36461 3043
rect 36461 3009 36495 3043
rect 36495 3009 36504 3043
rect 36452 3000 36504 3009
rect 37648 3000 37700 3052
rect 30288 2932 30340 2984
rect 31760 2932 31812 2984
rect 32496 2932 32548 2984
rect 33048 2932 33100 2984
rect 33968 2932 34020 2984
rect 3056 2796 3108 2848
rect 6000 2796 6052 2848
rect 6736 2839 6788 2848
rect 6736 2805 6745 2839
rect 6745 2805 6779 2839
rect 6779 2805 6788 2839
rect 6736 2796 6788 2805
rect 7472 2839 7524 2848
rect 7472 2805 7481 2839
rect 7481 2805 7515 2839
rect 7515 2805 7524 2839
rect 7472 2796 7524 2805
rect 9680 2796 9732 2848
rect 10416 2839 10468 2848
rect 10416 2805 10425 2839
rect 10425 2805 10459 2839
rect 10459 2805 10468 2839
rect 10416 2796 10468 2805
rect 10968 2839 11020 2848
rect 10968 2805 10977 2839
rect 10977 2805 11011 2839
rect 11011 2805 11020 2839
rect 10968 2796 11020 2805
rect 11888 2839 11940 2848
rect 11888 2805 11897 2839
rect 11897 2805 11931 2839
rect 11931 2805 11940 2839
rect 11888 2796 11940 2805
rect 12624 2839 12676 2848
rect 12624 2805 12633 2839
rect 12633 2805 12667 2839
rect 12667 2805 12676 2839
rect 12624 2796 12676 2805
rect 14924 2839 14976 2848
rect 14924 2805 14933 2839
rect 14933 2805 14967 2839
rect 14967 2805 14976 2839
rect 14924 2796 14976 2805
rect 15568 2839 15620 2848
rect 15568 2805 15577 2839
rect 15577 2805 15611 2839
rect 15611 2805 15620 2839
rect 15568 2796 15620 2805
rect 16304 2796 16356 2848
rect 17040 2839 17092 2848
rect 17040 2805 17049 2839
rect 17049 2805 17083 2839
rect 17083 2805 17092 2839
rect 17040 2796 17092 2805
rect 17776 2839 17828 2848
rect 17776 2805 17785 2839
rect 17785 2805 17819 2839
rect 17819 2805 17828 2839
rect 17776 2796 17828 2805
rect 18604 2839 18656 2848
rect 18604 2805 18613 2839
rect 18613 2805 18647 2839
rect 18647 2805 18656 2839
rect 18604 2796 18656 2805
rect 19248 2839 19300 2848
rect 19248 2805 19257 2839
rect 19257 2805 19291 2839
rect 19291 2805 19300 2839
rect 19248 2796 19300 2805
rect 19984 2839 20036 2848
rect 19984 2805 19993 2839
rect 19993 2805 20027 2839
rect 20027 2805 20036 2839
rect 19984 2796 20036 2805
rect 20812 2796 20864 2848
rect 24216 2839 24268 2848
rect 24216 2805 24225 2839
rect 24225 2805 24259 2839
rect 24259 2805 24268 2839
rect 24216 2796 24268 2805
rect 24400 2796 24452 2848
rect 25044 2796 25096 2848
rect 26976 2839 27028 2848
rect 26976 2805 26985 2839
rect 26985 2805 27019 2839
rect 27019 2805 27028 2839
rect 26976 2796 27028 2805
rect 27620 2839 27672 2848
rect 27620 2805 27629 2839
rect 27629 2805 27663 2839
rect 27663 2805 27672 2839
rect 27620 2796 27672 2805
rect 33232 2796 33284 2848
rect 34612 2796 34664 2848
rect 36636 2839 36688 2848
rect 36636 2805 36645 2839
rect 36645 2805 36679 2839
rect 36679 2805 36688 2839
rect 36636 2796 36688 2805
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 5172 2635 5224 2644
rect 5172 2601 5181 2635
rect 5181 2601 5215 2635
rect 5215 2601 5224 2635
rect 5172 2592 5224 2601
rect 7840 2592 7892 2644
rect 7932 2592 7984 2644
rect 9496 2635 9548 2644
rect 9496 2601 9505 2635
rect 9505 2601 9539 2635
rect 9539 2601 9548 2635
rect 9496 2592 9548 2601
rect 10324 2635 10376 2644
rect 10324 2601 10333 2635
rect 10333 2601 10367 2635
rect 10367 2601 10376 2635
rect 10324 2592 10376 2601
rect 13176 2592 13228 2644
rect 13636 2592 13688 2644
rect 14832 2635 14884 2644
rect 14832 2601 14841 2635
rect 14841 2601 14875 2635
rect 14875 2601 14884 2635
rect 14832 2592 14884 2601
rect 15384 2592 15436 2644
rect 16120 2635 16172 2644
rect 16120 2601 16129 2635
rect 16129 2601 16163 2635
rect 16163 2601 16172 2635
rect 16120 2592 16172 2601
rect 17316 2635 17368 2644
rect 17316 2601 17325 2635
rect 17325 2601 17359 2635
rect 17359 2601 17368 2635
rect 17316 2592 17368 2601
rect 18144 2592 18196 2644
rect 18512 2635 18564 2644
rect 18512 2601 18521 2635
rect 18521 2601 18555 2635
rect 18555 2601 18564 2635
rect 18512 2592 18564 2601
rect 20076 2635 20128 2644
rect 20076 2601 20085 2635
rect 20085 2601 20119 2635
rect 20119 2601 20128 2635
rect 20076 2592 20128 2601
rect 20720 2592 20772 2644
rect 23296 2592 23348 2644
rect 24584 2635 24636 2644
rect 24584 2601 24593 2635
rect 24593 2601 24627 2635
rect 24627 2601 24636 2635
rect 24584 2592 24636 2601
rect 25228 2635 25280 2644
rect 25228 2601 25237 2635
rect 25237 2601 25271 2635
rect 25271 2601 25280 2635
rect 25228 2592 25280 2601
rect 26240 2592 26292 2644
rect 27160 2635 27212 2644
rect 27160 2601 27169 2635
rect 27169 2601 27203 2635
rect 27203 2601 27212 2635
rect 27160 2592 27212 2601
rect 27804 2635 27856 2644
rect 27804 2601 27813 2635
rect 27813 2601 27847 2635
rect 27847 2601 27856 2635
rect 27804 2592 27856 2601
rect 28448 2635 28500 2644
rect 28448 2601 28457 2635
rect 28457 2601 28491 2635
rect 28491 2601 28500 2635
rect 28448 2592 28500 2601
rect 36544 2635 36596 2644
rect 36544 2601 36553 2635
rect 36553 2601 36587 2635
rect 36587 2601 36596 2635
rect 36544 2592 36596 2601
rect 5080 2524 5132 2576
rect 6920 2524 6972 2576
rect 7012 2567 7064 2576
rect 7012 2533 7021 2567
rect 7021 2533 7055 2567
rect 7055 2533 7064 2567
rect 7012 2524 7064 2533
rect 8116 2524 8168 2576
rect 13084 2524 13136 2576
rect 20352 2524 20404 2576
rect 35440 2524 35492 2576
rect 12992 2456 13044 2508
rect 30564 2456 30616 2508
rect 32312 2456 32364 2508
rect 33692 2456 33744 2508
rect 2320 2388 2372 2440
rect 3056 2431 3108 2440
rect 3056 2397 3065 2431
rect 3065 2397 3099 2431
rect 3099 2397 3108 2431
rect 3056 2388 3108 2397
rect 4896 2388 4948 2440
rect 5264 2388 5316 2440
rect 6000 2388 6052 2440
rect 6736 2388 6788 2440
rect 7472 2388 7524 2440
rect 8300 2388 8352 2440
rect 9680 2431 9732 2440
rect 9680 2397 9689 2431
rect 9689 2397 9723 2431
rect 9723 2397 9732 2431
rect 9680 2388 9732 2397
rect 10416 2388 10468 2440
rect 10968 2388 11020 2440
rect 11888 2388 11940 2440
rect 12624 2388 12676 2440
rect 13360 2431 13412 2440
rect 13360 2397 13369 2431
rect 13369 2397 13403 2431
rect 13403 2397 13412 2431
rect 13360 2388 13412 2397
rect 14832 2388 14884 2440
rect 15568 2388 15620 2440
rect 16304 2388 16356 2440
rect 17040 2388 17092 2440
rect 17776 2388 17828 2440
rect 18512 2388 18564 2440
rect 19340 2431 19392 2440
rect 19340 2397 19349 2431
rect 19349 2397 19383 2431
rect 19383 2397 19392 2431
rect 19340 2388 19392 2397
rect 19984 2388 20036 2440
rect 20720 2388 20772 2440
rect 22928 2388 22980 2440
rect 23020 2431 23072 2440
rect 23020 2397 23029 2431
rect 23029 2397 23063 2431
rect 23063 2397 23072 2431
rect 23020 2388 23072 2397
rect 23756 2388 23808 2440
rect 24216 2388 24268 2440
rect 25044 2431 25096 2440
rect 25044 2397 25053 2431
rect 25053 2397 25087 2431
rect 25087 2397 25096 2431
rect 25044 2388 25096 2397
rect 25136 2388 25188 2440
rect 26608 2388 26660 2440
rect 26976 2431 27028 2440
rect 26976 2397 26985 2431
rect 26985 2397 27019 2431
rect 27019 2397 27028 2431
rect 26976 2388 27028 2397
rect 27620 2431 27672 2440
rect 27620 2397 27629 2431
rect 27629 2397 27663 2431
rect 27663 2397 27672 2431
rect 27620 2388 27672 2397
rect 28080 2388 28132 2440
rect 29552 2388 29604 2440
rect 10508 2320 10560 2372
rect 3792 2252 3844 2304
rect 6920 2252 6972 2304
rect 13452 2320 13504 2372
rect 13268 2252 13320 2304
rect 22192 2252 22244 2304
rect 31024 2252 31076 2304
rect 34612 2388 34664 2440
rect 36728 2431 36780 2440
rect 36728 2397 36737 2431
rect 36737 2397 36771 2431
rect 36771 2397 36780 2431
rect 36728 2388 36780 2397
rect 35532 2320 35584 2372
rect 33968 2252 34020 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 2318 39200 2374 40000
rect 3054 39200 3110 40000
rect 3790 39200 3846 40000
rect 4526 39200 4582 40000
rect 5262 39200 5318 40000
rect 5998 39200 6054 40000
rect 6734 39200 6790 40000
rect 7470 39200 7526 40000
rect 8206 39200 8262 40000
rect 8942 39200 8998 40000
rect 9678 39200 9734 40000
rect 10414 39200 10470 40000
rect 11150 39200 11206 40000
rect 11886 39200 11942 40000
rect 12622 39200 12678 40000
rect 13358 39200 13414 40000
rect 14094 39200 14150 40000
rect 14830 39200 14886 40000
rect 15566 39200 15622 40000
rect 16302 39200 16358 40000
rect 17038 39200 17094 40000
rect 17774 39200 17830 40000
rect 18510 39200 18566 40000
rect 19246 39200 19302 40000
rect 19982 39200 20038 40000
rect 20718 39200 20774 40000
rect 21454 39200 21510 40000
rect 22190 39200 22246 40000
rect 22926 39200 22982 40000
rect 23662 39200 23718 40000
rect 24398 39200 24454 40000
rect 24504 39222 24808 39250
rect 2332 37330 2360 39200
rect 2320 37324 2372 37330
rect 2320 37266 2372 37272
rect 2688 37256 2740 37262
rect 2688 37198 2740 37204
rect 2700 11082 2728 37198
rect 3068 36786 3096 39200
rect 3804 37126 3832 39200
rect 4540 37754 4568 39200
rect 4540 37726 4660 37754
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 3792 37120 3844 37126
rect 3792 37062 3844 37068
rect 4632 36786 4660 37726
rect 5276 37330 5304 39200
rect 5264 37324 5316 37330
rect 5264 37266 5316 37272
rect 4988 37256 5040 37262
rect 4988 37198 5040 37204
rect 3056 36780 3108 36786
rect 3056 36722 3108 36728
rect 4620 36780 4672 36786
rect 4620 36722 4672 36728
rect 3424 36712 3476 36718
rect 3424 36654 3476 36660
rect 2688 11076 2740 11082
rect 2688 11018 2740 11024
rect 3436 9994 3464 36654
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4632 36378 4660 36722
rect 4896 36712 4948 36718
rect 4896 36654 4948 36660
rect 4620 36372 4672 36378
rect 4620 36314 4672 36320
rect 4712 36372 4764 36378
rect 4712 36314 4764 36320
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4724 13870 4752 36314
rect 4712 13864 4764 13870
rect 4712 13806 4764 13812
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 3424 9988 3476 9994
rect 3424 9930 3476 9936
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4908 5370 4936 36654
rect 5000 36378 5028 37198
rect 4988 36372 5040 36378
rect 4988 36314 5040 36320
rect 6012 36242 6040 39200
rect 6552 37256 6604 37262
rect 6552 37198 6604 37204
rect 6000 36236 6052 36242
rect 6000 36178 6052 36184
rect 6368 36168 6420 36174
rect 6368 36110 6420 36116
rect 5172 6724 5224 6730
rect 5172 6666 5224 6672
rect 4896 5364 4948 5370
rect 4896 5306 4948 5312
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 3056 2848 3108 2854
rect 3056 2790 3108 2796
rect 3068 2446 3096 2790
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 2320 2440 2372 2446
rect 2320 2382 2372 2388
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 2332 800 2360 2382
rect 3068 800 3096 2382
rect 3792 2304 3844 2310
rect 3792 2246 3844 2252
rect 3804 800 3832 2246
rect 4632 1986 4660 2994
rect 5184 2650 5212 6666
rect 6380 5914 6408 36110
rect 6564 6866 6592 37198
rect 6748 36786 6776 39200
rect 7484 37330 7512 39200
rect 7472 37324 7524 37330
rect 7472 37266 7524 37272
rect 8024 37256 8076 37262
rect 8024 37198 8076 37204
rect 6736 36780 6788 36786
rect 6736 36722 6788 36728
rect 6748 36378 6776 36722
rect 7104 36712 7156 36718
rect 7104 36654 7156 36660
rect 6736 36372 6788 36378
rect 6736 36314 6788 36320
rect 6552 6860 6604 6866
rect 6552 6802 6604 6808
rect 7116 6458 7144 36654
rect 7932 7744 7984 7750
rect 7932 7686 7984 7692
rect 7840 7336 7892 7342
rect 7840 7278 7892 7284
rect 7852 6866 7880 7278
rect 7840 6860 7892 6866
rect 7760 6820 7840 6848
rect 7104 6452 7156 6458
rect 7104 6394 7156 6400
rect 7012 6316 7064 6322
rect 7012 6258 7064 6264
rect 6368 5908 6420 5914
rect 6368 5850 6420 5856
rect 5540 5228 5592 5234
rect 5540 5170 5592 5176
rect 5264 3392 5316 3398
rect 5264 3334 5316 3340
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5080 2576 5132 2582
rect 4908 2524 5080 2530
rect 4908 2518 5132 2524
rect 4908 2502 5120 2518
rect 4908 2446 4936 2502
rect 5276 2446 5304 3334
rect 5552 3194 5580 5170
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 6000 2848 6052 2854
rect 6000 2790 6052 2796
rect 6736 2848 6788 2854
rect 6736 2790 6788 2796
rect 6012 2446 6040 2790
rect 6748 2446 6776 2790
rect 7024 2582 7052 6258
rect 7760 6254 7788 6820
rect 7840 6802 7892 6808
rect 7748 6248 7800 6254
rect 7748 6190 7800 6196
rect 7760 5778 7788 6190
rect 7748 5772 7800 5778
rect 7748 5714 7800 5720
rect 7760 5166 7788 5714
rect 7840 5568 7892 5574
rect 7840 5510 7892 5516
rect 7748 5160 7800 5166
rect 7748 5102 7800 5108
rect 7472 2848 7524 2854
rect 7472 2790 7524 2796
rect 6920 2576 6972 2582
rect 6920 2518 6972 2524
rect 7012 2576 7064 2582
rect 7012 2518 7064 2524
rect 4896 2440 4948 2446
rect 4896 2382 4948 2388
rect 5264 2440 5316 2446
rect 5264 2382 5316 2388
rect 6000 2440 6052 2446
rect 6000 2382 6052 2388
rect 6736 2440 6788 2446
rect 6736 2382 6788 2388
rect 4540 1958 4660 1986
rect 4540 800 4568 1958
rect 5276 800 5304 2382
rect 6012 800 6040 2382
rect 6748 800 6776 2382
rect 6932 2310 6960 2518
rect 7484 2446 7512 2790
rect 7852 2650 7880 5510
rect 7944 2650 7972 7686
rect 8036 7546 8064 37198
rect 8220 36786 8248 39200
rect 8208 36780 8260 36786
rect 8208 36722 8260 36728
rect 8220 36378 8248 36722
rect 8852 36712 8904 36718
rect 8852 36654 8904 36660
rect 8208 36372 8260 36378
rect 8208 36314 8260 36320
rect 8864 26234 8892 36654
rect 8956 36242 8984 39200
rect 9692 36786 9720 39200
rect 10428 37398 10456 39200
rect 10416 37392 10468 37398
rect 10416 37334 10468 37340
rect 10416 37256 10468 37262
rect 10416 37198 10468 37204
rect 9680 36780 9732 36786
rect 9680 36722 9732 36728
rect 9692 36378 9720 36722
rect 10048 36712 10100 36718
rect 10048 36654 10100 36660
rect 9680 36372 9732 36378
rect 9680 36314 9732 36320
rect 8944 36236 8996 36242
rect 8944 36178 8996 36184
rect 8956 35834 8984 36178
rect 9220 36168 9272 36174
rect 9220 36110 9272 36116
rect 8944 35828 8996 35834
rect 8944 35770 8996 35776
rect 8864 26206 8984 26234
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 8220 8430 8248 9454
rect 8208 8424 8260 8430
rect 8208 8366 8260 8372
rect 8220 7954 8248 8366
rect 8956 8090 8984 26206
rect 9232 8634 9260 36110
rect 10060 9654 10088 36654
rect 10428 10810 10456 37198
rect 11164 36786 11192 39200
rect 11900 37330 11928 39200
rect 11888 37324 11940 37330
rect 11888 37266 11940 37272
rect 11152 36780 11204 36786
rect 11152 36722 11204 36728
rect 11164 36378 11192 36722
rect 11900 36378 11928 37266
rect 12164 37256 12216 37262
rect 12164 37198 12216 37204
rect 11980 36712 12032 36718
rect 11980 36654 12032 36660
rect 11152 36372 11204 36378
rect 11152 36314 11204 36320
rect 11888 36372 11940 36378
rect 11888 36314 11940 36320
rect 11992 11354 12020 36654
rect 12072 13864 12124 13870
rect 12072 13806 12124 13812
rect 12084 13530 12112 13806
rect 12072 13524 12124 13530
rect 12072 13466 12124 13472
rect 12176 11898 12204 37198
rect 12636 36786 12664 39200
rect 13372 37262 13400 39200
rect 13360 37256 13412 37262
rect 13360 37198 13412 37204
rect 13544 37120 13596 37126
rect 13544 37062 13596 37068
rect 12624 36780 12676 36786
rect 12624 36722 12676 36728
rect 12636 36378 12664 36722
rect 12992 36576 13044 36582
rect 12992 36518 13044 36524
rect 12624 36372 12676 36378
rect 12624 36314 12676 36320
rect 12624 20936 12676 20942
rect 12624 20878 12676 20884
rect 12636 13394 12664 20878
rect 12900 13456 12952 13462
rect 12900 13398 12952 13404
rect 12624 13388 12676 13394
rect 12624 13330 12676 13336
rect 12636 12986 12664 13330
rect 12912 13190 12940 13398
rect 12900 13184 12952 13190
rect 12900 13126 12952 13132
rect 12624 12980 12676 12986
rect 12624 12922 12676 12928
rect 12164 11892 12216 11898
rect 12164 11834 12216 11840
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 11992 11150 12020 11290
rect 11980 11144 12032 11150
rect 11980 11086 12032 11092
rect 11336 11076 11388 11082
rect 11336 11018 11388 11024
rect 11348 10810 11376 11018
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 11336 10804 11388 10810
rect 11336 10746 11388 10752
rect 10140 10736 10192 10742
rect 10140 10678 10192 10684
rect 10152 10130 10180 10678
rect 10140 10124 10192 10130
rect 10140 10066 10192 10072
rect 10152 9654 10180 10066
rect 10428 10062 10456 10746
rect 12636 10674 12664 12922
rect 12808 12300 12860 12306
rect 12808 12242 12860 12248
rect 12820 11694 12848 12242
rect 12808 11688 12860 11694
rect 12808 11630 12860 11636
rect 12820 11286 12848 11630
rect 12808 11280 12860 11286
rect 12808 11222 12860 11228
rect 12912 10674 12940 13126
rect 13004 12238 13032 36518
rect 13360 13388 13412 13394
rect 13360 13330 13412 13336
rect 13372 12782 13400 13330
rect 13556 12986 13584 37062
rect 14108 36786 14136 39200
rect 14844 37262 14872 39200
rect 15580 37262 15608 39200
rect 16316 37262 16344 39200
rect 17052 37262 17080 39200
rect 17788 37262 17816 39200
rect 18524 37262 18552 39200
rect 19260 37262 19288 39200
rect 19996 37262 20024 39200
rect 20732 37262 20760 39200
rect 14832 37256 14884 37262
rect 14832 37198 14884 37204
rect 15568 37256 15620 37262
rect 15568 37198 15620 37204
rect 16304 37256 16356 37262
rect 16304 37198 16356 37204
rect 17040 37256 17092 37262
rect 17040 37198 17092 37204
rect 17776 37256 17828 37262
rect 17776 37198 17828 37204
rect 18512 37256 18564 37262
rect 18512 37198 18564 37204
rect 19248 37256 19300 37262
rect 19248 37198 19300 37204
rect 19984 37256 20036 37262
rect 19984 37198 20036 37204
rect 20720 37256 20772 37262
rect 20720 37198 20772 37204
rect 14844 36922 14872 37198
rect 15016 37120 15068 37126
rect 15016 37062 15068 37068
rect 14832 36916 14884 36922
rect 14832 36858 14884 36864
rect 14096 36780 14148 36786
rect 14096 36722 14148 36728
rect 14832 36576 14884 36582
rect 14832 36518 14884 36524
rect 14844 35894 14872 36518
rect 14844 35866 14964 35894
rect 14832 14272 14884 14278
rect 14832 14214 14884 14220
rect 14372 13184 14424 13190
rect 14372 13126 14424 13132
rect 13544 12980 13596 12986
rect 13544 12922 13596 12928
rect 13360 12776 13412 12782
rect 13360 12718 13412 12724
rect 13636 12776 13688 12782
rect 13636 12718 13688 12724
rect 13372 12374 13400 12718
rect 13360 12368 13412 12374
rect 13360 12310 13412 12316
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 13176 12164 13228 12170
rect 13176 12106 13228 12112
rect 13084 11688 13136 11694
rect 13084 11630 13136 11636
rect 10508 10668 10560 10674
rect 10508 10610 10560 10616
rect 12624 10668 12676 10674
rect 12624 10610 12676 10616
rect 12900 10668 12952 10674
rect 12900 10610 12952 10616
rect 10416 10056 10468 10062
rect 10416 9998 10468 10004
rect 10324 9920 10376 9926
rect 10324 9862 10376 9868
rect 10048 9648 10100 9654
rect 10048 9590 10100 9596
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9128 8424 9180 8430
rect 9128 8366 9180 8372
rect 8944 8084 8996 8090
rect 8944 8026 8996 8032
rect 8208 7948 8260 7954
rect 8208 7890 8260 7896
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 8220 7410 8248 7890
rect 8956 7886 8984 8026
rect 8944 7880 8996 7886
rect 8944 7822 8996 7828
rect 8208 7404 8260 7410
rect 8208 7346 8260 7352
rect 8116 7336 8168 7342
rect 8116 7278 8168 7284
rect 7840 2644 7892 2650
rect 7840 2586 7892 2592
rect 7932 2644 7984 2650
rect 7932 2586 7984 2592
rect 8128 2582 8156 7278
rect 8944 6792 8996 6798
rect 8944 6734 8996 6740
rect 8392 6656 8444 6662
rect 8392 6598 8444 6604
rect 8404 6322 8432 6598
rect 8956 6458 8984 6734
rect 8944 6452 8996 6458
rect 8944 6394 8996 6400
rect 8392 6316 8444 6322
rect 8392 6258 8444 6264
rect 8944 5704 8996 5710
rect 8944 5646 8996 5652
rect 8956 5370 8984 5646
rect 8944 5364 8996 5370
rect 8944 5306 8996 5312
rect 9140 3194 9168 8366
rect 9220 5704 9272 5710
rect 9220 5646 9272 5652
rect 9232 5234 9260 5646
rect 9220 5228 9272 5234
rect 9220 5170 9272 5176
rect 9128 3188 9180 3194
rect 9128 3130 9180 3136
rect 8944 3052 8996 3058
rect 8944 2994 8996 3000
rect 8116 2576 8168 2582
rect 8116 2518 8168 2524
rect 7472 2440 7524 2446
rect 8300 2440 8352 2446
rect 7472 2382 7524 2388
rect 8220 2400 8300 2428
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 7484 800 7512 2382
rect 8220 800 8248 2400
rect 8300 2382 8352 2388
rect 8956 800 8984 2994
rect 9508 2650 9536 9454
rect 10060 9178 10088 9590
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 9588 8968 9640 8974
rect 9588 8910 9640 8916
rect 9600 8634 9628 8910
rect 9588 8628 9640 8634
rect 9588 8570 9640 8576
rect 9772 8424 9824 8430
rect 9772 8366 9824 8372
rect 9784 7954 9812 8366
rect 9956 8356 10008 8362
rect 9956 8298 10008 8304
rect 9772 7948 9824 7954
rect 9772 7890 9824 7896
rect 9968 6458 9996 8298
rect 10232 6792 10284 6798
rect 10232 6734 10284 6740
rect 9956 6452 10008 6458
rect 9956 6394 10008 6400
rect 9968 5370 9996 6394
rect 10244 5914 10272 6734
rect 10232 5908 10284 5914
rect 10232 5850 10284 5856
rect 9956 5364 10008 5370
rect 9956 5306 10008 5312
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9496 2644 9548 2650
rect 9496 2586 9548 2592
rect 9692 2446 9720 2790
rect 10336 2650 10364 9862
rect 10416 2848 10468 2854
rect 10416 2790 10468 2796
rect 10324 2644 10376 2650
rect 10324 2586 10376 2592
rect 10428 2446 10456 2790
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 10416 2440 10468 2446
rect 10416 2382 10468 2388
rect 9692 800 9720 2382
rect 10428 800 10456 2382
rect 10520 2378 10548 10610
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 11980 9988 12032 9994
rect 11980 9930 12032 9936
rect 11992 9654 12020 9930
rect 11980 9648 12032 9654
rect 11980 9590 12032 9596
rect 12452 9586 12480 10406
rect 12636 10130 12664 10610
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12532 9920 12584 9926
rect 12532 9862 12584 9868
rect 12992 9920 13044 9926
rect 12992 9862 13044 9868
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12544 9042 12572 9862
rect 12808 9512 12860 9518
rect 12808 9454 12860 9460
rect 12532 9036 12584 9042
rect 12532 8978 12584 8984
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12360 4010 12388 8910
rect 12348 4004 12400 4010
rect 12348 3946 12400 3952
rect 12820 3126 12848 9454
rect 12808 3120 12860 3126
rect 12808 3062 12860 3068
rect 10968 2848 11020 2854
rect 10968 2790 11020 2796
rect 11888 2848 11940 2854
rect 11888 2790 11940 2796
rect 12624 2848 12676 2854
rect 12624 2790 12676 2796
rect 10980 2446 11008 2790
rect 11900 2446 11928 2790
rect 12636 2446 12664 2790
rect 13004 2514 13032 9862
rect 13096 2582 13124 11630
rect 13188 2650 13216 12106
rect 13268 11076 13320 11082
rect 13268 11018 13320 11024
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 13084 2576 13136 2582
rect 13084 2518 13136 2524
rect 12992 2508 13044 2514
rect 12992 2450 13044 2456
rect 10968 2440 11020 2446
rect 11888 2440 11940 2446
rect 11020 2400 11192 2428
rect 10968 2382 11020 2388
rect 10508 2372 10560 2378
rect 10508 2314 10560 2320
rect 11164 800 11192 2400
rect 11888 2382 11940 2388
rect 12624 2440 12676 2446
rect 12624 2382 12676 2388
rect 11900 800 11928 2382
rect 12636 800 12664 2382
rect 13280 2310 13308 11018
rect 13452 10464 13504 10470
rect 13452 10406 13504 10412
rect 13360 2440 13412 2446
rect 13360 2382 13412 2388
rect 13268 2304 13320 2310
rect 13268 2246 13320 2252
rect 13372 800 13400 2382
rect 13464 2378 13492 10406
rect 13648 2650 13676 12718
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 10130 13768 10406
rect 13728 10124 13780 10130
rect 13728 10066 13780 10072
rect 14384 3194 14412 13126
rect 14372 3188 14424 3194
rect 14372 3130 14424 3136
rect 14096 3052 14148 3058
rect 14096 2994 14148 3000
rect 13636 2644 13688 2650
rect 13636 2586 13688 2592
rect 13452 2372 13504 2378
rect 13452 2314 13504 2320
rect 14108 800 14136 2994
rect 14844 2650 14872 14214
rect 14936 14074 14964 35866
rect 15028 14414 15056 37062
rect 15580 36922 15608 37198
rect 15752 37120 15804 37126
rect 15752 37062 15804 37068
rect 15568 36916 15620 36922
rect 15568 36858 15620 36864
rect 15764 15162 15792 37062
rect 16316 36922 16344 37198
rect 16396 37120 16448 37126
rect 16396 37062 16448 37068
rect 16304 36916 16356 36922
rect 16304 36858 16356 36864
rect 16212 16040 16264 16046
rect 16212 15982 16264 15988
rect 16224 15570 16252 15982
rect 16212 15564 16264 15570
rect 16212 15506 16264 15512
rect 16120 15360 16172 15366
rect 16120 15302 16172 15308
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15200 14952 15252 14958
rect 15200 14894 15252 14900
rect 15212 14482 15240 14894
rect 15200 14476 15252 14482
rect 15200 14418 15252 14424
rect 15016 14408 15068 14414
rect 15016 14350 15068 14356
rect 15028 14074 15056 14350
rect 14924 14068 14976 14074
rect 14924 14010 14976 14016
rect 15016 14068 15068 14074
rect 15016 14010 15068 14016
rect 14936 13394 14964 14010
rect 15212 13818 15240 14418
rect 15120 13790 15240 13818
rect 15120 13462 15148 13790
rect 15108 13456 15160 13462
rect 15108 13398 15160 13404
rect 14924 13388 14976 13394
rect 14924 13330 14976 13336
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 14832 2644 14884 2650
rect 14832 2586 14884 2592
rect 14832 2440 14884 2446
rect 14936 2428 14964 2790
rect 15396 2650 15424 14962
rect 15764 14618 15792 15098
rect 15752 14612 15804 14618
rect 15752 14554 15804 14560
rect 15476 13932 15528 13938
rect 15476 13874 15528 13880
rect 15488 13530 15516 13874
rect 15476 13524 15528 13530
rect 15476 13466 15528 13472
rect 15568 2848 15620 2854
rect 15568 2790 15620 2796
rect 15384 2644 15436 2650
rect 15384 2586 15436 2592
rect 15580 2446 15608 2790
rect 16132 2650 16160 15302
rect 16224 14958 16252 15506
rect 16408 15502 16436 37062
rect 17052 36922 17080 37198
rect 17788 36922 17816 37198
rect 17868 37120 17920 37126
rect 17868 37062 17920 37068
rect 18052 37120 18104 37126
rect 18052 37062 18104 37068
rect 18236 37120 18288 37126
rect 18236 37062 18288 37068
rect 17040 36916 17092 36922
rect 17040 36858 17092 36864
rect 17776 36916 17828 36922
rect 17776 36858 17828 36864
rect 17880 16046 17908 37062
rect 17960 19168 18012 19174
rect 17960 19110 18012 19116
rect 17972 16726 18000 19110
rect 17960 16720 18012 16726
rect 17960 16662 18012 16668
rect 17316 16040 17368 16046
rect 17316 15982 17368 15988
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16408 15162 16436 15438
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 16212 14952 16264 14958
rect 16212 14894 16264 14900
rect 16304 2848 16356 2854
rect 16304 2790 16356 2796
rect 17040 2848 17092 2854
rect 17040 2790 17092 2796
rect 16120 2644 16172 2650
rect 16120 2586 16172 2592
rect 16316 2446 16344 2790
rect 17052 2446 17080 2790
rect 17328 2650 17356 15982
rect 17880 15706 17908 15982
rect 17972 15978 18000 16662
rect 18064 16522 18092 37062
rect 18248 18426 18276 37062
rect 18524 36922 18552 37198
rect 19260 36922 19288 37198
rect 19432 37120 19484 37126
rect 19432 37062 19484 37068
rect 18512 36916 18564 36922
rect 18512 36858 18564 36864
rect 19248 36916 19300 36922
rect 19248 36858 19300 36864
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 18236 18420 18288 18426
rect 18236 18362 18288 18368
rect 18248 17882 18276 18362
rect 19352 18358 19380 18770
rect 19444 18426 19472 37062
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19996 36922 20024 37198
rect 20536 37120 20588 37126
rect 20536 37062 20588 37068
rect 19984 36916 20036 36922
rect 19984 36858 20036 36864
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30427 19882 30436
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24987 19882 24996
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 20260 22228 20312 22234
rect 20260 22170 20312 22176
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 20168 19304 20220 19310
rect 20168 19246 20220 19252
rect 20076 18760 20128 18766
rect 20076 18702 20128 18708
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 19432 18420 19484 18426
rect 19432 18362 19484 18368
rect 19340 18352 19392 18358
rect 19340 18294 19392 18300
rect 18512 18216 18564 18222
rect 18512 18158 18564 18164
rect 18236 17876 18288 17882
rect 18236 17818 18288 17824
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 18156 16794 18184 17138
rect 18144 16788 18196 16794
rect 18144 16730 18196 16736
rect 18144 16652 18196 16658
rect 18144 16594 18196 16600
rect 18052 16516 18104 16522
rect 18052 16458 18104 16464
rect 17960 15972 18012 15978
rect 17960 15914 18012 15920
rect 17868 15700 17920 15706
rect 17868 15642 17920 15648
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 17316 2644 17368 2650
rect 17316 2586 17368 2592
rect 17788 2446 17816 2790
rect 18156 2650 18184 16594
rect 18524 2650 18552 18158
rect 19340 18080 19392 18086
rect 19340 18022 19392 18028
rect 19352 17678 19380 18022
rect 19444 17882 19472 18362
rect 19432 17876 19484 17882
rect 19432 17818 19484 17824
rect 19340 17672 19392 17678
rect 19340 17614 19392 17620
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 18604 2848 18656 2854
rect 18604 2790 18656 2796
rect 19248 2848 19300 2854
rect 19248 2790 19300 2796
rect 19984 2848 20036 2854
rect 19984 2790 20036 2796
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 14884 2400 14964 2428
rect 15568 2440 15620 2446
rect 14832 2382 14884 2388
rect 15568 2382 15620 2388
rect 16304 2440 16356 2446
rect 16304 2382 16356 2388
rect 17040 2440 17092 2446
rect 17040 2382 17092 2388
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 18512 2440 18564 2446
rect 18616 2428 18644 2790
rect 18564 2400 18644 2428
rect 19260 2428 19288 2790
rect 19996 2446 20024 2790
rect 20088 2650 20116 18702
rect 20180 18630 20208 19246
rect 20168 18624 20220 18630
rect 20168 18566 20220 18572
rect 20272 18442 20300 22170
rect 20444 20324 20496 20330
rect 20444 20266 20496 20272
rect 20456 19922 20484 20266
rect 20444 19916 20496 19922
rect 20444 19858 20496 19864
rect 20456 18834 20484 19858
rect 20548 19310 20576 37062
rect 20732 36922 20760 37198
rect 20812 37120 20864 37126
rect 20812 37062 20864 37068
rect 20720 36916 20772 36922
rect 20720 36858 20772 36864
rect 20824 19854 20852 37062
rect 21468 36786 21496 39200
rect 22204 37126 22232 39200
rect 22940 37262 22968 39200
rect 22284 37256 22336 37262
rect 22284 37198 22336 37204
rect 22928 37256 22980 37262
rect 22928 37198 22980 37204
rect 22192 37120 22244 37126
rect 22192 37062 22244 37068
rect 21456 36780 21508 36786
rect 21456 36722 21508 36728
rect 22192 36576 22244 36582
rect 22192 36518 22244 36524
rect 22204 20602 22232 36518
rect 22296 21894 22324 37198
rect 22836 37120 22888 37126
rect 22836 37062 22888 37068
rect 22744 22568 22796 22574
rect 22744 22510 22796 22516
rect 22376 22024 22428 22030
rect 22376 21966 22428 21972
rect 22284 21888 22336 21894
rect 22284 21830 22336 21836
rect 22388 21146 22416 21966
rect 22756 21486 22784 22510
rect 22848 21690 22876 37062
rect 23676 36922 23704 39200
rect 24412 39114 24440 39200
rect 24504 39114 24532 39222
rect 24412 39086 24532 39114
rect 24584 37256 24636 37262
rect 24780 37244 24808 39222
rect 25134 39200 25190 40000
rect 25870 39200 25926 40000
rect 26606 39200 26662 40000
rect 27342 39200 27398 40000
rect 28078 39200 28134 40000
rect 28814 39200 28870 40000
rect 29550 39200 29606 40000
rect 30286 39200 30342 40000
rect 31022 39200 31078 40000
rect 31758 39200 31814 40000
rect 32494 39200 32550 40000
rect 33230 39200 33286 40000
rect 33966 39200 34022 40000
rect 34072 39222 34468 39250
rect 25148 37330 25176 39200
rect 25136 37324 25188 37330
rect 25136 37266 25188 37272
rect 24860 37256 24912 37262
rect 24780 37216 24860 37244
rect 24584 37198 24636 37204
rect 24860 37198 24912 37204
rect 23756 37120 23808 37126
rect 23756 37062 23808 37068
rect 23664 36916 23716 36922
rect 23664 36858 23716 36864
rect 23020 23588 23072 23594
rect 23020 23530 23072 23536
rect 23032 23118 23060 23530
rect 23112 23180 23164 23186
rect 23112 23122 23164 23128
rect 23020 23112 23072 23118
rect 23020 23054 23072 23060
rect 22836 21684 22888 21690
rect 22836 21626 22888 21632
rect 22744 21480 22796 21486
rect 22744 21422 22796 21428
rect 22376 21140 22428 21146
rect 22376 21082 22428 21088
rect 22192 20596 22244 20602
rect 22192 20538 22244 20544
rect 22756 20398 22784 21422
rect 22008 20392 22060 20398
rect 22008 20334 22060 20340
rect 22744 20392 22796 20398
rect 22744 20334 22796 20340
rect 21824 20256 21876 20262
rect 21824 20198 21876 20204
rect 20904 20052 20956 20058
rect 20904 19994 20956 20000
rect 20812 19848 20864 19854
rect 20812 19790 20864 19796
rect 20720 19712 20772 19718
rect 20720 19654 20772 19660
rect 20536 19304 20588 19310
rect 20536 19246 20588 19252
rect 20444 18828 20496 18834
rect 20444 18770 20496 18776
rect 20180 18414 20300 18442
rect 20180 16522 20208 18414
rect 20352 18216 20404 18222
rect 20352 18158 20404 18164
rect 20168 16516 20220 16522
rect 20168 16458 20220 16464
rect 20180 10810 20208 16458
rect 20168 10804 20220 10810
rect 20168 10746 20220 10752
rect 20076 2644 20128 2650
rect 20076 2586 20128 2592
rect 20364 2582 20392 18158
rect 20732 2650 20760 19654
rect 20916 19446 20944 19994
rect 21836 19854 21864 20198
rect 21824 19848 21876 19854
rect 21824 19790 21876 19796
rect 21088 19712 21140 19718
rect 21088 19654 21140 19660
rect 20904 19440 20956 19446
rect 20904 19382 20956 19388
rect 20916 16794 20944 19382
rect 21100 19378 21128 19654
rect 21088 19372 21140 19378
rect 21088 19314 21140 19320
rect 20904 16788 20956 16794
rect 20904 16730 20956 16736
rect 20916 16590 20944 16730
rect 20904 16584 20956 16590
rect 20904 16526 20956 16532
rect 22020 3194 22048 20334
rect 22928 20256 22980 20262
rect 22928 20198 22980 20204
rect 22940 3194 22968 20198
rect 23032 20058 23060 23054
rect 23124 22982 23152 23122
rect 23112 22976 23164 22982
rect 23112 22918 23164 22924
rect 23124 22574 23152 22918
rect 23768 22778 23796 37062
rect 24596 36922 24624 37198
rect 24768 37120 24820 37126
rect 24768 37062 24820 37068
rect 24584 36916 24636 36922
rect 24584 36858 24636 36864
rect 23848 28144 23900 28150
rect 23848 28086 23900 28092
rect 23756 22772 23808 22778
rect 23756 22714 23808 22720
rect 23112 22568 23164 22574
rect 23112 22510 23164 22516
rect 23296 21888 23348 21894
rect 23296 21830 23348 21836
rect 23308 21486 23336 21830
rect 23296 21480 23348 21486
rect 23296 21422 23348 21428
rect 23204 20800 23256 20806
rect 23204 20742 23256 20748
rect 23216 20466 23244 20742
rect 23204 20460 23256 20466
rect 23204 20402 23256 20408
rect 23020 20052 23072 20058
rect 23020 19994 23072 20000
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 22928 3188 22980 3194
rect 22928 3130 22980 3136
rect 21456 3052 21508 3058
rect 21456 2994 21508 3000
rect 20812 2848 20864 2854
rect 20812 2790 20864 2796
rect 20720 2644 20772 2650
rect 20720 2586 20772 2592
rect 20352 2576 20404 2582
rect 20352 2518 20404 2524
rect 19340 2440 19392 2446
rect 19260 2400 19340 2428
rect 18512 2382 18564 2388
rect 14844 800 14872 2382
rect 15580 800 15608 2382
rect 16316 800 16344 2382
rect 17052 800 17080 2382
rect 17788 800 17816 2382
rect 18524 800 18552 2382
rect 19260 800 19288 2400
rect 19340 2382 19392 2388
rect 19984 2440 20036 2446
rect 19984 2382 20036 2388
rect 20720 2440 20772 2446
rect 20824 2428 20852 2790
rect 20772 2400 20852 2428
rect 20720 2382 20772 2388
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 19996 800 20024 2382
rect 20732 800 20760 2382
rect 21468 800 21496 2994
rect 22940 2446 22968 3130
rect 23308 2650 23336 21422
rect 23860 21146 23888 28086
rect 24492 24268 24544 24274
rect 24492 24210 24544 24216
rect 24504 23662 24532 24210
rect 24492 23656 24544 23662
rect 24492 23598 24544 23604
rect 24504 23186 24532 23598
rect 24492 23180 24544 23186
rect 24492 23122 24544 23128
rect 24780 23118 24808 37062
rect 24872 36922 24900 37198
rect 25320 37120 25372 37126
rect 25320 37062 25372 37068
rect 24860 36916 24912 36922
rect 24860 36858 24912 36864
rect 25332 23866 25360 37062
rect 25884 36922 25912 39200
rect 26620 37262 26648 39200
rect 27356 37262 27384 39200
rect 28092 37262 28120 39200
rect 26608 37256 26660 37262
rect 26608 37198 26660 37204
rect 26976 37256 27028 37262
rect 26976 37198 27028 37204
rect 27344 37256 27396 37262
rect 27344 37198 27396 37204
rect 27620 37256 27672 37262
rect 27620 37198 27672 37204
rect 28080 37256 28132 37262
rect 28080 37198 28132 37204
rect 26988 36922 27016 37198
rect 27344 37120 27396 37126
rect 27344 37062 27396 37068
rect 27528 37120 27580 37126
rect 27528 37062 27580 37068
rect 25872 36916 25924 36922
rect 25872 36858 25924 36864
rect 26976 36916 27028 36922
rect 26976 36858 27028 36864
rect 25780 36576 25832 36582
rect 25780 36518 25832 36524
rect 25792 24206 25820 36518
rect 27356 26042 27384 37062
rect 27344 26036 27396 26042
rect 27344 25978 27396 25984
rect 27160 25968 27212 25974
rect 27160 25910 27212 25916
rect 26792 24812 26844 24818
rect 26792 24754 26844 24760
rect 26056 24608 26108 24614
rect 26056 24550 26108 24556
rect 25780 24200 25832 24206
rect 25780 24142 25832 24148
rect 26068 24070 26096 24550
rect 26804 24410 26832 24754
rect 26792 24404 26844 24410
rect 26792 24346 26844 24352
rect 26056 24064 26108 24070
rect 26056 24006 26108 24012
rect 25320 23860 25372 23866
rect 25320 23802 25372 23808
rect 25228 23180 25280 23186
rect 25228 23122 25280 23128
rect 24768 23112 24820 23118
rect 24768 23054 24820 23060
rect 24584 22500 24636 22506
rect 24584 22442 24636 22448
rect 24596 21894 24624 22442
rect 25240 22438 25268 23122
rect 25228 22432 25280 22438
rect 25228 22374 25280 22380
rect 25320 22432 25372 22438
rect 25320 22374 25372 22380
rect 24584 21888 24636 21894
rect 24584 21830 24636 21836
rect 24032 21344 24084 21350
rect 24032 21286 24084 21292
rect 24044 21146 24072 21286
rect 23848 21140 23900 21146
rect 23848 21082 23900 21088
rect 24032 21140 24084 21146
rect 24032 21082 24084 21088
rect 23860 20874 23888 21082
rect 23848 20868 23900 20874
rect 23848 20810 23900 20816
rect 23860 20602 23888 20810
rect 23848 20596 23900 20602
rect 23848 20538 23900 20544
rect 24216 2848 24268 2854
rect 24216 2790 24268 2796
rect 24400 2848 24452 2854
rect 24400 2790 24452 2796
rect 23296 2644 23348 2650
rect 23296 2586 23348 2592
rect 24228 2446 24256 2790
rect 22928 2440 22980 2446
rect 22928 2382 22980 2388
rect 23020 2440 23072 2446
rect 23756 2440 23808 2446
rect 23020 2382 23072 2388
rect 23676 2400 23756 2428
rect 22192 2304 22244 2310
rect 22192 2246 22244 2252
rect 22204 800 22232 2246
rect 23032 1578 23060 2382
rect 22940 1550 23060 1578
rect 22940 800 22968 1550
rect 23676 800 23704 2400
rect 23756 2382 23808 2388
rect 24216 2440 24268 2446
rect 24216 2382 24268 2388
rect 24412 800 24440 2790
rect 24596 2650 24624 21830
rect 25044 2848 25096 2854
rect 25044 2790 25096 2796
rect 24584 2644 24636 2650
rect 24584 2586 24636 2592
rect 25056 2446 25084 2790
rect 25240 2650 25268 22374
rect 25332 22234 25360 22374
rect 25320 22228 25372 22234
rect 25320 22170 25372 22176
rect 26068 3194 26096 24006
rect 26240 23656 26292 23662
rect 26240 23598 26292 23604
rect 26252 22982 26280 23598
rect 26240 22976 26292 22982
rect 26240 22918 26292 22924
rect 26056 3188 26108 3194
rect 26056 3130 26108 3136
rect 25872 3052 25924 3058
rect 25872 2994 25924 3000
rect 25228 2644 25280 2650
rect 25228 2586 25280 2592
rect 25044 2440 25096 2446
rect 25044 2382 25096 2388
rect 25136 2440 25188 2446
rect 25136 2382 25188 2388
rect 25148 800 25176 2382
rect 25884 800 25912 2994
rect 26252 2650 26280 22918
rect 26976 2848 27028 2854
rect 26976 2790 27028 2796
rect 26240 2644 26292 2650
rect 26240 2586 26292 2592
rect 26988 2446 27016 2790
rect 27172 2650 27200 25910
rect 27540 25294 27568 37062
rect 27632 36922 27660 37198
rect 28264 37120 28316 37126
rect 28264 37062 28316 37068
rect 28724 37120 28776 37126
rect 28724 37062 28776 37068
rect 27620 36916 27672 36922
rect 27620 36858 27672 36864
rect 28172 28076 28224 28082
rect 28172 28018 28224 28024
rect 27988 26920 28040 26926
rect 27988 26862 28040 26868
rect 28000 26450 28028 26862
rect 27988 26444 28040 26450
rect 27988 26386 28040 26392
rect 27896 25900 27948 25906
rect 27896 25842 27948 25848
rect 27712 25696 27764 25702
rect 27712 25638 27764 25644
rect 27724 25294 27752 25638
rect 27908 25498 27936 25842
rect 28000 25770 28028 26386
rect 27988 25764 28040 25770
rect 27988 25706 28040 25712
rect 27896 25492 27948 25498
rect 27896 25434 27948 25440
rect 28000 25362 28028 25706
rect 27988 25356 28040 25362
rect 27988 25298 28040 25304
rect 27528 25288 27580 25294
rect 27528 25230 27580 25236
rect 27712 25288 27764 25294
rect 27712 25230 27764 25236
rect 27804 25152 27856 25158
rect 27804 25094 27856 25100
rect 27816 24614 27844 25094
rect 27804 24608 27856 24614
rect 27804 24550 27856 24556
rect 27620 2848 27672 2854
rect 27620 2790 27672 2796
rect 27160 2644 27212 2650
rect 27160 2586 27212 2592
rect 27632 2446 27660 2790
rect 27816 2650 27844 24550
rect 28184 23594 28212 28018
rect 28276 26382 28304 37062
rect 28736 27130 28764 37062
rect 28828 35834 28856 39200
rect 29368 37256 29420 37262
rect 29368 37198 29420 37204
rect 29380 36582 29408 37198
rect 29564 36922 29592 39200
rect 30012 37256 30064 37262
rect 30300 37244 30328 39200
rect 30472 37256 30524 37262
rect 30300 37216 30472 37244
rect 30012 37198 30064 37204
rect 30472 37198 30524 37204
rect 29644 37120 29696 37126
rect 29644 37062 29696 37068
rect 29552 36916 29604 36922
rect 29552 36858 29604 36864
rect 29368 36576 29420 36582
rect 29368 36518 29420 36524
rect 29380 35834 29408 36518
rect 28816 35828 28868 35834
rect 28816 35770 28868 35776
rect 29368 35828 29420 35834
rect 29368 35770 29420 35776
rect 29656 28218 29684 37062
rect 30024 36922 30052 37198
rect 30380 37120 30432 37126
rect 30380 37062 30432 37068
rect 30012 36916 30064 36922
rect 30012 36858 30064 36864
rect 30196 29708 30248 29714
rect 30196 29650 30248 29656
rect 30208 29102 30236 29650
rect 30196 29096 30248 29102
rect 30196 29038 30248 29044
rect 30208 28626 30236 29038
rect 30196 28620 30248 28626
rect 30196 28562 30248 28568
rect 29644 28212 29696 28218
rect 29644 28154 29696 28160
rect 28816 28076 28868 28082
rect 28816 28018 28868 28024
rect 28828 27674 28856 28018
rect 29184 28008 29236 28014
rect 29184 27950 29236 27956
rect 28816 27668 28868 27674
rect 28816 27610 28868 27616
rect 28724 27124 28776 27130
rect 28724 27066 28776 27072
rect 29196 26994 29224 27950
rect 30208 27946 30236 28562
rect 30392 28558 30420 37062
rect 31036 36922 31064 39200
rect 31772 37262 31800 39200
rect 32508 37262 32536 39200
rect 33244 37262 33272 39200
rect 33980 39114 34008 39200
rect 34072 39114 34100 39222
rect 33980 39086 34100 39114
rect 31760 37256 31812 37262
rect 31760 37198 31812 37204
rect 32220 37256 32272 37262
rect 32220 37198 32272 37204
rect 32496 37256 32548 37262
rect 32496 37198 32548 37204
rect 33232 37256 33284 37262
rect 33232 37198 33284 37204
rect 34440 37210 34468 39222
rect 34702 39200 34758 40000
rect 35438 39200 35494 40000
rect 35544 39222 35848 39250
rect 34716 37330 34744 39200
rect 35452 39114 35480 39200
rect 35544 39114 35572 39222
rect 35452 39086 35572 39114
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 34704 37324 34756 37330
rect 34532 37262 34560 37293
rect 34704 37266 34756 37272
rect 34520 37256 34572 37262
rect 34440 37204 34520 37210
rect 34440 37198 34572 37204
rect 35820 37210 35848 39222
rect 36174 39200 36230 40000
rect 36910 39200 36966 40000
rect 37646 39200 37702 40000
rect 36188 37466 36216 39200
rect 36176 37460 36228 37466
rect 36176 37402 36228 37408
rect 35900 37256 35952 37262
rect 35820 37204 35900 37210
rect 35820 37198 35952 37204
rect 32128 37120 32180 37126
rect 32128 37062 32180 37068
rect 31024 36916 31076 36922
rect 31024 36858 31076 36864
rect 31116 36576 31168 36582
rect 31116 36518 31168 36524
rect 31128 29306 31156 36518
rect 31668 32224 31720 32230
rect 31668 32166 31720 32172
rect 31116 29300 31168 29306
rect 31116 29242 31168 29248
rect 30656 28620 30708 28626
rect 30656 28562 30708 28568
rect 30380 28552 30432 28558
rect 30380 28494 30432 28500
rect 30472 28008 30524 28014
rect 30472 27950 30524 27956
rect 30196 27940 30248 27946
rect 30196 27882 30248 27888
rect 29920 27872 29972 27878
rect 29920 27814 29972 27820
rect 29932 27470 29960 27814
rect 30484 27538 30512 27950
rect 30472 27532 30524 27538
rect 30472 27474 30524 27480
rect 29920 27464 29972 27470
rect 29920 27406 29972 27412
rect 29184 26988 29236 26994
rect 29184 26930 29236 26936
rect 29092 26920 29144 26926
rect 29092 26862 29144 26868
rect 28264 26376 28316 26382
rect 28264 26318 28316 26324
rect 28448 26308 28500 26314
rect 28448 26250 28500 26256
rect 28172 23588 28224 23594
rect 28172 23530 28224 23536
rect 28460 2650 28488 26250
rect 28540 26240 28592 26246
rect 28540 26182 28592 26188
rect 28552 25906 28580 26182
rect 28540 25900 28592 25906
rect 28540 25842 28592 25848
rect 29104 3194 29132 26862
rect 30484 26234 30512 27474
rect 30484 26206 30604 26234
rect 30288 3392 30340 3398
rect 30288 3334 30340 3340
rect 29092 3188 29144 3194
rect 29092 3130 29144 3136
rect 28816 3052 28868 3058
rect 28816 2994 28868 3000
rect 27804 2644 27856 2650
rect 27804 2586 27856 2592
rect 28448 2644 28500 2650
rect 28448 2586 28500 2592
rect 26608 2440 26660 2446
rect 26608 2382 26660 2388
rect 26976 2440 27028 2446
rect 26976 2382 27028 2388
rect 27620 2440 27672 2446
rect 27620 2382 27672 2388
rect 28080 2440 28132 2446
rect 28080 2382 28132 2388
rect 26620 800 26648 2382
rect 27632 1986 27660 2382
rect 27356 1958 27660 1986
rect 27356 800 27384 1958
rect 28092 800 28120 2382
rect 28828 800 28856 2994
rect 30300 2990 30328 3334
rect 30288 2984 30340 2990
rect 30288 2926 30340 2932
rect 29552 2440 29604 2446
rect 29552 2382 29604 2388
rect 29564 800 29592 2382
rect 30300 800 30328 2926
rect 30576 2514 30604 26206
rect 30668 3058 30696 28562
rect 31680 28150 31708 32166
rect 32140 29646 32168 37062
rect 32232 36922 32260 37198
rect 32508 36922 32536 37198
rect 34440 37182 34560 37198
rect 32588 37120 32640 37126
rect 32588 37062 32640 37068
rect 33416 37120 33468 37126
rect 33416 37062 33468 37068
rect 33784 37120 33836 37126
rect 33784 37062 33836 37068
rect 32220 36916 32272 36922
rect 32220 36858 32272 36864
rect 32496 36916 32548 36922
rect 32496 36858 32548 36864
rect 32496 30592 32548 30598
rect 32496 30534 32548 30540
rect 32508 30190 32536 30534
rect 32600 30326 32628 37062
rect 32588 30320 32640 30326
rect 32588 30262 32640 30268
rect 32312 30184 32364 30190
rect 32312 30126 32364 30132
rect 32496 30184 32548 30190
rect 32496 30126 32548 30132
rect 32324 29714 32352 30126
rect 32312 29708 32364 29714
rect 32312 29650 32364 29656
rect 32128 29640 32180 29646
rect 32128 29582 32180 29588
rect 32404 29572 32456 29578
rect 32404 29514 32456 29520
rect 32312 29096 32364 29102
rect 32312 29038 32364 29044
rect 32324 28422 32352 29038
rect 32312 28416 32364 28422
rect 32312 28358 32364 28364
rect 31668 28144 31720 28150
rect 31668 28086 31720 28092
rect 31024 20460 31076 20466
rect 31024 20402 31076 20408
rect 31036 19718 31064 20402
rect 31024 19712 31076 19718
rect 31024 19654 31076 19660
rect 31760 3392 31812 3398
rect 31760 3334 31812 3340
rect 30656 3052 30708 3058
rect 30656 2994 30708 3000
rect 31772 2990 31800 3334
rect 31760 2984 31812 2990
rect 31760 2926 31812 2932
rect 30564 2508 30616 2514
rect 30564 2450 30616 2456
rect 31024 2304 31076 2310
rect 31024 2246 31076 2252
rect 31036 800 31064 2246
rect 31772 800 31800 2926
rect 32324 2514 32352 28358
rect 32416 3058 32444 29514
rect 32508 16574 32536 30126
rect 33428 29646 33456 37062
rect 33600 31884 33652 31890
rect 33600 31826 33652 31832
rect 33612 31210 33640 31826
rect 33796 31754 33824 37062
rect 34532 36922 34560 37182
rect 35820 37182 35940 37198
rect 34796 37120 34848 37126
rect 34796 37062 34848 37068
rect 35532 37120 35584 37126
rect 35532 37062 35584 37068
rect 34520 36916 34572 36922
rect 34520 36858 34572 36864
rect 34520 33312 34572 33318
rect 34520 33254 34572 33260
rect 34532 32978 34560 33254
rect 34520 32972 34572 32978
rect 34520 32914 34572 32920
rect 34532 32366 34560 32914
rect 34808 32570 34836 37062
rect 35348 36712 35400 36718
rect 35348 36654 35400 36660
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35360 36378 35388 36654
rect 35348 36372 35400 36378
rect 35348 36314 35400 36320
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35440 34944 35492 34950
rect 35440 34886 35492 34892
rect 35452 34746 35480 34886
rect 35440 34740 35492 34746
rect 35440 34682 35492 34688
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35544 32910 35572 37062
rect 35820 35834 35848 37182
rect 36188 36786 36216 37402
rect 36452 37256 36504 37262
rect 36452 37198 36504 37204
rect 36268 36916 36320 36922
rect 36268 36858 36320 36864
rect 36176 36780 36228 36786
rect 36176 36722 36228 36728
rect 36174 36680 36230 36689
rect 36174 36615 36230 36624
rect 36188 36174 36216 36615
rect 36176 36168 36228 36174
rect 36176 36110 36228 36116
rect 35992 36032 36044 36038
rect 35992 35974 36044 35980
rect 35808 35828 35860 35834
rect 35808 35770 35860 35776
rect 35900 35488 35952 35494
rect 35900 35430 35952 35436
rect 35912 34950 35940 35430
rect 35900 34944 35952 34950
rect 35900 34886 35952 34892
rect 35912 34066 35940 34886
rect 36004 34610 36032 35974
rect 36188 35834 36216 36110
rect 36176 35828 36228 35834
rect 36176 35770 36228 35776
rect 35992 34604 36044 34610
rect 35992 34546 36044 34552
rect 35900 34060 35952 34066
rect 35900 34002 35952 34008
rect 35532 32904 35584 32910
rect 35532 32846 35584 32852
rect 35440 32836 35492 32842
rect 35440 32778 35492 32784
rect 34796 32564 34848 32570
rect 34796 32506 34848 32512
rect 34520 32360 34572 32366
rect 34520 32302 34572 32308
rect 34704 32360 34756 32366
rect 34704 32302 34756 32308
rect 34716 32026 34744 32302
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34704 32020 34756 32026
rect 34704 31962 34756 31968
rect 34716 31754 34744 31962
rect 33784 31748 33836 31754
rect 34716 31726 34836 31754
rect 33784 31690 33836 31696
rect 33968 31680 34020 31686
rect 33968 31622 34020 31628
rect 33600 31204 33652 31210
rect 33652 31164 33732 31192
rect 33600 31146 33652 31152
rect 33508 30252 33560 30258
rect 33508 30194 33560 30200
rect 33520 29850 33548 30194
rect 33508 29844 33560 29850
rect 33508 29786 33560 29792
rect 33416 29640 33468 29646
rect 33416 29582 33468 29588
rect 33508 29640 33560 29646
rect 33508 29582 33560 29588
rect 32772 29504 32824 29510
rect 32772 29446 32824 29452
rect 32784 29170 32812 29446
rect 33520 29306 33548 29582
rect 33600 29504 33652 29510
rect 33600 29446 33652 29452
rect 33508 29300 33560 29306
rect 33508 29242 33560 29248
rect 32772 29164 32824 29170
rect 32772 29106 32824 29112
rect 33612 29034 33640 29446
rect 33600 29028 33652 29034
rect 33600 28970 33652 28976
rect 33612 16574 33640 28970
rect 33704 28218 33732 31164
rect 33980 31142 34008 31622
rect 34612 31340 34664 31346
rect 34612 31282 34664 31288
rect 33968 31136 34020 31142
rect 33968 31078 34020 31084
rect 33692 28212 33744 28218
rect 33692 28154 33744 28160
rect 33980 16574 34008 31078
rect 34520 30728 34572 30734
rect 34520 30670 34572 30676
rect 34152 30252 34204 30258
rect 34152 30194 34204 30200
rect 34164 29102 34192 30194
rect 34532 30122 34560 30670
rect 34520 30116 34572 30122
rect 34520 30058 34572 30064
rect 34624 30054 34652 31282
rect 34612 30048 34664 30054
rect 34612 29990 34664 29996
rect 34152 29096 34204 29102
rect 34152 29038 34204 29044
rect 34520 19372 34572 19378
rect 34520 19314 34572 19320
rect 34532 18630 34560 19314
rect 34520 18624 34572 18630
rect 34520 18566 34572 18572
rect 32508 16546 32628 16574
rect 33612 16546 33732 16574
rect 33980 16546 34100 16574
rect 32600 3058 32628 16546
rect 33048 3392 33100 3398
rect 33048 3334 33100 3340
rect 32404 3052 32456 3058
rect 32404 2994 32456 3000
rect 32588 3052 32640 3058
rect 32588 2994 32640 3000
rect 33060 2990 33088 3334
rect 32496 2984 32548 2990
rect 32496 2926 32548 2932
rect 33048 2984 33100 2990
rect 33048 2926 33100 2932
rect 32312 2508 32364 2514
rect 32312 2450 32364 2456
rect 32508 800 32536 2926
rect 33232 2848 33284 2854
rect 33232 2790 33284 2796
rect 33244 800 33272 2790
rect 33704 2514 33732 16546
rect 34072 3058 34100 16546
rect 34704 3936 34756 3942
rect 34704 3878 34756 3884
rect 34716 3534 34744 3878
rect 34808 3670 34836 31726
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35452 16574 35480 32778
rect 35912 31210 35940 34002
rect 36280 33998 36308 36858
rect 36360 36644 36412 36650
rect 36360 36586 36412 36592
rect 36268 33992 36320 33998
rect 36268 33934 36320 33940
rect 35992 33312 36044 33318
rect 35992 33254 36044 33260
rect 36004 32842 36032 33254
rect 35992 32836 36044 32842
rect 35992 32778 36044 32784
rect 35900 31204 35952 31210
rect 35900 31146 35952 31152
rect 36372 22778 36400 36586
rect 36464 36106 36492 37198
rect 36924 36922 36952 39200
rect 36912 36916 36964 36922
rect 36912 36858 36964 36864
rect 36544 36780 36596 36786
rect 36544 36722 36596 36728
rect 36452 36100 36504 36106
rect 36452 36042 36504 36048
rect 36464 35494 36492 36042
rect 36452 35488 36504 35494
rect 36452 35430 36504 35436
rect 36556 34746 36584 36722
rect 37660 36718 37688 39200
rect 38106 37360 38162 37369
rect 38106 37295 38162 37304
rect 38016 37120 38068 37126
rect 38016 37062 38068 37068
rect 37648 36712 37700 36718
rect 37648 36654 37700 36660
rect 37188 36644 37240 36650
rect 37188 36586 37240 36592
rect 36728 35692 36780 35698
rect 36728 35634 36780 35640
rect 36544 34740 36596 34746
rect 36544 34682 36596 34688
rect 36452 33856 36504 33862
rect 36452 33798 36504 33804
rect 36544 33856 36596 33862
rect 36544 33798 36596 33804
rect 36464 26234 36492 33798
rect 36556 33522 36584 33798
rect 36740 33658 36768 35634
rect 37096 35556 37148 35562
rect 37096 35498 37148 35504
rect 36820 35080 36872 35086
rect 36820 35022 36872 35028
rect 36728 33652 36780 33658
rect 36728 33594 36780 33600
rect 36544 33516 36596 33522
rect 36544 33458 36596 33464
rect 36464 26206 36584 26234
rect 36360 22772 36412 22778
rect 36360 22714 36412 22720
rect 35452 16546 35572 16574
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 34796 3664 34848 3670
rect 34796 3606 34848 3612
rect 34704 3528 34756 3534
rect 34704 3470 34756 3476
rect 34060 3052 34112 3058
rect 34060 2994 34112 3000
rect 33968 2984 34020 2990
rect 33968 2926 34020 2932
rect 33692 2508 33744 2514
rect 33692 2450 33744 2456
rect 33980 2310 34008 2926
rect 34612 2848 34664 2854
rect 34612 2790 34664 2796
rect 34624 2446 34652 2790
rect 34612 2440 34664 2446
rect 34612 2382 34664 2388
rect 33968 2304 34020 2310
rect 33968 2246 34020 2252
rect 33980 800 34008 2246
rect 34716 800 34744 3470
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 35440 2576 35492 2582
rect 35440 2518 35492 2524
rect 35452 800 35480 2518
rect 35544 2378 35572 16546
rect 36176 3936 36228 3942
rect 36176 3878 36228 3884
rect 36452 3936 36504 3942
rect 36452 3878 36504 3884
rect 36188 3534 36216 3878
rect 36176 3528 36228 3534
rect 36176 3470 36228 3476
rect 35532 2372 35584 2378
rect 35532 2314 35584 2320
rect 36188 800 36216 3470
rect 36464 3194 36492 3878
rect 36556 3602 36584 26206
rect 36832 23322 36860 35022
rect 37004 34944 37056 34950
rect 37004 34886 37056 34892
rect 37016 34649 37044 34886
rect 37002 34640 37058 34649
rect 37002 34575 37058 34584
rect 37108 33969 37136 35498
rect 37200 35329 37228 36586
rect 37464 36576 37516 36582
rect 37464 36518 37516 36524
rect 37186 35320 37242 35329
rect 37186 35255 37242 35264
rect 37476 33998 37504 36518
rect 37832 36168 37884 36174
rect 37832 36110 37884 36116
rect 37648 35624 37700 35630
rect 37648 35566 37700 35572
rect 37556 34944 37608 34950
rect 37556 34886 37608 34892
rect 37568 34678 37596 34886
rect 37556 34672 37608 34678
rect 37556 34614 37608 34620
rect 37660 34610 37688 35566
rect 37740 35080 37792 35086
rect 37740 35022 37792 35028
rect 37648 34604 37700 34610
rect 37648 34546 37700 34552
rect 37464 33992 37516 33998
rect 37094 33960 37150 33969
rect 37464 33934 37516 33940
rect 37094 33895 37150 33904
rect 37476 33658 37504 33934
rect 37464 33652 37516 33658
rect 37464 33594 37516 33600
rect 37660 33454 37688 34546
rect 37752 34202 37780 35022
rect 37844 34746 37872 36110
rect 38028 36009 38056 37062
rect 38120 36242 38148 37295
rect 38108 36236 38160 36242
rect 38108 36178 38160 36184
rect 38014 36000 38070 36009
rect 38014 35935 38070 35944
rect 37924 35080 37976 35086
rect 37924 35022 37976 35028
rect 37832 34740 37884 34746
rect 37832 34682 37884 34688
rect 37936 34610 37964 35022
rect 38016 35012 38068 35018
rect 38016 34954 38068 34960
rect 38028 34678 38056 34954
rect 38016 34672 38068 34678
rect 38016 34614 38068 34620
rect 37924 34604 37976 34610
rect 37924 34546 37976 34552
rect 37740 34196 37792 34202
rect 37740 34138 37792 34144
rect 38028 34066 38056 34614
rect 38200 34604 38252 34610
rect 38200 34546 38252 34552
rect 38016 34060 38068 34066
rect 38016 34002 38068 34008
rect 38028 33522 38056 34002
rect 38212 33658 38240 34546
rect 38200 33652 38252 33658
rect 38200 33594 38252 33600
rect 38016 33516 38068 33522
rect 38016 33458 38068 33464
rect 37648 33448 37700 33454
rect 37648 33390 37700 33396
rect 37278 33280 37334 33289
rect 37278 33215 37334 33224
rect 37292 33114 37320 33215
rect 37280 33108 37332 33114
rect 37280 33050 37332 33056
rect 37660 32298 37688 33390
rect 37832 32904 37884 32910
rect 37832 32846 37884 32852
rect 38028 32858 38056 33458
rect 37844 32570 37872 32846
rect 38028 32830 38148 32858
rect 38016 32768 38068 32774
rect 38016 32710 38068 32716
rect 38028 32609 38056 32710
rect 38014 32600 38070 32609
rect 37832 32564 37884 32570
rect 38014 32535 38070 32544
rect 37832 32506 37884 32512
rect 37832 32428 37884 32434
rect 37832 32370 37884 32376
rect 37648 32292 37700 32298
rect 37648 32234 37700 32240
rect 37740 32020 37792 32026
rect 37740 31962 37792 31968
rect 36820 23316 36872 23322
rect 36820 23258 36872 23264
rect 36728 23112 36780 23118
rect 36728 23054 36780 23060
rect 36740 22778 36768 23054
rect 36728 22772 36780 22778
rect 36728 22714 36780 22720
rect 36636 22568 36688 22574
rect 36636 22510 36688 22516
rect 36544 3596 36596 3602
rect 36544 3538 36596 3544
rect 36648 3482 36676 22510
rect 37280 16448 37332 16454
rect 37280 16390 37332 16396
rect 37292 16182 37320 16390
rect 37280 16176 37332 16182
rect 37280 16118 37332 16124
rect 37280 15904 37332 15910
rect 37280 15846 37332 15852
rect 37292 15366 37320 15846
rect 37280 15360 37332 15366
rect 37280 15302 37332 15308
rect 37280 13184 37332 13190
rect 37280 13126 37332 13132
rect 37292 12646 37320 13126
rect 37280 12640 37332 12646
rect 37280 12582 37332 12588
rect 37280 10464 37332 10470
rect 37280 10406 37332 10412
rect 37292 10062 37320 10406
rect 37280 10056 37332 10062
rect 37280 9998 37332 10004
rect 37280 7744 37332 7750
rect 37280 7686 37332 7692
rect 37292 7342 37320 7686
rect 37280 7336 37332 7342
rect 37280 7278 37332 7284
rect 37188 6724 37240 6730
rect 37188 6666 37240 6672
rect 37200 6458 37228 6666
rect 37188 6452 37240 6458
rect 37188 6394 37240 6400
rect 37280 6248 37332 6254
rect 37280 6190 37332 6196
rect 37292 5914 37320 6190
rect 37280 5908 37332 5914
rect 37280 5850 37332 5856
rect 36728 4480 36780 4486
rect 36728 4422 36780 4428
rect 37648 4480 37700 4486
rect 37648 4422 37700 4428
rect 36556 3454 36676 3482
rect 36452 3188 36504 3194
rect 36452 3130 36504 3136
rect 36464 3058 36492 3130
rect 36452 3052 36504 3058
rect 36452 2994 36504 3000
rect 36556 2650 36584 3454
rect 36636 2848 36688 2854
rect 36636 2790 36688 2796
rect 36648 2689 36676 2790
rect 36634 2680 36690 2689
rect 36544 2644 36596 2650
rect 36634 2615 36690 2624
rect 36544 2586 36596 2592
rect 36740 2446 36768 4422
rect 37660 3058 37688 4422
rect 37752 3194 37780 31962
rect 37844 31958 37872 32370
rect 38016 32224 38068 32230
rect 38016 32166 38068 32172
rect 37832 31952 37884 31958
rect 38028 31929 38056 32166
rect 38120 32026 38148 32830
rect 38108 32020 38160 32026
rect 38108 31962 38160 31968
rect 37832 31894 37884 31900
rect 38014 31920 38070 31929
rect 38014 31855 38070 31864
rect 38014 31240 38070 31249
rect 38014 31175 38016 31184
rect 38068 31175 38070 31184
rect 38016 31146 38068 31152
rect 38016 30592 38068 30598
rect 38014 30560 38016 30569
rect 38068 30560 38070 30569
rect 38014 30495 38070 30504
rect 38016 30048 38068 30054
rect 38016 29990 38068 29996
rect 38028 29889 38056 29990
rect 38014 29880 38070 29889
rect 38014 29815 38070 29824
rect 38016 29504 38068 29510
rect 38016 29446 38068 29452
rect 38028 29209 38056 29446
rect 38014 29200 38070 29209
rect 38014 29135 38070 29144
rect 38014 28520 38070 28529
rect 38014 28455 38070 28464
rect 38028 28422 38056 28455
rect 38016 28416 38068 28422
rect 38016 28358 38068 28364
rect 37832 28076 37884 28082
rect 37832 28018 37884 28024
rect 37844 27606 37872 28018
rect 38016 27872 38068 27878
rect 38014 27840 38016 27849
rect 38068 27840 38070 27849
rect 38014 27775 38070 27784
rect 37832 27600 37884 27606
rect 37832 27542 37884 27548
rect 37832 27464 37884 27470
rect 37832 27406 37884 27412
rect 37844 27130 37872 27406
rect 38016 27328 38068 27334
rect 38016 27270 38068 27276
rect 38028 27169 38056 27270
rect 38014 27160 38070 27169
rect 37832 27124 37884 27130
rect 38014 27095 38070 27104
rect 37832 27066 37884 27072
rect 37832 26988 37884 26994
rect 37832 26930 37884 26936
rect 37844 26042 37872 26930
rect 38016 26784 38068 26790
rect 38016 26726 38068 26732
rect 38028 26489 38056 26726
rect 38014 26480 38070 26489
rect 38014 26415 38070 26424
rect 37832 26036 37884 26042
rect 37832 25978 37884 25984
rect 38014 25800 38070 25809
rect 38014 25735 38016 25744
rect 38068 25735 38070 25744
rect 38016 25706 38068 25712
rect 38016 25152 38068 25158
rect 38014 25120 38016 25129
rect 38068 25120 38070 25129
rect 38014 25055 38070 25064
rect 38016 24608 38068 24614
rect 38016 24550 38068 24556
rect 38028 24449 38056 24550
rect 38014 24440 38070 24449
rect 38014 24375 38070 24384
rect 37832 24200 37884 24206
rect 37832 24142 37884 24148
rect 37844 23526 37872 24142
rect 38016 24064 38068 24070
rect 38016 24006 38068 24012
rect 38028 23769 38056 24006
rect 38014 23760 38070 23769
rect 38014 23695 38070 23704
rect 37832 23520 37884 23526
rect 37832 23462 37884 23468
rect 38014 23080 38070 23089
rect 38014 23015 38070 23024
rect 38028 22982 38056 23015
rect 38016 22976 38068 22982
rect 38016 22918 38068 22924
rect 38016 22432 38068 22438
rect 38014 22400 38016 22409
rect 38068 22400 38070 22409
rect 38014 22335 38070 22344
rect 37832 22024 37884 22030
rect 37832 21966 37884 21972
rect 37844 21146 37872 21966
rect 38016 21888 38068 21894
rect 38016 21830 38068 21836
rect 38028 21729 38056 21830
rect 38014 21720 38070 21729
rect 38014 21655 38070 21664
rect 38108 21548 38160 21554
rect 38108 21490 38160 21496
rect 37924 21344 37976 21350
rect 37924 21286 37976 21292
rect 37832 21140 37884 21146
rect 37832 21082 37884 21088
rect 37936 20942 37964 21286
rect 38120 21049 38148 21490
rect 38106 21040 38162 21049
rect 38106 20975 38162 20984
rect 37924 20936 37976 20942
rect 37924 20878 37976 20884
rect 38014 20360 38070 20369
rect 38014 20295 38016 20304
rect 38068 20295 38070 20304
rect 38016 20266 38068 20272
rect 37832 19848 37884 19854
rect 37832 19790 37884 19796
rect 37844 19514 37872 19790
rect 38016 19712 38068 19718
rect 38014 19680 38016 19689
rect 38068 19680 38070 19689
rect 38014 19615 38070 19624
rect 37832 19508 37884 19514
rect 37832 19450 37884 19456
rect 38016 19168 38068 19174
rect 38016 19110 38068 19116
rect 38028 19009 38056 19110
rect 38014 19000 38070 19009
rect 38014 18935 38070 18944
rect 37832 18760 37884 18766
rect 37832 18702 37884 18708
rect 37844 18086 37872 18702
rect 38016 18624 38068 18630
rect 38016 18566 38068 18572
rect 38028 18329 38056 18566
rect 38014 18320 38070 18329
rect 38014 18255 38070 18264
rect 37832 18080 37884 18086
rect 37832 18022 37884 18028
rect 38014 17640 38070 17649
rect 38014 17575 38070 17584
rect 38028 17542 38056 17575
rect 38016 17536 38068 17542
rect 38016 17478 38068 17484
rect 38016 16992 38068 16998
rect 38014 16960 38016 16969
rect 38068 16960 38070 16969
rect 38014 16895 38070 16904
rect 38016 16448 38068 16454
rect 38016 16390 38068 16396
rect 38028 16289 38056 16390
rect 38014 16280 38070 16289
rect 38014 16215 38070 16224
rect 38016 15904 38068 15910
rect 38016 15846 38068 15852
rect 38028 15609 38056 15846
rect 38014 15600 38070 15609
rect 38014 15535 38070 15544
rect 38014 14920 38070 14929
rect 38014 14855 38016 14864
rect 38068 14855 38070 14864
rect 38016 14826 38068 14832
rect 38016 14272 38068 14278
rect 38014 14240 38016 14249
rect 38068 14240 38070 14249
rect 38014 14175 38070 14184
rect 38016 13728 38068 13734
rect 38016 13670 38068 13676
rect 38028 13569 38056 13670
rect 38014 13560 38070 13569
rect 38014 13495 38070 13504
rect 38016 13184 38068 13190
rect 38016 13126 38068 13132
rect 38028 12889 38056 13126
rect 38014 12880 38070 12889
rect 38014 12815 38070 12824
rect 38014 12200 38070 12209
rect 38014 12135 38070 12144
rect 38028 12102 38056 12135
rect 38016 12096 38068 12102
rect 38016 12038 38068 12044
rect 38016 11552 38068 11558
rect 38014 11520 38016 11529
rect 38068 11520 38070 11529
rect 38014 11455 38070 11464
rect 38016 11280 38068 11286
rect 38016 11222 38068 11228
rect 38028 10849 38056 11222
rect 38014 10840 38070 10849
rect 38014 10775 38070 10784
rect 37924 10736 37976 10742
rect 37924 10678 37976 10684
rect 37936 4146 37964 10678
rect 38016 10464 38068 10470
rect 38016 10406 38068 10412
rect 38028 10169 38056 10406
rect 38014 10160 38070 10169
rect 38014 10095 38070 10104
rect 38014 9480 38070 9489
rect 38014 9415 38016 9424
rect 38068 9415 38070 9424
rect 38016 9386 38068 9392
rect 38016 8832 38068 8838
rect 38014 8800 38016 8809
rect 38068 8800 38070 8809
rect 38014 8735 38070 8744
rect 38016 8356 38068 8362
rect 38016 8298 38068 8304
rect 38028 8129 38056 8298
rect 38014 8120 38070 8129
rect 38014 8055 38070 8064
rect 38016 7744 38068 7750
rect 38016 7686 38068 7692
rect 38028 7449 38056 7686
rect 38014 7440 38070 7449
rect 38014 7375 38070 7384
rect 38014 6760 38070 6769
rect 38014 6695 38070 6704
rect 38028 6662 38056 6695
rect 38016 6656 38068 6662
rect 38016 6598 38068 6604
rect 38016 6112 38068 6118
rect 38014 6080 38016 6089
rect 38068 6080 38070 6089
rect 38014 6015 38070 6024
rect 38016 5568 38068 5574
rect 38016 5510 38068 5516
rect 38028 5409 38056 5510
rect 38014 5400 38070 5409
rect 38014 5335 38070 5344
rect 38016 5024 38068 5030
rect 38016 4966 38068 4972
rect 38028 4729 38056 4966
rect 38014 4720 38070 4729
rect 38014 4655 38070 4664
rect 38016 4480 38068 4486
rect 38016 4422 38068 4428
rect 38028 4214 38056 4422
rect 38016 4208 38068 4214
rect 38016 4150 38068 4156
rect 37924 4140 37976 4146
rect 37924 4082 37976 4088
rect 38028 4049 38056 4150
rect 38014 4040 38070 4049
rect 37832 4004 37884 4010
rect 38014 3975 38070 3984
rect 37832 3946 37884 3952
rect 37844 3534 37872 3946
rect 37832 3528 37884 3534
rect 37832 3470 37884 3476
rect 38016 3392 38068 3398
rect 38014 3360 38016 3369
rect 38068 3360 38070 3369
rect 38014 3295 38070 3304
rect 37740 3188 37792 3194
rect 37740 3130 37792 3136
rect 37648 3052 37700 3058
rect 37648 2994 37700 3000
rect 36728 2440 36780 2446
rect 36780 2388 36952 2394
rect 36728 2382 36952 2388
rect 36740 2366 36952 2382
rect 36924 800 36952 2366
rect 37660 800 37688 2994
rect 2318 0 2374 800
rect 3054 0 3110 800
rect 3790 0 3846 800
rect 4526 0 4582 800
rect 5262 0 5318 800
rect 5998 0 6054 800
rect 6734 0 6790 800
rect 7470 0 7526 800
rect 8206 0 8262 800
rect 8942 0 8998 800
rect 9678 0 9734 800
rect 10414 0 10470 800
rect 11150 0 11206 800
rect 11886 0 11942 800
rect 12622 0 12678 800
rect 13358 0 13414 800
rect 14094 0 14150 800
rect 14830 0 14886 800
rect 15566 0 15622 800
rect 16302 0 16358 800
rect 17038 0 17094 800
rect 17774 0 17830 800
rect 18510 0 18566 800
rect 19246 0 19302 800
rect 19982 0 20038 800
rect 20718 0 20774 800
rect 21454 0 21510 800
rect 22190 0 22246 800
rect 22926 0 22982 800
rect 23662 0 23718 800
rect 24398 0 24454 800
rect 25134 0 25190 800
rect 25870 0 25926 800
rect 26606 0 26662 800
rect 27342 0 27398 800
rect 28078 0 28134 800
rect 28814 0 28870 800
rect 29550 0 29606 800
rect 30286 0 30342 800
rect 31022 0 31078 800
rect 31758 0 31814 800
rect 32494 0 32550 800
rect 33230 0 33286 800
rect 33966 0 34022 800
rect 34702 0 34758 800
rect 35438 0 35494 800
rect 36174 0 36230 800
rect 36910 0 36966 800
rect 37646 0 37702 800
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 36174 36624 36230 36680
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 38106 37304 38162 37360
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 37002 34584 37058 34640
rect 37186 35264 37242 35320
rect 37094 33904 37150 33960
rect 38014 35944 38070 36000
rect 37278 33224 37334 33280
rect 38014 32544 38070 32600
rect 36634 2624 36690 2680
rect 38014 31864 38070 31920
rect 38014 31204 38070 31240
rect 38014 31184 38016 31204
rect 38016 31184 38068 31204
rect 38068 31184 38070 31204
rect 38014 30540 38016 30560
rect 38016 30540 38068 30560
rect 38068 30540 38070 30560
rect 38014 30504 38070 30540
rect 38014 29824 38070 29880
rect 38014 29144 38070 29200
rect 38014 28464 38070 28520
rect 38014 27820 38016 27840
rect 38016 27820 38068 27840
rect 38068 27820 38070 27840
rect 38014 27784 38070 27820
rect 38014 27104 38070 27160
rect 38014 26424 38070 26480
rect 38014 25764 38070 25800
rect 38014 25744 38016 25764
rect 38016 25744 38068 25764
rect 38068 25744 38070 25764
rect 38014 25100 38016 25120
rect 38016 25100 38068 25120
rect 38068 25100 38070 25120
rect 38014 25064 38070 25100
rect 38014 24384 38070 24440
rect 38014 23704 38070 23760
rect 38014 23024 38070 23080
rect 38014 22380 38016 22400
rect 38016 22380 38068 22400
rect 38068 22380 38070 22400
rect 38014 22344 38070 22380
rect 38014 21664 38070 21720
rect 38106 20984 38162 21040
rect 38014 20324 38070 20360
rect 38014 20304 38016 20324
rect 38016 20304 38068 20324
rect 38068 20304 38070 20324
rect 38014 19660 38016 19680
rect 38016 19660 38068 19680
rect 38068 19660 38070 19680
rect 38014 19624 38070 19660
rect 38014 18944 38070 19000
rect 38014 18264 38070 18320
rect 38014 17584 38070 17640
rect 38014 16940 38016 16960
rect 38016 16940 38068 16960
rect 38068 16940 38070 16960
rect 38014 16904 38070 16940
rect 38014 16224 38070 16280
rect 38014 15544 38070 15600
rect 38014 14884 38070 14920
rect 38014 14864 38016 14884
rect 38016 14864 38068 14884
rect 38068 14864 38070 14884
rect 38014 14220 38016 14240
rect 38016 14220 38068 14240
rect 38068 14220 38070 14240
rect 38014 14184 38070 14220
rect 38014 13504 38070 13560
rect 38014 12824 38070 12880
rect 38014 12144 38070 12200
rect 38014 11500 38016 11520
rect 38016 11500 38068 11520
rect 38068 11500 38070 11520
rect 38014 11464 38070 11500
rect 38014 10784 38070 10840
rect 38014 10104 38070 10160
rect 38014 9444 38070 9480
rect 38014 9424 38016 9444
rect 38016 9424 38068 9444
rect 38068 9424 38070 9444
rect 38014 8780 38016 8800
rect 38016 8780 38068 8800
rect 38068 8780 38070 8800
rect 38014 8744 38070 8780
rect 38014 8064 38070 8120
rect 38014 7384 38070 7440
rect 38014 6704 38070 6760
rect 38014 6060 38016 6080
rect 38016 6060 38068 6080
rect 38068 6060 38070 6080
rect 38014 6024 38070 6060
rect 38014 5344 38070 5400
rect 38014 4664 38070 4720
rect 38014 3984 38070 4040
rect 38014 3340 38016 3360
rect 38016 3340 38068 3360
rect 38068 3340 38070 3360
rect 38014 3304 38070 3340
<< metal3 >>
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 38101 37362 38167 37365
rect 39200 37362 40000 37392
rect 38101 37360 40000 37362
rect 38101 37304 38106 37360
rect 38162 37304 40000 37360
rect 38101 37302 40000 37304
rect 38101 37299 38167 37302
rect 39200 37272 40000 37302
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 36169 36682 36235 36685
rect 39200 36682 40000 36712
rect 36169 36680 40000 36682
rect 36169 36624 36174 36680
rect 36230 36624 40000 36680
rect 36169 36622 40000 36624
rect 36169 36619 36235 36622
rect 39200 36592 40000 36622
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 38009 36002 38075 36005
rect 39200 36002 40000 36032
rect 38009 36000 40000 36002
rect 38009 35944 38014 36000
rect 38070 35944 40000 36000
rect 38009 35942 40000 35944
rect 38009 35939 38075 35942
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 39200 35912 40000 35942
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 37181 35322 37247 35325
rect 39200 35322 40000 35352
rect 37181 35320 40000 35322
rect 37181 35264 37186 35320
rect 37242 35264 40000 35320
rect 37181 35262 40000 35264
rect 37181 35259 37247 35262
rect 39200 35232 40000 35262
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 36997 34642 37063 34645
rect 39200 34642 40000 34672
rect 36997 34640 40000 34642
rect 36997 34584 37002 34640
rect 37058 34584 40000 34640
rect 36997 34582 40000 34584
rect 36997 34579 37063 34582
rect 39200 34552 40000 34582
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 37089 33962 37155 33965
rect 39200 33962 40000 33992
rect 37089 33960 40000 33962
rect 37089 33904 37094 33960
rect 37150 33904 40000 33960
rect 37089 33902 40000 33904
rect 37089 33899 37155 33902
rect 39200 33872 40000 33902
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 37273 33282 37339 33285
rect 39200 33282 40000 33312
rect 37273 33280 40000 33282
rect 37273 33224 37278 33280
rect 37334 33224 40000 33280
rect 37273 33222 40000 33224
rect 37273 33219 37339 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 39200 33192 40000 33222
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 38009 32602 38075 32605
rect 39200 32602 40000 32632
rect 38009 32600 40000 32602
rect 38009 32544 38014 32600
rect 38070 32544 40000 32600
rect 38009 32542 40000 32544
rect 38009 32539 38075 32542
rect 39200 32512 40000 32542
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 38009 31922 38075 31925
rect 39200 31922 40000 31952
rect 38009 31920 40000 31922
rect 38009 31864 38014 31920
rect 38070 31864 40000 31920
rect 38009 31862 40000 31864
rect 38009 31859 38075 31862
rect 39200 31832 40000 31862
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 38009 31242 38075 31245
rect 39200 31242 40000 31272
rect 38009 31240 40000 31242
rect 38009 31184 38014 31240
rect 38070 31184 40000 31240
rect 38009 31182 40000 31184
rect 38009 31179 38075 31182
rect 39200 31152 40000 31182
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 38009 30562 38075 30565
rect 39200 30562 40000 30592
rect 38009 30560 40000 30562
rect 38009 30504 38014 30560
rect 38070 30504 40000 30560
rect 38009 30502 40000 30504
rect 38009 30499 38075 30502
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 39200 30472 40000 30502
rect 19570 30431 19886 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 38009 29882 38075 29885
rect 39200 29882 40000 29912
rect 38009 29880 40000 29882
rect 38009 29824 38014 29880
rect 38070 29824 40000 29880
rect 38009 29822 40000 29824
rect 38009 29819 38075 29822
rect 39200 29792 40000 29822
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 38009 29202 38075 29205
rect 39200 29202 40000 29232
rect 38009 29200 40000 29202
rect 38009 29144 38014 29200
rect 38070 29144 40000 29200
rect 38009 29142 40000 29144
rect 38009 29139 38075 29142
rect 39200 29112 40000 29142
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 38009 28522 38075 28525
rect 39200 28522 40000 28552
rect 38009 28520 40000 28522
rect 38009 28464 38014 28520
rect 38070 28464 40000 28520
rect 38009 28462 40000 28464
rect 38009 28459 38075 28462
rect 39200 28432 40000 28462
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 38009 27842 38075 27845
rect 39200 27842 40000 27872
rect 38009 27840 40000 27842
rect 38009 27784 38014 27840
rect 38070 27784 40000 27840
rect 38009 27782 40000 27784
rect 38009 27779 38075 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 39200 27752 40000 27782
rect 34930 27711 35246 27712
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 38009 27162 38075 27165
rect 39200 27162 40000 27192
rect 38009 27160 40000 27162
rect 38009 27104 38014 27160
rect 38070 27104 40000 27160
rect 38009 27102 40000 27104
rect 38009 27099 38075 27102
rect 39200 27072 40000 27102
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 38009 26482 38075 26485
rect 39200 26482 40000 26512
rect 38009 26480 40000 26482
rect 38009 26424 38014 26480
rect 38070 26424 40000 26480
rect 38009 26422 40000 26424
rect 38009 26419 38075 26422
rect 39200 26392 40000 26422
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 38009 25802 38075 25805
rect 39200 25802 40000 25832
rect 38009 25800 40000 25802
rect 38009 25744 38014 25800
rect 38070 25744 40000 25800
rect 38009 25742 40000 25744
rect 38009 25739 38075 25742
rect 39200 25712 40000 25742
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 38009 25122 38075 25125
rect 39200 25122 40000 25152
rect 38009 25120 40000 25122
rect 38009 25064 38014 25120
rect 38070 25064 40000 25120
rect 38009 25062 40000 25064
rect 38009 25059 38075 25062
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 39200 25032 40000 25062
rect 19570 24991 19886 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 38009 24442 38075 24445
rect 39200 24442 40000 24472
rect 38009 24440 40000 24442
rect 38009 24384 38014 24440
rect 38070 24384 40000 24440
rect 38009 24382 40000 24384
rect 38009 24379 38075 24382
rect 39200 24352 40000 24382
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 38009 23762 38075 23765
rect 39200 23762 40000 23792
rect 38009 23760 40000 23762
rect 38009 23704 38014 23760
rect 38070 23704 40000 23760
rect 38009 23702 40000 23704
rect 38009 23699 38075 23702
rect 39200 23672 40000 23702
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 38009 23082 38075 23085
rect 39200 23082 40000 23112
rect 38009 23080 40000 23082
rect 38009 23024 38014 23080
rect 38070 23024 40000 23080
rect 38009 23022 40000 23024
rect 38009 23019 38075 23022
rect 39200 22992 40000 23022
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 38009 22402 38075 22405
rect 39200 22402 40000 22432
rect 38009 22400 40000 22402
rect 38009 22344 38014 22400
rect 38070 22344 40000 22400
rect 38009 22342 40000 22344
rect 38009 22339 38075 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 39200 22312 40000 22342
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 38009 21722 38075 21725
rect 39200 21722 40000 21752
rect 38009 21720 40000 21722
rect 38009 21664 38014 21720
rect 38070 21664 40000 21720
rect 38009 21662 40000 21664
rect 38009 21659 38075 21662
rect 39200 21632 40000 21662
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 38101 21042 38167 21045
rect 39200 21042 40000 21072
rect 38101 21040 40000 21042
rect 38101 20984 38106 21040
rect 38162 20984 40000 21040
rect 38101 20982 40000 20984
rect 38101 20979 38167 20982
rect 39200 20952 40000 20982
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 38009 20362 38075 20365
rect 39200 20362 40000 20392
rect 38009 20360 40000 20362
rect 38009 20304 38014 20360
rect 38070 20304 40000 20360
rect 38009 20302 40000 20304
rect 38009 20299 38075 20302
rect 39200 20272 40000 20302
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 38009 19682 38075 19685
rect 39200 19682 40000 19712
rect 38009 19680 40000 19682
rect 38009 19624 38014 19680
rect 38070 19624 40000 19680
rect 38009 19622 40000 19624
rect 38009 19619 38075 19622
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 39200 19592 40000 19622
rect 19570 19551 19886 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 38009 19002 38075 19005
rect 39200 19002 40000 19032
rect 38009 19000 40000 19002
rect 38009 18944 38014 19000
rect 38070 18944 40000 19000
rect 38009 18942 40000 18944
rect 38009 18939 38075 18942
rect 39200 18912 40000 18942
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 38009 18322 38075 18325
rect 39200 18322 40000 18352
rect 38009 18320 40000 18322
rect 38009 18264 38014 18320
rect 38070 18264 40000 18320
rect 38009 18262 40000 18264
rect 38009 18259 38075 18262
rect 39200 18232 40000 18262
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 38009 17642 38075 17645
rect 39200 17642 40000 17672
rect 38009 17640 40000 17642
rect 38009 17584 38014 17640
rect 38070 17584 40000 17640
rect 38009 17582 40000 17584
rect 38009 17579 38075 17582
rect 39200 17552 40000 17582
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 38009 16962 38075 16965
rect 39200 16962 40000 16992
rect 38009 16960 40000 16962
rect 38009 16904 38014 16960
rect 38070 16904 40000 16960
rect 38009 16902 40000 16904
rect 38009 16899 38075 16902
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 39200 16872 40000 16902
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 38009 16282 38075 16285
rect 39200 16282 40000 16312
rect 38009 16280 40000 16282
rect 38009 16224 38014 16280
rect 38070 16224 40000 16280
rect 38009 16222 40000 16224
rect 38009 16219 38075 16222
rect 39200 16192 40000 16222
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 38009 15602 38075 15605
rect 39200 15602 40000 15632
rect 38009 15600 40000 15602
rect 38009 15544 38014 15600
rect 38070 15544 40000 15600
rect 38009 15542 40000 15544
rect 38009 15539 38075 15542
rect 39200 15512 40000 15542
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 38009 14922 38075 14925
rect 39200 14922 40000 14952
rect 38009 14920 40000 14922
rect 38009 14864 38014 14920
rect 38070 14864 40000 14920
rect 38009 14862 40000 14864
rect 38009 14859 38075 14862
rect 39200 14832 40000 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 38009 14242 38075 14245
rect 39200 14242 40000 14272
rect 38009 14240 40000 14242
rect 38009 14184 38014 14240
rect 38070 14184 40000 14240
rect 38009 14182 40000 14184
rect 38009 14179 38075 14182
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 39200 14152 40000 14182
rect 19570 14111 19886 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 38009 13562 38075 13565
rect 39200 13562 40000 13592
rect 38009 13560 40000 13562
rect 38009 13504 38014 13560
rect 38070 13504 40000 13560
rect 38009 13502 40000 13504
rect 38009 13499 38075 13502
rect 39200 13472 40000 13502
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 38009 12882 38075 12885
rect 39200 12882 40000 12912
rect 38009 12880 40000 12882
rect 38009 12824 38014 12880
rect 38070 12824 40000 12880
rect 38009 12822 40000 12824
rect 38009 12819 38075 12822
rect 39200 12792 40000 12822
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 38009 12202 38075 12205
rect 39200 12202 40000 12232
rect 38009 12200 40000 12202
rect 38009 12144 38014 12200
rect 38070 12144 40000 12200
rect 38009 12142 40000 12144
rect 38009 12139 38075 12142
rect 39200 12112 40000 12142
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 38009 11522 38075 11525
rect 39200 11522 40000 11552
rect 38009 11520 40000 11522
rect 38009 11464 38014 11520
rect 38070 11464 40000 11520
rect 38009 11462 40000 11464
rect 38009 11459 38075 11462
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 39200 11432 40000 11462
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 38009 10842 38075 10845
rect 39200 10842 40000 10872
rect 38009 10840 40000 10842
rect 38009 10784 38014 10840
rect 38070 10784 40000 10840
rect 38009 10782 40000 10784
rect 38009 10779 38075 10782
rect 39200 10752 40000 10782
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 38009 10162 38075 10165
rect 39200 10162 40000 10192
rect 38009 10160 40000 10162
rect 38009 10104 38014 10160
rect 38070 10104 40000 10160
rect 38009 10102 40000 10104
rect 38009 10099 38075 10102
rect 39200 10072 40000 10102
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 38009 9482 38075 9485
rect 39200 9482 40000 9512
rect 38009 9480 40000 9482
rect 38009 9424 38014 9480
rect 38070 9424 40000 9480
rect 38009 9422 40000 9424
rect 38009 9419 38075 9422
rect 39200 9392 40000 9422
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 38009 8802 38075 8805
rect 39200 8802 40000 8832
rect 38009 8800 40000 8802
rect 38009 8744 38014 8800
rect 38070 8744 40000 8800
rect 38009 8742 40000 8744
rect 38009 8739 38075 8742
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 39200 8712 40000 8742
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 38009 8122 38075 8125
rect 39200 8122 40000 8152
rect 38009 8120 40000 8122
rect 38009 8064 38014 8120
rect 38070 8064 40000 8120
rect 38009 8062 40000 8064
rect 38009 8059 38075 8062
rect 39200 8032 40000 8062
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 38009 7442 38075 7445
rect 39200 7442 40000 7472
rect 38009 7440 40000 7442
rect 38009 7384 38014 7440
rect 38070 7384 40000 7440
rect 38009 7382 40000 7384
rect 38009 7379 38075 7382
rect 39200 7352 40000 7382
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 38009 6762 38075 6765
rect 39200 6762 40000 6792
rect 38009 6760 40000 6762
rect 38009 6704 38014 6760
rect 38070 6704 40000 6760
rect 38009 6702 40000 6704
rect 38009 6699 38075 6702
rect 39200 6672 40000 6702
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 38009 6082 38075 6085
rect 39200 6082 40000 6112
rect 38009 6080 40000 6082
rect 38009 6024 38014 6080
rect 38070 6024 40000 6080
rect 38009 6022 40000 6024
rect 38009 6019 38075 6022
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 39200 5992 40000 6022
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 38009 5402 38075 5405
rect 39200 5402 40000 5432
rect 38009 5400 40000 5402
rect 38009 5344 38014 5400
rect 38070 5344 40000 5400
rect 38009 5342 40000 5344
rect 38009 5339 38075 5342
rect 39200 5312 40000 5342
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 38009 4722 38075 4725
rect 39200 4722 40000 4752
rect 38009 4720 40000 4722
rect 38009 4664 38014 4720
rect 38070 4664 40000 4720
rect 38009 4662 40000 4664
rect 38009 4659 38075 4662
rect 39200 4632 40000 4662
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 38009 4042 38075 4045
rect 39200 4042 40000 4072
rect 38009 4040 40000 4042
rect 38009 3984 38014 4040
rect 38070 3984 40000 4040
rect 38009 3982 40000 3984
rect 38009 3979 38075 3982
rect 39200 3952 40000 3982
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 38009 3362 38075 3365
rect 39200 3362 40000 3392
rect 38009 3360 40000 3362
rect 38009 3304 38014 3360
rect 38070 3304 40000 3360
rect 38009 3302 40000 3304
rect 38009 3299 38075 3302
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 39200 3272 40000 3302
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 36629 2682 36695 2685
rect 39200 2682 40000 2712
rect 36629 2680 40000 2682
rect 36629 2624 36634 2680
rect 36690 2624 40000 2680
rect 36629 2622 40000 2624
rect 36629 2619 36695 2622
rect 39200 2592 40000 2622
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__060__A opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 28612 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__A0
timestamp 1649977179
transform -1 0 12144 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__061__S
timestamp 1649977179
transform -1 0 14260 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__A0
timestamp 1649977179
transform 1 0 11316 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__063__S
timestamp 1649977179
transform -1 0 11040 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__065__A_N
timestamp 1649977179
transform 1 0 23644 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__A_N
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__067__B
timestamp 1649977179
transform 1 0 12972 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__A1
timestamp 1649977179
transform -1 0 35512 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__069__S
timestamp 1649977179
transform 1 0 33856 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__A1
timestamp 1649977179
transform -1 0 36156 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__071__S
timestamp 1649977179
transform 1 0 34960 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__073__A
timestamp 1649977179
transform 1 0 20884 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__A1
timestamp 1649977179
transform -1 0 37444 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__074__S
timestamp 1649977179
transform -1 0 35604 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__A0
timestamp 1649977179
transform -1 0 7176 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__076__S
timestamp 1649977179
transform 1 0 9292 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__A0
timestamp 1649977179
transform 1 0 6532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__078__S
timestamp 1649977179
transform -1 0 7268 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__A0
timestamp 1649977179
transform 1 0 6992 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__080__S
timestamp 1649977179
transform 1 0 8740 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__A0
timestamp 1649977179
transform -1 0 7268 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__082__S
timestamp 1649977179
transform 1 0 10120 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__A0
timestamp 1649977179
transform -1 0 10580 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__084__S
timestamp 1649977179
transform 1 0 7268 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__A0
timestamp 1649977179
transform -1 0 9108 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__086__S
timestamp 1649977179
transform 1 0 8280 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__A0
timestamp 1649977179
transform -1 0 10212 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__088__S
timestamp 1649977179
transform 1 0 10580 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__A0
timestamp 1649977179
transform -1 0 9660 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__090__S
timestamp 1649977179
transform 1 0 9752 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__A0
timestamp 1649977179
transform -1 0 10488 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__092__S
timestamp 1649977179
transform 1 0 9476 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__094__A
timestamp 1649977179
transform 1 0 19780 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__095__A0
timestamp 1649977179
transform 1 0 11868 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__097__A0
timestamp 1649977179
transform -1 0 12236 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__099__A0
timestamp 1649977179
transform -1 0 14904 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__101__A0
timestamp 1649977179
transform -1 0 15180 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__103__A0
timestamp 1649977179
transform -1 0 15088 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__105__A0
timestamp 1649977179
transform -1 0 15640 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__107__A0
timestamp 1649977179
transform -1 0 16652 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__109__A0
timestamp 1649977179
transform -1 0 17480 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__111__A0
timestamp 1649977179
transform -1 0 18032 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__113__A0
timestamp 1649977179
transform -1 0 19412 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1649977179
transform 1 0 23460 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__116__A0
timestamp 1649977179
transform -1 0 18768 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__A0
timestamp 1649977179
transform -1 0 20148 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__120__A0
timestamp 1649977179
transform -1 0 20700 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__A1
timestamp 1649977179
transform -1 0 23644 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__128__A1
timestamp 1649977179
transform -1 0 24564 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__130__A1
timestamp 1649977179
transform -1 0 25392 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__A1
timestamp 1649977179
transform -1 0 26404 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A1
timestamp 1649977179
transform -1 0 26404 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__136__A
timestamp 1649977179
transform 1 0 31372 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__A1
timestamp 1649977179
transform -1 0 29624 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A1
timestamp 1649977179
transform -1 0 28152 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__141__A1
timestamp 1649977179
transform -1 0 29716 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A1
timestamp 1649977179
transform -1 0 30544 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A1
timestamp 1649977179
transform -1 0 30728 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A1
timestamp 1649977179
transform -1 0 32016 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__A1
timestamp 1649977179
transform -1 0 32568 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__151__A1
timestamp 1649977179
transform -1 0 34132 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__A1
timestamp 1649977179
transform -1 0 33212 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__155__A1
timestamp 1649977179
transform 1 0 33580 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A1
timestamp 1649977179
transform 1 0 34224 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__S
timestamp 1649977179
transform 1 0 34776 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A1
timestamp 1649977179
transform -1 0 35512 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__S
timestamp 1649977179
transform 1 0 36248 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__A1
timestamp 1649977179
transform -1 0 35512 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__S
timestamp 1649977179
transform 1 0 37260 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__165__A
timestamp 1649977179
transform 1 0 23644 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__A
timestamp 1649977179
transform 1 0 14720 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__167__B
timestamp 1649977179
transform 1 0 14168 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__A1
timestamp 1649977179
transform 1 0 37260 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__169__A2
timestamp 1649977179
transform -1 0 38180 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A1
timestamp 1649977179
transform -1 0 36800 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__A2
timestamp 1649977179
transform -1 0 35880 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__171__CLK
timestamp 1649977179
transform -1 0 34868 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 36248 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 35420 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 37628 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 38180 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 37536 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 2024 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 2760 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1649977179
transform -1 0 4600 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1649977179
transform -1 0 12052 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1649977179
transform -1 0 12788 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1649977179
transform -1 0 14260 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1649977179
transform -1 0 13800 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1649977179
transform -1 0 15088 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1649977179
transform -1 0 15640 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1649977179
transform -1 0 16192 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1649977179
transform -1 0 17112 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1649977179
transform -1 0 17848 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1649977179
transform -1 0 18768 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1649977179
transform -1 0 6532 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1649977179
transform -1 0 19320 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1649977179
transform -1 0 20056 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1649977179
transform -1 0 20792 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1649977179
transform -1 0 22632 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1649977179
transform -1 0 5704 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1649977179
transform -1 0 7544 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1649977179
transform -1 0 7176 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1649977179
transform -1 0 8280 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1649977179
transform -1 0 9016 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1649977179
transform -1 0 10488 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1649977179
transform -1 0 9752 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1649977179
transform -1 0 11500 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1649977179
transform -1 0 23828 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1649977179
transform -1 0 31648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1649977179
transform -1 0 30728 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1649977179
transform -1 0 32292 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1649977179
transform -1 0 32844 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1649977179
transform -1 0 34224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1649977179
transform -1 0 34592 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1649977179
transform -1 0 24380 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1649977179
transform -1 0 25024 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1649977179
transform -1 0 26496 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1649977179
transform -1 0 25576 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1649977179
transform -1 0 27140 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1649977179
transform -1 0 27692 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1649977179
transform -1 0 29072 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1649977179
transform -1 0 29532 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1649977179
transform -1 0 30176 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1649977179
transform -1 0 36800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1649977179
transform -1 0 35696 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1649977179
transform -1 0 37444 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1649977179
transform -1 0 37444 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1649977179
transform -1 0 2024 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1649977179
transform -1 0 3496 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1649977179
transform -1 0 4232 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1649977179
transform -1 0 11960 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1649977179
transform -1 0 12696 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1649977179
transform -1 0 14260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1649977179
transform -1 0 13800 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1649977179
transform -1 0 15088 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1649977179
transform -1 0 15640 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1649977179
transform -1 0 16192 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1649977179
transform -1 0 17112 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1649977179
transform -1 0 17848 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1649977179
transform -1 0 18768 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input65_A
timestamp 1649977179
transform -1 0 5428 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input66_A
timestamp 1649977179
transform -1 0 19320 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input67_A
timestamp 1649977179
transform -1 0 20056 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input68_A
timestamp 1649977179
transform -1 0 20792 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input69_A
timestamp 1649977179
transform -1 0 22632 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input70_A
timestamp 1649977179
transform -1 0 5888 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input71_A
timestamp 1649977179
transform -1 0 6808 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input72_A
timestamp 1649977179
transform -1 0 7544 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input73_A
timestamp 1649977179
transform -1 0 9108 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input74_A
timestamp 1649977179
transform -1 0 8648 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input75_A
timestamp 1649977179
transform -1 0 9936 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input76_A
timestamp 1649977179
transform -1 0 10488 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input77_A
timestamp 1649977179
transform -1 0 11040 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input78_A
timestamp 1649977179
transform -1 0 23828 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input79_A
timestamp 1649977179
transform -1 0 30360 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input80_A
timestamp 1649977179
transform -1 0 31648 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input81_A
timestamp 1649977179
transform -1 0 32108 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input82_A
timestamp 1649977179
transform -1 0 33396 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input83_A
timestamp 1649977179
transform -1 0 36156 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input84_A
timestamp 1649977179
transform 1 0 34040 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input85_A
timestamp 1649977179
transform -1 0 24380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input86_A
timestamp 1649977179
transform -1 0 25024 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input87_A
timestamp 1649977179
transform -1 0 26496 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input88_A
timestamp 1649977179
transform -1 0 25576 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input89_A
timestamp 1649977179
transform -1 0 27140 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input90_A
timestamp 1649977179
transform -1 0 27692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input91_A
timestamp 1649977179
transform -1 0 29072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input92_A
timestamp 1649977179
transform -1 0 29716 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input93_A
timestamp 1649977179
transform -1 0 31096 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input94_A
timestamp 1649977179
transform -1 0 34776 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input95_A
timestamp 1649977179
transform -1 0 33672 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input96_A
timestamp 1649977179
transform -1 0 36248 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input97_A
timestamp 1649977179
transform -1 0 36984 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output98_A
timestamp 1649977179
transform 1 0 34960 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output100_A
timestamp 1649977179
transform -1 0 36800 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output101_A
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output102_A
timestamp 1649977179
transform -1 0 37444 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output103_A
timestamp 1649977179
transform -1 0 37444 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output104_A
timestamp 1649977179
transform -1 0 37444 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output105_A
timestamp 1649977179
transform -1 0 37444 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output106_A
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output107_A
timestamp 1649977179
transform -1 0 37444 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output108_A
timestamp 1649977179
transform -1 0 37444 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output109_A
timestamp 1649977179
transform 1 0 37260 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output110_A
timestamp 1649977179
transform -1 0 37444 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output111_A
timestamp 1649977179
transform -1 0 37444 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output112_A
timestamp 1649977179
transform -1 0 37444 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output113_A
timestamp 1649977179
transform 1 0 37260 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output118_A
timestamp 1649977179
transform -1 0 37444 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output119_A
timestamp 1649977179
transform -1 0 37444 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output120_A
timestamp 1649977179
transform -1 0 37444 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output121_A
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output122_A
timestamp 1649977179
transform -1 0 37444 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output123_A
timestamp 1649977179
transform -1 0 37444 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output124_A
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output125_A
timestamp 1649977179
transform -1 0 37444 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output146_A
timestamp 1649977179
transform 1 0 4968 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output149_A
timestamp 1649977179
transform -1 0 23184 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1748 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10
timestamp 1649977179
transform 1 0 2024 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17
timestamp 1649977179
transform 1 0 2668 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24
timestamp 1649977179
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 4232 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45
timestamp 1649977179
transform 1 0 5244 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52
timestamp 1649977179
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61
timestamp 1649977179
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65
timestamp 1649977179
transform 1 0 7084 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_73
timestamp 1649977179
transform 1 0 7820 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1649977179
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_87
timestamp 1649977179
transform 1 0 9108 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_94
timestamp 1649977179
transform 1 0 9752 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_101
timestamp 1649977179
transform 1 0 10396 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_108
timestamp 1649977179
transform 1 0 11040 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_117
timestamp 1649977179
transform 1 0 11868 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_121
timestamp 1649977179
transform 1 0 12236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_129
timestamp 1649977179
transform 1 0 12972 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_136
timestamp 1649977179
transform 1 0 13616 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_143
timestamp 1649977179
transform 1 0 14260 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_150
timestamp 1649977179
transform 1 0 14904 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_157
timestamp 1649977179
transform 1 0 15548 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1649977179
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_169
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_173
timestamp 1649977179
transform 1 0 17020 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_177
timestamp 1649977179
transform 1 0 17388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_181
timestamp 1649977179
transform 1 0 17756 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_185
timestamp 1649977179
transform 1 0 18124 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1649977179
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_201
timestamp 1649977179
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1649977179
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_213
timestamp 1649977179
transform 1 0 20700 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_217 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_223
timestamp 1649977179
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_229
timestamp 1649977179
transform 1 0 22172 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_234
timestamp 1649977179
transform 1 0 22632 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_241
timestamp 1649977179
transform 1 0 23276 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1649977179
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1649977179
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_256
timestamp 1649977179
transform 1 0 24656 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_263
timestamp 1649977179
transform 1 0 25300 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_270
timestamp 1649977179
transform 1 0 25944 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1649977179
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_284
timestamp 1649977179
transform 1 0 27232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_291
timestamp 1649977179
transform 1 0 27876 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_298
timestamp 1649977179
transform 1 0 28520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1649977179
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_320
timestamp 1649977179
transform 1 0 30544 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_326
timestamp 1649977179
transform 1 0 31096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1649977179
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_347
timestamp 1649977179
transform 1 0 33028 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_351
timestamp 1649977179
transform 1 0 33396 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_354
timestamp 1649977179
transform 1 0 33672 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1649977179
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_375
timestamp 1649977179
transform 1 0 35604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_381
timestamp 1649977179
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_388
timestamp 1649977179
transform 1 0 36800 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_403
timestamp 1649977179
transform 1 0 38180 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_3 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_15
timestamp 1649977179
transform 1 0 2484 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_23
timestamp 1649977179
transform 1 0 3220 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_26
timestamp 1649977179
transform 1 0 3496 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_34
timestamp 1649977179
transform 1 0 4232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_41
timestamp 1649977179
transform 1 0 4876 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_49
timestamp 1649977179
transform 1 0 5612 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_52
timestamp 1649977179
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_57 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_62
timestamp 1649977179
transform 1 0 6808 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_70
timestamp 1649977179
transform 1 0 7544 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_78 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 8280 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_82
timestamp 1649977179
transform 1 0 8648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_89
timestamp 1649977179
transform 1 0 9292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_96
timestamp 1649977179
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_102
timestamp 1649977179
transform 1 0 10488 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1649977179
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_118
timestamp 1649977179
transform 1 0 11960 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_126
timestamp 1649977179
transform 1 0 12696 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_134
timestamp 1649977179
transform 1 0 13432 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_138
timestamp 1649977179
transform 1 0 13800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_145
timestamp 1649977179
transform 1 0 14444 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_152
timestamp 1649977179
transform 1 0 15088 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_158
timestamp 1649977179
transform 1 0 15640 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_164
timestamp 1649977179
transform 1 0 16192 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_174
timestamp 1649977179
transform 1 0 17112 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_182
timestamp 1649977179
transform 1 0 17848 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_192
timestamp 1649977179
transform 1 0 18768 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_198
timestamp 1649977179
transform 1 0 19320 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_206
timestamp 1649977179
transform 1 0 20056 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_1_214
timestamp 1649977179
transform 1 0 20792 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_222
timestamp 1649977179
transform 1 0 21528 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_228
timestamp 1649977179
transform 1 0 22080 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_234
timestamp 1649977179
transform 1 0 22632 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_240
timestamp 1649977179
transform 1 0 23184 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_248
timestamp 1649977179
transform 1 0 23920 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_253
timestamp 1649977179
transform 1 0 24380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_257
timestamp 1649977179
transform 1 0 24748 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_260
timestamp 1649977179
transform 1 0 25024 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_266
timestamp 1649977179
transform 1 0 25576 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1649977179
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1649977179
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_283
timestamp 1649977179
transform 1 0 27140 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_1_289
timestamp 1649977179
transform 1 0 27692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_301
timestamp 1649977179
transform 1 0 28796 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_305
timestamp 1649977179
transform 1 0 29164 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_311
timestamp 1649977179
transform 1 0 29716 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_317
timestamp 1649977179
transform 1 0 30268 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_328
timestamp 1649977179
transform 1 0 31280 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_347
timestamp 1649977179
transform 1 0 33028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_361
timestamp 1649977179
transform 1 0 34316 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_375
timestamp 1649977179
transform 1 0 35604 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_383
timestamp 1649977179
transform 1 0 36340 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1649977179
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_393
timestamp 1649977179
transform 1 0 37260 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_397
timestamp 1649977179
transform 1 0 37628 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_402
timestamp 1649977179
transform 1 0 38088 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_406
timestamp 1649977179
transform 1 0 38456 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_2_47
timestamp 1649977179
transform 1 0 5428 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_59
timestamp 1649977179
transform 1 0 6532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_71
timestamp 1649977179
transform 1 0 7636 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1649977179
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1649977179
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1649977179
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1649977179
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1649977179
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1649977179
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1649977179
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1649977179
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_315
timestamp 1649977179
transform 1 0 30084 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_318
timestamp 1649977179
transform 1 0 30360 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_330
timestamp 1649977179
transform 1 0 31464 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_334
timestamp 1649977179
transform 1 0 31832 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_337
timestamp 1649977179
transform 1 0 32108 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_351
timestamp 1649977179
transform 1 0 33396 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1649977179
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_376
timestamp 1649977179
transform 1 0 35696 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_392
timestamp 1649977179
transform 1 0 37168 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_398
timestamp 1649977179
transform 1 0 37720 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_403
timestamp 1649977179
transform 1 0 38180 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1649977179
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1649977179
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1649977179
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1649977179
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1649977179
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1649977179
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1649977179
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1649977179
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_361
timestamp 1649977179
transform 1 0 34316 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_3_366
timestamp 1649977179
transform 1 0 34776 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_378
timestamp 1649977179
transform 1 0 35880 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_382
timestamp 1649977179
transform 1 0 36248 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_388
timestamp 1649977179
transform 1 0 36800 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_395
timestamp 1649977179
transform 1 0 37444 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_403
timestamp 1649977179
transform 1 0 38180 0 -1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1649977179
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1649977179
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1649977179
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1649977179
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1649977179
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1649977179
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1649977179
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1649977179
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1649977179
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1649977179
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1649977179
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1649977179
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_385
timestamp 1649977179
transform 1 0 36524 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_390
timestamp 1649977179
transform 1 0 36984 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_394
timestamp 1649977179
transform 1 0 37352 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_397
timestamp 1649977179
transform 1 0 37628 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_403
timestamp 1649977179
transform 1 0 38180 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_63
timestamp 1649977179
transform 1 0 6900 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_66
timestamp 1649977179
transform 1 0 7176 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_79
timestamp 1649977179
transform 1 0 8372 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_85
timestamp 1649977179
transform 1 0 8924 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_5_91
timestamp 1649977179
transform 1 0 9476 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_103
timestamp 1649977179
transform 1 0 10580 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1649977179
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1649977179
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1649977179
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1649977179
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1649977179
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1649977179
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1649977179
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1649977179
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1649977179
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1649977179
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1649977179
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_395
timestamp 1649977179
transform 1 0 37444 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_403
timestamp 1649977179
transform 1 0 38180 0 -1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_6_61
timestamp 1649977179
transform 1 0 6716 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_66
timestamp 1649977179
transform 1 0 7176 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp 1649977179
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_95
timestamp 1649977179
transform 1 0 9844 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_107
timestamp 1649977179
transform 1 0 10948 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_119
timestamp 1649977179
transform 1 0 12052 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_131
timestamp 1649977179
transform 1 0 13156 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1649977179
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1649977179
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1649977179
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1649977179
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1649977179
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1649977179
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1649977179
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1649977179
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1649977179
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_389
timestamp 1649977179
transform 1 0 36892 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_395
timestamp 1649977179
transform 1 0 37444 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_403
timestamp 1649977179
transform 1 0 38180 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_67
timestamp 1649977179
transform 1 0 7268 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_80
timestamp 1649977179
transform 1 0 8464 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_94
timestamp 1649977179
transform 1 0 9752 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_7_100
timestamp 1649977179
transform 1 0 10304 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1649977179
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1649977179
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1649977179
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1649977179
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1649977179
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1649977179
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1649977179
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_395
timestamp 1649977179
transform 1 0 37444 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_403
timestamp 1649977179
transform 1 0 38180 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_61
timestamp 1649977179
transform 1 0 6716 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_67
timestamp 1649977179
transform 1 0 7268 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_80
timestamp 1649977179
transform 1 0 8464 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_95
timestamp 1649977179
transform 1 0 9844 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1649977179
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1649977179
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1649977179
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1649977179
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1649977179
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1649977179
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1649977179
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1649977179
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1649977179
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1649977179
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1649977179
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1649977179
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_389
timestamp 1649977179
transform 1 0 36892 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_395
timestamp 1649977179
transform 1 0 37444 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_403
timestamp 1649977179
transform 1 0 38180 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_65
timestamp 1649977179
transform 1 0 7084 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_82
timestamp 1649977179
transform 1 0 8648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_86
timestamp 1649977179
transform 1 0 9016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_97
timestamp 1649977179
transform 1 0 10028 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_103
timestamp 1649977179
transform 1 0 10580 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1649977179
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1649977179
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1649977179
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1649977179
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1649977179
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1649977179
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1649977179
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1649977179
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1649977179
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1649977179
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1649977179
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_80
timestamp 1649977179
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_87
timestamp 1649977179
transform 1 0 9108 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_10_101
timestamp 1649977179
transform 1 0 10396 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_113
timestamp 1649977179
transform 1 0 11500 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_125
timestamp 1649977179
transform 1 0 12604 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_137
timestamp 1649977179
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1649977179
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1649977179
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1649977179
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1649977179
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1649977179
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1649977179
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1649977179
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1649977179
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1649977179
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1649977179
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1649977179
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1649977179
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1649977179
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_389
timestamp 1649977179
transform 1 0 36892 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_395
timestamp 1649977179
transform 1 0 37444 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_403
timestamp 1649977179
transform 1 0 38180 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_77
timestamp 1649977179
transform 1 0 8188 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_80
timestamp 1649977179
transform 1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_99
timestamp 1649977179
transform 1 0 10212 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1649977179
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1649977179
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1649977179
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1649977179
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1649977179
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1649977179
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1649977179
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1649977179
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1649977179
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1649977179
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1649977179
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_395
timestamp 1649977179
transform 1 0 37444 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_403
timestamp 1649977179
transform 1 0 38180 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1649977179
transform 1 0 9660 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_107
timestamp 1649977179
transform 1 0 10948 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_115
timestamp 1649977179
transform 1 0 11684 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_126
timestamp 1649977179
transform 1 0 12696 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_138
timestamp 1649977179
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1649977179
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1649977179
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1649977179
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1649977179
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1649977179
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1649977179
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1649977179
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1649977179
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1649977179
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1649977179
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1649977179
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1649977179
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1649977179
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_389
timestamp 1649977179
transform 1 0 36892 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_395
timestamp 1649977179
transform 1 0 37444 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_403
timestamp 1649977179
transform 1 0 38180 0 1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_94
timestamp 1649977179
transform 1 0 9752 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_108
timestamp 1649977179
transform 1 0 11040 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_117
timestamp 1649977179
transform 1 0 11868 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_120
timestamp 1649977179
transform 1 0 12144 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_13_134
timestamp 1649977179
transform 1 0 13432 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_146
timestamp 1649977179
transform 1 0 14536 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_158
timestamp 1649977179
transform 1 0 15640 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_166
timestamp 1649977179
transform 1 0 16376 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1649977179
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1649977179
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1649977179
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1649977179
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1649977179
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1649977179
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1649977179
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1649977179
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1649977179
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1649977179
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1649977179
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1649977179
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_395
timestamp 1649977179
transform 1 0 37444 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_403
timestamp 1649977179
transform 1 0 38180 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_93
timestamp 1649977179
transform 1 0 9660 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_106
timestamp 1649977179
transform 1 0 10856 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_120
timestamp 1649977179
transform 1 0 12144 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_143
timestamp 1649977179
transform 1 0 14260 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_155
timestamp 1649977179
transform 1 0 15364 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_167
timestamp 1649977179
transform 1 0 16468 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_179
timestamp 1649977179
transform 1 0 17572 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_191
timestamp 1649977179
transform 1 0 18676 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1649977179
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1649977179
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1649977179
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1649977179
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1649977179
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1649977179
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1649977179
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1649977179
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1649977179
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1649977179
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1649977179
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1649977179
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_96
timestamp 1649977179
transform 1 0 9936 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_102
timestamp 1649977179
transform 1 0 10488 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_108
timestamp 1649977179
transform 1 0 11040 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_122
timestamp 1649977179
transform 1 0 12328 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_131
timestamp 1649977179
transform 1 0 13156 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_138
timestamp 1649977179
transform 1 0 13800 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_144
timestamp 1649977179
transform 1 0 14352 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_15_150
timestamp 1649977179
transform 1 0 14904 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_162
timestamp 1649977179
transform 1 0 16008 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1649977179
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1649977179
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1649977179
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1649977179
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1649977179
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1649977179
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1649977179
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1649977179
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1649977179
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1649977179
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1649977179
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1649977179
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1649977179
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_395
timestamp 1649977179
transform 1 0 37444 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_403
timestamp 1649977179
transform 1 0 38180 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_113
timestamp 1649977179
transform 1 0 11500 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_119
timestamp 1649977179
transform 1 0 12052 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_16_132
timestamp 1649977179
transform 1 0 13248 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_16_144
timestamp 1649977179
transform 1 0 14352 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_156
timestamp 1649977179
transform 1 0 15456 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_168
timestamp 1649977179
transform 1 0 16560 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_180
timestamp 1649977179
transform 1 0 17664 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1649977179
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1649977179
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1649977179
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1649977179
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1649977179
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1649977179
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1649977179
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1649977179
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1649977179
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1649977179
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1649977179
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1649977179
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1649977179
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1649977179
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1649977179
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_389
timestamp 1649977179
transform 1 0 36892 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_395
timestamp 1649977179
transform 1 0 37444 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_403
timestamp 1649977179
transform 1 0 38180 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1649977179
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_121
timestamp 1649977179
transform 1 0 12236 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_134
timestamp 1649977179
transform 1 0 13432 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_17_141
timestamp 1649977179
transform 1 0 14076 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_153
timestamp 1649977179
transform 1 0 15180 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_17_165
timestamp 1649977179
transform 1 0 16284 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1649977179
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1649977179
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1649977179
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1649977179
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1649977179
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1649977179
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1649977179
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1649977179
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1649977179
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1649977179
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1649977179
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_395
timestamp 1649977179
transform 1 0 37444 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_403
timestamp 1649977179
transform 1 0 38180 0 -1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_134
timestamp 1649977179
transform 1 0 13432 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_144
timestamp 1649977179
transform 1 0 14352 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_18_150
timestamp 1649977179
transform 1 0 14904 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_162
timestamp 1649977179
transform 1 0 16008 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_174
timestamp 1649977179
transform 1 0 17112 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_186
timestamp 1649977179
transform 1 0 18216 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_194
timestamp 1649977179
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1649977179
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1649977179
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1649977179
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1649977179
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1649977179
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1649977179
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1649977179
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1649977179
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1649977179
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1649977179
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1649977179
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1649977179
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_389
timestamp 1649977179
transform 1 0 36892 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_395
timestamp 1649977179
transform 1 0 37444 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_403
timestamp 1649977179
transform 1 0 38180 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_127
timestamp 1649977179
transform 1 0 12788 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_140
timestamp 1649977179
transform 1 0 13984 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_147
timestamp 1649977179
transform 1 0 14628 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_153
timestamp 1649977179
transform 1 0 15180 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_165
timestamp 1649977179
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1649977179
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1649977179
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1649977179
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1649977179
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1649977179
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1649977179
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1649977179
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1649977179
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1649977179
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1649977179
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1649977179
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1649977179
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1649977179
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1649977179
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_393
timestamp 1649977179
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_405
timestamp 1649977179
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_117
timestamp 1649977179
transform 1 0 11868 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_125
timestamp 1649977179
transform 1 0 12604 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_131
timestamp 1649977179
transform 1 0 13156 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_150
timestamp 1649977179
transform 1 0 14904 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_20_157
timestamp 1649977179
transform 1 0 15548 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_169
timestamp 1649977179
transform 1 0 16652 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_181
timestamp 1649977179
transform 1 0 17756 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1649977179
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1649977179
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1649977179
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1649977179
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1649977179
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1649977179
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1649977179
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1649977179
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1649977179
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1649977179
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1649977179
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1649977179
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1649977179
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1649977179
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_389
timestamp 1649977179
transform 1 0 36892 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_395
timestamp 1649977179
transform 1 0 37444 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_403
timestamp 1649977179
transform 1 0 38180 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_129
timestamp 1649977179
transform 1 0 12972 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_141
timestamp 1649977179
transform 1 0 14076 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_152
timestamp 1649977179
transform 1 0 15088 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_158
timestamp 1649977179
transform 1 0 15640 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_166
timestamp 1649977179
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1649977179
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1649977179
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1649977179
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1649977179
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1649977179
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1649977179
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1649977179
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1649977179
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1649977179
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1649977179
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1649977179
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1649977179
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1649977179
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1649977179
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1649977179
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_395
timestamp 1649977179
transform 1 0 37444 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_403
timestamp 1649977179
transform 1 0 38180 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_156
timestamp 1649977179
transform 1 0 15456 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_163
timestamp 1649977179
transform 1 0 16100 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_22_169
timestamp 1649977179
transform 1 0 16652 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_181
timestamp 1649977179
transform 1 0 17756 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_193
timestamp 1649977179
transform 1 0 18860 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1649977179
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1649977179
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1649977179
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1649977179
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1649977179
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1649977179
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1649977179
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1649977179
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1649977179
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1649977179
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1649977179
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_389
timestamp 1649977179
transform 1 0 36892 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_395
timestamp 1649977179
transform 1 0 37444 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_403
timestamp 1649977179
transform 1 0 38180 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1649977179
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_172
timestamp 1649977179
transform 1 0 16928 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_23_178
timestamp 1649977179
transform 1 0 17480 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_190
timestamp 1649977179
transform 1 0 18584 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_202
timestamp 1649977179
transform 1 0 19688 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_214
timestamp 1649977179
transform 1 0 20792 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_222
timestamp 1649977179
transform 1 0 21528 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1649977179
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1649977179
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1649977179
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1649977179
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1649977179
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1649977179
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1649977179
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1649977179
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1649977179
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1649977179
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1649977179
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1649977179
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_395
timestamp 1649977179
transform 1 0 37444 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_403
timestamp 1649977179
transform 1 0 38180 0 -1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_161
timestamp 1649977179
transform 1 0 15916 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_171
timestamp 1649977179
transform 1 0 16836 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_178
timestamp 1649977179
transform 1 0 17480 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_24_184
timestamp 1649977179
transform 1 0 18032 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1649977179
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1649977179
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1649977179
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1649977179
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1649977179
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1649977179
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1649977179
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1649977179
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1649977179
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1649977179
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1649977179
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1649977179
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1649977179
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1649977179
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_179
timestamp 1649977179
transform 1 0 17572 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_25_186
timestamp 1649977179
transform 1 0 18216 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_198
timestamp 1649977179
transform 1 0 19320 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_210
timestamp 1649977179
transform 1 0 20424 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1649977179
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1649977179
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1649977179
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1649977179
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1649977179
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1649977179
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1649977179
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1649977179
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1649977179
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1649977179
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1649977179
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1649977179
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1649977179
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_395
timestamp 1649977179
transform 1 0 37444 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_403
timestamp 1649977179
transform 1 0 38180 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_188
timestamp 1649977179
transform 1 0 18400 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_199
timestamp 1649977179
transform 1 0 19412 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_211
timestamp 1649977179
transform 1 0 20516 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_26_217
timestamp 1649977179
transform 1 0 21068 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_229
timestamp 1649977179
transform 1 0 22172 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_241
timestamp 1649977179
transform 1 0 23276 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_249
timestamp 1649977179
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1649977179
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1649977179
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1649977179
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1649977179
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1649977179
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1649977179
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1649977179
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1649977179
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1649977179
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_389
timestamp 1649977179
transform 1 0 36892 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_395
timestamp 1649977179
transform 1 0 37444 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_403
timestamp 1649977179
transform 1 0 38180 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1649977179
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_27_188
timestamp 1649977179
transform 1 0 18400 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_200
timestamp 1649977179
transform 1 0 19504 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_212
timestamp 1649977179
transform 1 0 20608 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1649977179
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1649977179
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1649977179
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1649977179
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1649977179
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1649977179
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1649977179
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1649977179
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1649977179
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1649977179
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1649977179
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1649977179
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1649977179
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_395
timestamp 1649977179
transform 1 0 37444 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_403
timestamp 1649977179
transform 1 0 38180 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1649977179
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_201
timestamp 1649977179
transform 1 0 19596 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_28_207
timestamp 1649977179
transform 1 0 20148 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_219
timestamp 1649977179
transform 1 0 21252 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_231
timestamp 1649977179
transform 1 0 22356 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_243
timestamp 1649977179
transform 1 0 23460 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1649977179
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1649977179
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1649977179
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1649977179
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1649977179
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1649977179
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1649977179
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1649977179
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1649977179
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1649977179
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_389
timestamp 1649977179
transform 1 0 36892 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_395
timestamp 1649977179
transform 1 0 37444 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_403
timestamp 1649977179
transform 1 0 38180 0 1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_3
timestamp 1649977179
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_15
timestamp 1649977179
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_27
timestamp 1649977179
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_39
timestamp 1649977179
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_51
timestamp 1649977179
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_55
timestamp 1649977179
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_191
timestamp 1649977179
transform 1 0 18676 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_204
timestamp 1649977179
transform 1 0 19872 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_211
timestamp 1649977179
transform 1 0 20516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1649977179
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1649977179
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1649977179
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1649977179
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1649977179
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1649977179
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1649977179
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1649977179
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1649977179
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1649977179
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1649977179
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1649977179
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1649977179
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1649977179
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1649977179
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_201
timestamp 1649977179
transform 1 0 19596 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_211
timestamp 1649977179
transform 1 0 20516 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_30_218
timestamp 1649977179
transform 1 0 21160 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_230
timestamp 1649977179
transform 1 0 22264 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_242
timestamp 1649977179
transform 1 0 23368 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_250
timestamp 1649977179
transform 1 0 24104 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1649977179
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1649977179
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1649977179
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1649977179
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1649977179
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1649977179
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1649977179
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1649977179
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1649977179
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1649977179
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_389
timestamp 1649977179
transform 1 0 36892 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_397
timestamp 1649977179
transform 1 0 37628 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_403
timestamp 1649977179
transform 1 0 38180 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_203
timestamp 1649977179
transform 1 0 19780 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_213
timestamp 1649977179
transform 1 0 20700 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1649977179
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1649977179
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1649977179
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1649977179
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1649977179
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1649977179
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1649977179
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1649977179
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1649977179
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1649977179
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1649977179
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1649977179
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1649977179
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_393
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_403
timestamp 1649977179
transform 1 0 38180 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1649977179
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1649977179
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_205
timestamp 1649977179
transform 1 0 19964 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_32_219
timestamp 1649977179
transform 1 0 21252 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_32_228
timestamp 1649977179
transform 1 0 22080 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_240
timestamp 1649977179
transform 1 0 23184 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1649977179
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1649977179
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1649977179
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1649977179
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1649977179
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1649977179
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1649977179
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1649977179
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1649977179
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1649977179
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_389
timestamp 1649977179
transform 1 0 36892 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_397
timestamp 1649977179
transform 1 0 37628 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_403
timestamp 1649977179
transform 1 0 38180 0 1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1649977179
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_205
timestamp 1649977179
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_217
timestamp 1649977179
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1649977179
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_234
timestamp 1649977179
transform 1 0 22632 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_241
timestamp 1649977179
transform 1 0 23276 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_247
timestamp 1649977179
transform 1 0 23828 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_259
timestamp 1649977179
transform 1 0 24932 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_271
timestamp 1649977179
transform 1 0 26036 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1649977179
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1649977179
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1649977179
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1649977179
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1649977179
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1649977179
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1649977179
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1649977179
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1649977179
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1649977179
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1649977179
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_393
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_33_403
timestamp 1649977179
transform 1 0 38180 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1649977179
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1649977179
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1649977179
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1649977179
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1649977179
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_189
timestamp 1649977179
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1649977179
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_209
timestamp 1649977179
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_221
timestamp 1649977179
transform 1 0 21436 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_225
timestamp 1649977179
transform 1 0 21804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_232
timestamp 1649977179
transform 1 0 22448 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_241
timestamp 1649977179
transform 1 0 23276 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_247
timestamp 1649977179
transform 1 0 23828 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_251
timestamp 1649977179
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1649977179
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1649977179
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1649977179
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1649977179
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1649977179
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1649977179
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1649977179
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1649977179
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1649977179
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1649977179
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1649977179
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1649977179
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1649977179
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1649977179
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1649977179
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1649977179
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1649977179
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1649977179
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1649977179
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1649977179
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_181
timestamp 1649977179
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_193
timestamp 1649977179
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_205
timestamp 1649977179
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_217
timestamp 1649977179
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1649977179
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_225
timestamp 1649977179
transform 1 0 21804 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_233
timestamp 1649977179
transform 1 0 22540 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_243
timestamp 1649977179
transform 1 0 23460 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_250
timestamp 1649977179
transform 1 0 24104 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_262
timestamp 1649977179
transform 1 0 25208 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_274
timestamp 1649977179
transform 1 0 26312 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1649977179
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1649977179
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1649977179
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1649977179
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1649977179
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1649977179
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1649977179
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1649977179
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1649977179
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_396
timestamp 1649977179
transform 1 0 37536 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_403
timestamp 1649977179
transform 1 0 38180 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1649977179
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1649977179
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1649977179
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1649977179
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1649977179
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1649977179
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1649977179
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1649977179
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1649977179
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_165
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_177
timestamp 1649977179
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_189
timestamp 1649977179
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_195
timestamp 1649977179
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_209
timestamp 1649977179
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_221
timestamp 1649977179
transform 1 0 21436 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_229
timestamp 1649977179
transform 1 0 22172 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_233
timestamp 1649977179
transform 1 0 22540 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_241
timestamp 1649977179
transform 1 0 23276 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_36_245
timestamp 1649977179
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_251
timestamp 1649977179
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_255
timestamp 1649977179
transform 1 0 24564 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_267
timestamp 1649977179
transform 1 0 25668 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_279
timestamp 1649977179
transform 1 0 26772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_291
timestamp 1649977179
transform 1 0 27876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_303
timestamp 1649977179
transform 1 0 28980 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1649977179
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1649977179
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1649977179
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1649977179
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1649977179
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1649977179
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1649977179
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_389
timestamp 1649977179
transform 1 0 36892 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_397
timestamp 1649977179
transform 1 0 37628 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_403
timestamp 1649977179
transform 1 0 38180 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1649977179
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1649977179
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1649977179
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1649977179
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1649977179
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1649977179
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1649977179
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1649977179
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1649977179
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_149
timestamp 1649977179
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1649977179
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_181
timestamp 1649977179
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_193
timestamp 1649977179
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_205
timestamp 1649977179
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_217
timestamp 1649977179
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_223
timestamp 1649977179
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_225
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_237
timestamp 1649977179
transform 1 0 22908 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_241
timestamp 1649977179
transform 1 0 23276 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_251
timestamp 1649977179
transform 1 0 24196 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_258
timestamp 1649977179
transform 1 0 24840 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_264
timestamp 1649977179
transform 1 0 25392 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_276
timestamp 1649977179
transform 1 0 26496 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1649977179
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1649977179
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1649977179
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1649977179
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1649977179
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1649977179
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1649977179
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1649977179
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_375
timestamp 1649977179
transform 1 0 35604 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_388
timestamp 1649977179
transform 1 0 36800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_395
timestamp 1649977179
transform 1 0 37444 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_403
timestamp 1649977179
transform 1 0 38180 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1649977179
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1649977179
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1649977179
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1649977179
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_121
timestamp 1649977179
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_133
timestamp 1649977179
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_153
timestamp 1649977179
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_165
timestamp 1649977179
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_177
timestamp 1649977179
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_189
timestamp 1649977179
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1649977179
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_197
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_209
timestamp 1649977179
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_221
timestamp 1649977179
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_233
timestamp 1649977179
transform 1 0 22540 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_243
timestamp 1649977179
transform 1 0 23460 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1649977179
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_262
timestamp 1649977179
transform 1 0 25208 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_269
timestamp 1649977179
transform 1 0 25852 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_38_275
timestamp 1649977179
transform 1 0 26404 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_287
timestamp 1649977179
transform 1 0 27508 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_299
timestamp 1649977179
transform 1 0 28612 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1649977179
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1649977179
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1649977179
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1649977179
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1649977179
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1649977179
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_377
timestamp 1649977179
transform 1 0 35788 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_385
timestamp 1649977179
transform 1 0 36524 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_391
timestamp 1649977179
transform 1 0 37076 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_403
timestamp 1649977179
transform 1 0 38180 0 1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1649977179
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1649977179
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1649977179
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1649977179
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1649977179
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1649977179
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1649977179
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1649977179
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_137
timestamp 1649977179
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_149
timestamp 1649977179
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1649977179
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_169
timestamp 1649977179
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_181
timestamp 1649977179
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_193
timestamp 1649977179
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_205
timestamp 1649977179
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1649977179
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1649977179
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_225
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_237
timestamp 1649977179
transform 1 0 22908 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_245
timestamp 1649977179
transform 1 0 23644 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_257
timestamp 1649977179
transform 1 0 24748 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_267
timestamp 1649977179
transform 1 0 25668 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_274
timestamp 1649977179
transform 1 0 26312 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1649977179
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1649977179
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1649977179
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1649977179
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1649977179
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1649977179
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1649977179
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1649977179
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1649977179
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1649977179
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1649977179
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1649977179
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1649977179
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1649977179
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1649977179
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1649977179
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1649977179
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1649977179
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1649977179
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_121
timestamp 1649977179
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_133
timestamp 1649977179
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1649977179
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_141
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_153
timestamp 1649977179
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_165
timestamp 1649977179
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_177
timestamp 1649977179
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_189
timestamp 1649977179
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1649977179
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_197
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_209
timestamp 1649977179
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_221
timestamp 1649977179
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_233
timestamp 1649977179
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1649977179
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1649977179
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_253
timestamp 1649977179
transform 1 0 24380 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_261
timestamp 1649977179
transform 1 0 25116 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_273
timestamp 1649977179
transform 1 0 26220 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_280
timestamp 1649977179
transform 1 0 26864 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_292
timestamp 1649977179
transform 1 0 27968 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1649977179
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1649977179
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1649977179
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1649977179
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1649977179
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1649977179
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_389
timestamp 1649977179
transform 1 0 36892 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_397
timestamp 1649977179
transform 1 0 37628 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_403
timestamp 1649977179
transform 1 0 38180 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1649977179
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1649977179
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1649977179
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1649977179
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1649977179
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_81
timestamp 1649977179
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_93
timestamp 1649977179
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_105
timestamp 1649977179
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1649977179
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_125
timestamp 1649977179
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_137
timestamp 1649977179
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_149
timestamp 1649977179
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_161
timestamp 1649977179
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1649977179
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_169
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_181
timestamp 1649977179
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_193
timestamp 1649977179
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_205
timestamp 1649977179
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_217
timestamp 1649977179
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_223
timestamp 1649977179
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_225
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_237
timestamp 1649977179
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_249
timestamp 1649977179
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_261
timestamp 1649977179
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_275
timestamp 1649977179
transform 1 0 26404 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_279
timestamp 1649977179
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_289
timestamp 1649977179
transform 1 0 27692 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_294
timestamp 1649977179
transform 1 0 28152 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_306
timestamp 1649977179
transform 1 0 29256 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_318
timestamp 1649977179
transform 1 0 30360 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_330
timestamp 1649977179
transform 1 0 31464 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1649977179
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1649977179
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1649977179
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1649977179
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1649977179
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_403
timestamp 1649977179
transform 1 0 38180 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1649977179
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1649977179
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1649977179
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1649977179
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_97
timestamp 1649977179
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_109
timestamp 1649977179
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_121
timestamp 1649977179
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1649977179
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1649977179
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_153
timestamp 1649977179
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_165
timestamp 1649977179
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_177
timestamp 1649977179
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_189
timestamp 1649977179
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1649977179
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_209
timestamp 1649977179
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_221
timestamp 1649977179
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_233
timestamp 1649977179
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1649977179
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1649977179
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1649977179
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_277
timestamp 1649977179
transform 1 0 26588 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_292
timestamp 1649977179
transform 1 0 27968 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_299
timestamp 1649977179
transform 1 0 28612 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1649977179
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1649977179
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1649977179
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1649977179
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1649977179
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1649977179
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1649977179
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_389
timestamp 1649977179
transform 1 0 36892 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_42_397
timestamp 1649977179
transform 1 0 37628 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_403
timestamp 1649977179
transform 1 0 38180 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1649977179
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1649977179
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1649977179
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1649977179
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1649977179
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_69
timestamp 1649977179
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_81
timestamp 1649977179
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_93
timestamp 1649977179
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_105
timestamp 1649977179
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1649977179
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_125
timestamp 1649977179
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_137
timestamp 1649977179
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_149
timestamp 1649977179
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_161
timestamp 1649977179
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1649977179
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_181
timestamp 1649977179
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_193
timestamp 1649977179
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_205
timestamp 1649977179
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_217
timestamp 1649977179
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_223
timestamp 1649977179
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_225
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_237
timestamp 1649977179
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_249
timestamp 1649977179
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_261
timestamp 1649977179
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_273
timestamp 1649977179
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_279
timestamp 1649977179
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_290
timestamp 1649977179
transform 1 0 27784 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_297
timestamp 1649977179
transform 1 0 28428 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_304
timestamp 1649977179
transform 1 0 29072 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_310
timestamp 1649977179
transform 1 0 29624 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_322
timestamp 1649977179
transform 1 0 30728 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_334
timestamp 1649977179
transform 1 0 31832 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1649977179
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1649977179
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1649977179
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1649977179
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1649977179
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_403
timestamp 1649977179
transform 1 0 38180 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_3
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_15
timestamp 1649977179
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1649977179
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_29
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_41
timestamp 1649977179
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_53
timestamp 1649977179
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_65
timestamp 1649977179
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_77
timestamp 1649977179
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_83
timestamp 1649977179
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_85
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_97
timestamp 1649977179
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_109
timestamp 1649977179
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_121
timestamp 1649977179
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_133
timestamp 1649977179
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_139
timestamp 1649977179
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_165
timestamp 1649977179
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_177
timestamp 1649977179
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_189
timestamp 1649977179
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1649977179
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_209
timestamp 1649977179
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_221
timestamp 1649977179
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_233
timestamp 1649977179
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_245
timestamp 1649977179
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_251
timestamp 1649977179
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1649977179
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1649977179
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_289
timestamp 1649977179
transform 1 0 27692 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_44_299
timestamp 1649977179
transform 1 0 28612 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1649977179
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_311
timestamp 1649977179
transform 1 0 29716 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_323
timestamp 1649977179
transform 1 0 30820 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_335
timestamp 1649977179
transform 1 0 31924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_347
timestamp 1649977179
transform 1 0 33028 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_359
timestamp 1649977179
transform 1 0 34132 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1649977179
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1649977179
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1649977179
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1649977179
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1649977179
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1649977179
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1649977179
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1649977179
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1649977179
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_69
timestamp 1649977179
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_81
timestamp 1649977179
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_93
timestamp 1649977179
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1649977179
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1649977179
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_113
timestamp 1649977179
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_125
timestamp 1649977179
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_137
timestamp 1649977179
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_149
timestamp 1649977179
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_161
timestamp 1649977179
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1649977179
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_169
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_181
timestamp 1649977179
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_193
timestamp 1649977179
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_205
timestamp 1649977179
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_217
timestamp 1649977179
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1649977179
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_225
timestamp 1649977179
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_237
timestamp 1649977179
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_249
timestamp 1649977179
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_261
timestamp 1649977179
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_273
timestamp 1649977179
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1649977179
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_293
timestamp 1649977179
transform 1 0 28060 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_297
timestamp 1649977179
transform 1 0 28428 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_307
timestamp 1649977179
transform 1 0 29348 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_314
timestamp 1649977179
transform 1 0 29992 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_320
timestamp 1649977179
transform 1 0 30544 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_332
timestamp 1649977179
transform 1 0 31648 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1649977179
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1649977179
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1649977179
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1649977179
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1649977179
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_403
timestamp 1649977179
transform 1 0 38180 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_3
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_15
timestamp 1649977179
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_27
timestamp 1649977179
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1649977179
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_65
timestamp 1649977179
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_77
timestamp 1649977179
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_83
timestamp 1649977179
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_85
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_97
timestamp 1649977179
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_109
timestamp 1649977179
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_121
timestamp 1649977179
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1649977179
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1649977179
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_141
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_153
timestamp 1649977179
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_165
timestamp 1649977179
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_177
timestamp 1649977179
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_189
timestamp 1649977179
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_195
timestamp 1649977179
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_209
timestamp 1649977179
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_221
timestamp 1649977179
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_233
timestamp 1649977179
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_245
timestamp 1649977179
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_251
timestamp 1649977179
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1649977179
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1649977179
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_289
timestamp 1649977179
transform 1 0 27692 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_297
timestamp 1649977179
transform 1 0 28428 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1649977179
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1649977179
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_309
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_316
timestamp 1649977179
transform 1 0 30176 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_322
timestamp 1649977179
transform 1 0 30728 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_334
timestamp 1649977179
transform 1 0 31832 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_346
timestamp 1649977179
transform 1 0 32936 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_358
timestamp 1649977179
transform 1 0 34040 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1649977179
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_389
timestamp 1649977179
transform 1 0 36892 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_397
timestamp 1649977179
transform 1 0 37628 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_403
timestamp 1649977179
transform 1 0 38180 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_15
timestamp 1649977179
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_27
timestamp 1649977179
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_39
timestamp 1649977179
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1649977179
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1649977179
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1649977179
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_81
timestamp 1649977179
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_93
timestamp 1649977179
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_105
timestamp 1649977179
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1649977179
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_113
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_125
timestamp 1649977179
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_137
timestamp 1649977179
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_149
timestamp 1649977179
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_161
timestamp 1649977179
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1649977179
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_181
timestamp 1649977179
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_193
timestamp 1649977179
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_205
timestamp 1649977179
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_217
timestamp 1649977179
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1649977179
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1649977179
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1649977179
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1649977179
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1649977179
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1649977179
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_299
timestamp 1649977179
transform 1 0 28612 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_305
timestamp 1649977179
transform 1 0 29164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_315
timestamp 1649977179
transform 1 0 30084 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_325
timestamp 1649977179
transform 1 0 31004 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_331
timestamp 1649977179
transform 1 0 31556 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1649977179
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1649977179
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1649977179
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1649977179
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1649977179
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1649977179
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1649977179
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_393
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_403
timestamp 1649977179
transform 1 0 38180 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1649977179
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_41
timestamp 1649977179
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_53
timestamp 1649977179
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1649977179
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1649977179
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1649977179
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_85
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_97
timestamp 1649977179
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_109
timestamp 1649977179
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_121
timestamp 1649977179
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_133
timestamp 1649977179
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_139
timestamp 1649977179
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_153
timestamp 1649977179
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_165
timestamp 1649977179
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_177
timestamp 1649977179
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_189
timestamp 1649977179
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_195
timestamp 1649977179
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_197
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1649977179
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1649977179
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1649977179
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1649977179
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1649977179
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1649977179
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1649977179
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1649977179
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1649977179
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1649977179
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_309
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_313
timestamp 1649977179
transform 1 0 29900 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_323
timestamp 1649977179
transform 1 0 30820 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_330
timestamp 1649977179
transform 1 0 31464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_336
timestamp 1649977179
transform 1 0 32016 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_342
timestamp 1649977179
transform 1 0 32568 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_354
timestamp 1649977179
transform 1 0 33672 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_362
timestamp 1649977179
transform 1 0 34408 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1649977179
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1649977179
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_389
timestamp 1649977179
transform 1 0 36892 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_397
timestamp 1649977179
transform 1 0 37628 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_403
timestamp 1649977179
transform 1 0 38180 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1649977179
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1649977179
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1649977179
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1649977179
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1649977179
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1649977179
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_69
timestamp 1649977179
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_81
timestamp 1649977179
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_93
timestamp 1649977179
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_105
timestamp 1649977179
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1649977179
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_113
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_125
timestamp 1649977179
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_137
timestamp 1649977179
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_149
timestamp 1649977179
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_161
timestamp 1649977179
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_167
timestamp 1649977179
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_169
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_181
timestamp 1649977179
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_193
timestamp 1649977179
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1649977179
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1649977179
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1649977179
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1649977179
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1649977179
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1649977179
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1649977179
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1649977179
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1649977179
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1649977179
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_317
timestamp 1649977179
transform 1 0 30268 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_321
timestamp 1649977179
transform 1 0 30636 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_331
timestamp 1649977179
transform 1 0 31556 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1649977179
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_340
timestamp 1649977179
transform 1 0 32384 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_347
timestamp 1649977179
transform 1 0 33028 0 -1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_355
timestamp 1649977179
transform 1 0 33764 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_367
timestamp 1649977179
transform 1 0 34868 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_379
timestamp 1649977179
transform 1 0 35972 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1649977179
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1649977179
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1649977179
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1649977179
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1649977179
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1649977179
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1649977179
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1649977179
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1649977179
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1649977179
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1649977179
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_109
timestamp 1649977179
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_121
timestamp 1649977179
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_133
timestamp 1649977179
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1649977179
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_153
timestamp 1649977179
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_165
timestamp 1649977179
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_177
timestamp 1649977179
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_189
timestamp 1649977179
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1649977179
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_197
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_209
timestamp 1649977179
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_221
timestamp 1649977179
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_233
timestamp 1649977179
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_245
timestamp 1649977179
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_251
timestamp 1649977179
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1649977179
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1649977179
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1649977179
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1649977179
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1649977179
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1649977179
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_321
timestamp 1649977179
transform 1 0 30636 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_329
timestamp 1649977179
transform 1 0 31372 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_340
timestamp 1649977179
transform 1 0 32384 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_353
timestamp 1649977179
transform 1 0 33580 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_359
timestamp 1649977179
transform 1 0 34132 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1649977179
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1649977179
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1649977179
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_389
timestamp 1649977179
transform 1 0 36892 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_397
timestamp 1649977179
transform 1 0 37628 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_403
timestamp 1649977179
transform 1 0 38180 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1649977179
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1649977179
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1649977179
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1649977179
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1649977179
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1649977179
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_81
timestamp 1649977179
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_93
timestamp 1649977179
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_105
timestamp 1649977179
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_111
timestamp 1649977179
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1649977179
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1649977179
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1649977179
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1649977179
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1649977179
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_169
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_181
timestamp 1649977179
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_193
timestamp 1649977179
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1649977179
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1649977179
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1649977179
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1649977179
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1649977179
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1649977179
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1649977179
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1649977179
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1649977179
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1649977179
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1649977179
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1649977179
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1649977179
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_347
timestamp 1649977179
transform 1 0 33028 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_354
timestamp 1649977179
transform 1 0 33672 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1649977179
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1649977179
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1649977179
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1649977179
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_393
timestamp 1649977179
transform 1 0 37260 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_403
timestamp 1649977179
transform 1 0 38180 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1649977179
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1649977179
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1649977179
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1649977179
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1649977179
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1649977179
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1649977179
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_85
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_97
timestamp 1649977179
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_109
timestamp 1649977179
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_121
timestamp 1649977179
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_133
timestamp 1649977179
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_139
timestamp 1649977179
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_141
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_153
timestamp 1649977179
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_165
timestamp 1649977179
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_177
timestamp 1649977179
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1649977179
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1649977179
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_197
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_209
timestamp 1649977179
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_221
timestamp 1649977179
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_233
timestamp 1649977179
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_245
timestamp 1649977179
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_251
timestamp 1649977179
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1649977179
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1649977179
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1649977179
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1649977179
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1649977179
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1649977179
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1649977179
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_345
timestamp 1649977179
transform 1 0 32844 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_349
timestamp 1649977179
transform 1 0 33212 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_361
timestamp 1649977179
transform 1 0 34316 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1649977179
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_389
timestamp 1649977179
transform 1 0 36892 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_397
timestamp 1649977179
transform 1 0 37628 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_403
timestamp 1649977179
transform 1 0 38180 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_3
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_15
timestamp 1649977179
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_27
timestamp 1649977179
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_39
timestamp 1649977179
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_51
timestamp 1649977179
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1649977179
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_69
timestamp 1649977179
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_81
timestamp 1649977179
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_93
timestamp 1649977179
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1649977179
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1649977179
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1649977179
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1649977179
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1649977179
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1649977179
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1649977179
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_169
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_181
timestamp 1649977179
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_193
timestamp 1649977179
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_205
timestamp 1649977179
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_217
timestamp 1649977179
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1649977179
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1649977179
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1649977179
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1649977179
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1649977179
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1649977179
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1649977179
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1649977179
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1649977179
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1649977179
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1649977179
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_349
timestamp 1649977179
transform 1 0 33212 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_357
timestamp 1649977179
transform 1 0 33948 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_362
timestamp 1649977179
transform 1 0 34408 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_368
timestamp 1649977179
transform 1 0 34960 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_380
timestamp 1649977179
transform 1 0 36064 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_393
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_403
timestamp 1649977179
transform 1 0 38180 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1649977179
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1649977179
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1649977179
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1649977179
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1649977179
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1649977179
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_97
timestamp 1649977179
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1649977179
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1649977179
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1649977179
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1649977179
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_141
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_153
timestamp 1649977179
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_165
timestamp 1649977179
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_177
timestamp 1649977179
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1649977179
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1649977179
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_197
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_209
timestamp 1649977179
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_221
timestamp 1649977179
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_233
timestamp 1649977179
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_245
timestamp 1649977179
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1649977179
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1649977179
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1649977179
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1649977179
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1649977179
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1649977179
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1649977179
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1649977179
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1649977179
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_345
timestamp 1649977179
transform 1 0 32844 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_360
timestamp 1649977179
transform 1 0 34224 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_368
timestamp 1649977179
transform 1 0 34960 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_374
timestamp 1649977179
transform 1 0 35512 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_386
timestamp 1649977179
transform 1 0 36616 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_398
timestamp 1649977179
transform 1 0 37720 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_403
timestamp 1649977179
transform 1 0 38180 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1649977179
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1649977179
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1649977179
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1649977179
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1649977179
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1649977179
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1649977179
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1649977179
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1649977179
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1649977179
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1649977179
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1649977179
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_137
timestamp 1649977179
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_149
timestamp 1649977179
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_161
timestamp 1649977179
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1649977179
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_169
timestamp 1649977179
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_181
timestamp 1649977179
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_193
timestamp 1649977179
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_205
timestamp 1649977179
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1649977179
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1649977179
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1649977179
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1649977179
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1649977179
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1649977179
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1649977179
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1649977179
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1649977179
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1649977179
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1649977179
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1649977179
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_349
timestamp 1649977179
transform 1 0 33212 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_355
timestamp 1649977179
transform 1 0 33764 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_358
timestamp 1649977179
transform 1 0 34040 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_371
timestamp 1649977179
transform 1 0 35236 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_378
timestamp 1649977179
transform 1 0 35880 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_390
timestamp 1649977179
transform 1 0 36984 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_395
timestamp 1649977179
transform 1 0 37444 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_403
timestamp 1649977179
transform 1 0 38180 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1649977179
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1649977179
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1649977179
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1649977179
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1649977179
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1649977179
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1649977179
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_109
timestamp 1649977179
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_121
timestamp 1649977179
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_133
timestamp 1649977179
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_139
timestamp 1649977179
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_141
timestamp 1649977179
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_153
timestamp 1649977179
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_165
timestamp 1649977179
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_177
timestamp 1649977179
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_189
timestamp 1649977179
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_195
timestamp 1649977179
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1649977179
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1649977179
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1649977179
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1649977179
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1649977179
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1649977179
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1649977179
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1649977179
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1649977179
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1649977179
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1649977179
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1649977179
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1649977179
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1649977179
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1649977179
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_369
timestamp 1649977179
transform 1 0 35052 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_379
timestamp 1649977179
transform 1 0 35972 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_386
timestamp 1649977179
transform 1 0 36616 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_390
timestamp 1649977179
transform 1 0 36984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_395
timestamp 1649977179
transform 1 0 37444 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_403
timestamp 1649977179
transform 1 0 38180 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1649977179
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1649977179
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1649977179
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1649977179
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1649977179
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1649977179
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1649977179
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1649977179
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1649977179
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1649977179
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1649977179
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_137
timestamp 1649977179
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_149
timestamp 1649977179
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_161
timestamp 1649977179
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_167
timestamp 1649977179
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_169
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1649977179
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1649977179
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1649977179
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1649977179
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1649977179
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1649977179
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1649977179
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1649977179
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1649977179
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1649977179
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1649977179
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1649977179
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1649977179
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1649977179
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1649977179
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1649977179
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_361
timestamp 1649977179
transform 1 0 34316 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_367
timestamp 1649977179
transform 1 0 34868 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_370
timestamp 1649977179
transform 1 0 35144 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_378
timestamp 1649977179
transform 1 0 35880 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_381
timestamp 1649977179
transform 1 0 36156 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_388
timestamp 1649977179
transform 1 0 36800 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_401
timestamp 1649977179
transform 1 0 37996 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1649977179
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1649977179
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1649977179
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1649977179
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1649977179
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1649977179
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1649977179
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1649977179
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1649977179
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1649977179
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1649977179
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1649977179
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_153
timestamp 1649977179
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_165
timestamp 1649977179
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_177
timestamp 1649977179
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_189
timestamp 1649977179
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1649977179
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1649977179
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1649977179
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1649977179
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1649977179
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1649977179
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1649977179
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1649977179
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1649977179
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1649977179
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1649977179
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1649977179
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1649977179
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1649977179
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1649977179
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1649977179
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_365
timestamp 1649977179
transform 1 0 34684 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_371
timestamp 1649977179
transform 1 0 35236 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_374
timestamp 1649977179
transform 1 0 35512 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_387
timestamp 1649977179
transform 1 0 36708 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_400
timestamp 1649977179
transform 1 0 37904 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_406
timestamp 1649977179
transform 1 0 38456 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1649977179
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1649977179
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1649977179
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1649977179
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1649977179
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1649977179
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1649977179
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1649977179
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1649977179
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1649977179
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1649977179
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1649977179
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1649977179
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1649977179
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1649977179
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1649977179
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_169
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_181
timestamp 1649977179
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_193
timestamp 1649977179
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_205
timestamp 1649977179
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_217
timestamp 1649977179
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_223
timestamp 1649977179
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1649977179
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1649977179
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1649977179
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1649977179
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1649977179
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1649977179
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1649977179
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1649977179
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1649977179
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1649977179
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1649977179
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1649977179
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1649977179
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_361
timestamp 1649977179
transform 1 0 34316 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_59_369
timestamp 1649977179
transform 1 0 35052 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_374
timestamp 1649977179
transform 1 0 35512 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_381
timestamp 1649977179
transform 1 0 36156 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_388
timestamp 1649977179
transform 1 0 36800 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_59_393
timestamp 1649977179
transform 1 0 37260 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_403
timestamp 1649977179
transform 1 0 38180 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1649977179
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1649977179
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1649977179
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1649977179
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1649977179
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1649977179
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1649977179
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1649977179
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1649977179
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1649977179
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1649977179
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1649977179
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1649977179
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_153
timestamp 1649977179
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_165
timestamp 1649977179
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_177
timestamp 1649977179
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_189
timestamp 1649977179
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_195
timestamp 1649977179
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1649977179
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1649977179
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1649977179
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1649977179
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1649977179
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1649977179
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1649977179
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1649977179
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1649977179
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1649977179
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1649977179
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1649977179
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1649977179
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1649977179
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1649977179
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_365
timestamp 1649977179
transform 1 0 34684 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_373
timestamp 1649977179
transform 1 0 35420 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_378
timestamp 1649977179
transform 1 0 35880 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_384
timestamp 1649977179
transform 1 0 36432 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_392
timestamp 1649977179
transform 1 0 37168 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_401
timestamp 1649977179
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1649977179
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1649977179
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1649977179
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1649977179
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1649977179
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1649977179
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_57
timestamp 1649977179
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_69
timestamp 1649977179
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_61_81
timestamp 1649977179
transform 1 0 8556 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_61_86
timestamp 1649977179
transform 1 0 9016 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_98
timestamp 1649977179
transform 1 0 10120 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1649977179
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1649977179
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1649977179
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1649977179
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1649977179
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1649977179
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1649977179
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1649977179
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1649977179
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1649977179
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1649977179
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1649977179
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1649977179
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1649977179
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1649977179
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1649977179
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1649977179
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1649977179
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1649977179
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1649977179
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1649977179
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1649977179
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1649977179
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1649977179
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_361
timestamp 1649977179
transform 1 0 34316 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_367
timestamp 1649977179
transform 1 0 34868 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_370
timestamp 1649977179
transform 1 0 35144 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_376
timestamp 1649977179
transform 1 0 35696 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_382
timestamp 1649977179
transform 1 0 36248 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_388
timestamp 1649977179
transform 1 0 36800 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_395
timestamp 1649977179
transform 1 0 37444 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_403
timestamp 1649977179
transform 1 0 38180 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1649977179
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1649977179
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1649977179
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_29
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_35
timestamp 1649977179
transform 1 0 4324 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_38
timestamp 1649977179
transform 1 0 4600 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_44
timestamp 1649977179
transform 1 0 5152 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_50
timestamp 1649977179
transform 1 0 5704 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_64
timestamp 1649977179
transform 1 0 6992 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_70
timestamp 1649977179
transform 1 0 7544 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_78
timestamp 1649977179
transform 1 0 8280 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_96
timestamp 1649977179
transform 1 0 9936 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_102
timestamp 1649977179
transform 1 0 10488 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_110
timestamp 1649977179
transform 1 0 11224 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_113
timestamp 1649977179
transform 1 0 11500 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_119
timestamp 1649977179
transform 1 0 12052 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_62_127
timestamp 1649977179
transform 1 0 12788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1649977179
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1649977179
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1649977179
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1649977179
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1649977179
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1649977179
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1649977179
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1649977179
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1649977179
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1649977179
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1649977179
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1649977179
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1649977179
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1649977179
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1649977179
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1649977179
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1649977179
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1649977179
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1649977179
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1649977179
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1649977179
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1649977179
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1649977179
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_367
timestamp 1649977179
transform 1 0 34868 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_373
timestamp 1649977179
transform 1 0 35420 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_380
timestamp 1649977179
transform 1 0 36064 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_403
timestamp 1649977179
transform 1 0 38180 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_15
timestamp 1649977179
transform 1 0 2484 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_18
timestamp 1649977179
transform 1 0 2760 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_32
timestamp 1649977179
transform 1 0 4048 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_48
timestamp 1649977179
transform 1 0 5520 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_57
timestamp 1649977179
transform 1 0 6348 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_61
timestamp 1649977179
transform 1 0 6716 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_63_72
timestamp 1649977179
transform 1 0 7728 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_88
timestamp 1649977179
transform 1 0 9200 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_104
timestamp 1649977179
transform 1 0 10672 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_123
timestamp 1649977179
transform 1 0 12420 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_130
timestamp 1649977179
transform 1 0 13064 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_138
timestamp 1649977179
transform 1 0 13800 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_145
timestamp 1649977179
transform 1 0 14444 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_149
timestamp 1649977179
transform 1 0 14812 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_152
timestamp 1649977179
transform 1 0 15088 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_158
timestamp 1649977179
transform 1 0 15640 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_164
timestamp 1649977179
transform 1 0 16192 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_63_169
timestamp 1649977179
transform 1 0 16652 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_63_174
timestamp 1649977179
transform 1 0 17112 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_182
timestamp 1649977179
transform 1 0 17848 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_192
timestamp 1649977179
transform 1 0 18768 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_198
timestamp 1649977179
transform 1 0 19320 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_63_206
timestamp 1649977179
transform 1 0 20056 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_214
timestamp 1649977179
transform 1 0 20792 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1649977179
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_63_228
timestamp 1649977179
transform 1 0 22080 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_234
timestamp 1649977179
transform 1 0 22632 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_246
timestamp 1649977179
transform 1 0 23736 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_250
timestamp 1649977179
transform 1 0 24104 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_253
timestamp 1649977179
transform 1 0 24380 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_257
timestamp 1649977179
transform 1 0 24748 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_260
timestamp 1649977179
transform 1 0 25024 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_266
timestamp 1649977179
transform 1 0 25576 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1649977179
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1649977179
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_283
timestamp 1649977179
transform 1 0 27140 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_289
timestamp 1649977179
transform 1 0 27692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_301
timestamp 1649977179
transform 1 0 28796 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_309
timestamp 1649977179
transform 1 0 29532 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_313
timestamp 1649977179
transform 1 0 29900 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_316
timestamp 1649977179
transform 1 0 30176 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_322
timestamp 1649977179
transform 1 0 30728 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1649977179
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1649977179
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_339
timestamp 1649977179
transform 1 0 32292 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_63_345
timestamp 1649977179
transform 1 0 32844 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_357
timestamp 1649977179
transform 1 0 33948 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_361
timestamp 1649977179
transform 1 0 34316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_364
timestamp 1649977179
transform 1 0 34592 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_371
timestamp 1649977179
transform 1 0 35236 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_378
timestamp 1649977179
transform 1 0 35880 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1649977179
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1649977179
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_395
timestamp 1649977179
transform 1 0 37444 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_403
timestamp 1649977179
transform 1 0 38180 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_3
timestamp 1649977179
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_7
timestamp 1649977179
transform 1 0 1748 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_10
timestamp 1649977179
transform 1 0 2024 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_24
timestamp 1649977179
transform 1 0 3312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_29
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_64_34
timestamp 1649977179
transform 1 0 4232 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_52
timestamp 1649977179
transform 1 0 5888 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_59
timestamp 1649977179
transform 1 0 6532 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_63
timestamp 1649977179
transform 1 0 6900 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_66
timestamp 1649977179
transform 1 0 7176 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_80
timestamp 1649977179
transform 1 0 8464 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_91
timestamp 1649977179
transform 1 0 9476 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_94
timestamp 1649977179
transform 1 0 9752 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_108
timestamp 1649977179
transform 1 0 11040 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_113
timestamp 1649977179
transform 1 0 11500 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_117
timestamp 1649977179
transform 1 0 11868 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_128
timestamp 1649977179
transform 1 0 12880 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_132
timestamp 1649977179
transform 1 0 13248 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_136
timestamp 1649977179
transform 1 0 13616 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_143
timestamp 1649977179
transform 1 0 14260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_150
timestamp 1649977179
transform 1 0 14904 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_157
timestamp 1649977179
transform 1 0 15548 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_164
timestamp 1649977179
transform 1 0 16192 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_169
timestamp 1649977179
transform 1 0 16652 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_173
timestamp 1649977179
transform 1 0 17020 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_177
timestamp 1649977179
transform 1 0 17388 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_181
timestamp 1649977179
transform 1 0 17756 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_185
timestamp 1649977179
transform 1 0 18124 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_192
timestamp 1649977179
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_197
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_201
timestamp 1649977179
transform 1 0 19596 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_205
timestamp 1649977179
transform 1 0 19964 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_209
timestamp 1649977179
transform 1 0 20332 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_213
timestamp 1649977179
transform 1 0 20700 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_217
timestamp 1649977179
transform 1 0 21068 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_223
timestamp 1649977179
transform 1 0 21620 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_225
timestamp 1649977179
transform 1 0 21804 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_229
timestamp 1649977179
transform 1 0 22172 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_234
timestamp 1649977179
transform 1 0 22632 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_241
timestamp 1649977179
transform 1 0 23276 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_247
timestamp 1649977179
transform 1 0 23828 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_251
timestamp 1649977179
transform 1 0 24196 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_256
timestamp 1649977179
transform 1 0 24656 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_263
timestamp 1649977179
transform 1 0 25300 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_270
timestamp 1649977179
transform 1 0 25944 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_276
timestamp 1649977179
transform 1 0 26496 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_284
timestamp 1649977179
transform 1 0 27232 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_291
timestamp 1649977179
transform 1 0 27876 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_298
timestamp 1649977179
transform 1 0 28520 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_304
timestamp 1649977179
transform 1 0 29072 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_312
timestamp 1649977179
transform 1 0 29808 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_319
timestamp 1649977179
transform 1 0 30452 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_326
timestamp 1649977179
transform 1 0 31096 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_332
timestamp 1649977179
transform 1 0 31648 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_340
timestamp 1649977179
transform 1 0 32384 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_347
timestamp 1649977179
transform 1 0 33028 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_354
timestamp 1649977179
transform 1 0 33672 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_360
timestamp 1649977179
transform 1 0 34224 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_368
timestamp 1649977179
transform 1 0 34960 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_375
timestamp 1649977179
transform 1 0 35604 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_382
timestamp 1649977179
transform 1 0 36248 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_388
timestamp 1649977179
transform 1 0 36800 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_395
timestamp 1649977179
transform 1 0 37444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_403
timestamp 1649977179
transform 1 0 38180 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_4  _060_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 28060 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _061_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12512 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _062_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12696 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _063_
timestamp 1649977179
transform -1 0 12328 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _064_
timestamp 1649977179
transform 1 0 12512 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _065_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21896 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _066_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22264 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _067_
timestamp 1649977179
transform -1 0 12604 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _068_
timestamp 1649977179
transform 1 0 12052 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _069_
timestamp 1649977179
transform -1 0 35236 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1649977179
transform -1 0 35880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _071_
timestamp 1649977179
transform -1 0 35972 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1649977179
transform -1 0 36616 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _073_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20516 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _074_
timestamp 1649977179
transform -1 0 36800 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1649977179
transform 1 0 36800 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _076_
timestamp 1649977179
transform -1 0 8372 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _077_
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _078_
timestamp 1649977179
transform -1 0 8464 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _079_
timestamp 1649977179
transform 1 0 8832 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _080_
timestamp 1649977179
transform -1 0 8372 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _081_
timestamp 1649977179
transform 1 0 10212 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _082_
timestamp 1649977179
transform -1 0 8464 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _083_
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _084_
timestamp 1649977179
transform -1 0 8648 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _085_
timestamp 1649977179
transform 1 0 9108 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _086_
timestamp 1649977179
transform -1 0 8464 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _087_
timestamp 1649977179
transform 1 0 9476 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _088_
timestamp 1649977179
transform -1 0 9660 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _089_
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _090_
timestamp 1649977179
transform -1 0 9752 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _091_
timestamp 1649977179
transform 1 0 10120 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _092_
timestamp 1649977179
transform -1 0 10856 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _093_
timestamp 1649977179
transform 1 0 11224 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _094_
timestamp 1649977179
transform -1 0 19780 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _095_
timestamp 1649977179
transform -1 0 13248 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1649977179
transform -1 0 14352 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _097_
timestamp 1649977179
transform -1 0 13432 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1649977179
transform -1 0 14076 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _099_
timestamp 1649977179
transform -1 0 13432 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1649977179
transform -1 0 14352 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _101_
timestamp 1649977179
transform -1 0 13984 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1649977179
transform -1 0 14628 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _103_
timestamp 1649977179
transform -1 0 14904 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1649977179
transform -1 0 15548 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _105_
timestamp 1649977179
transform -1 0 15456 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1649977179
transform -1 0 16100 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _107_
timestamp 1649977179
transform -1 0 16192 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1649977179
transform -1 0 16928 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _109_
timestamp 1649977179
transform -1 0 16836 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1649977179
transform -1 0 17480 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _111_
timestamp 1649977179
transform -1 0 17572 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1649977179
transform -1 0 18216 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _113_
timestamp 1649977179
transform -1 0 18400 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1649977179
transform -1 0 18400 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _115_
timestamp 1649977179
transform 1 0 22908 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _116_
timestamp 1649977179
transform -1 0 18676 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1649977179
transform -1 0 19596 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _118_
timestamp 1649977179
transform -1 0 19872 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1649977179
transform -1 0 20516 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _120_
timestamp 1649977179
transform -1 0 20516 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1649977179
transform -1 0 21160 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _122_
timestamp 1649977179
transform -1 0 21252 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1649977179
transform -1 0 21344 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _124_
timestamp 1649977179
transform 1 0 21804 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1649977179
transform -1 0 22080 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _126_
timestamp 1649977179
transform -1 0 23460 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _127_
timestamp 1649977179
transform -1 0 24104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _128_
timestamp 1649977179
transform -1 0 24196 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1649977179
transform -1 0 24840 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _130_
timestamp 1649977179
transform -1 0 25208 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1649977179
transform -1 0 25852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _132_
timestamp 1649977179
transform -1 0 25668 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1649977179
transform -1 0 26312 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _134_
timestamp 1649977179
transform -1 0 26220 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 1649977179
transform -1 0 26864 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _136_
timestamp 1649977179
transform 1 0 30452 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _137_
timestamp 1649977179
transform -1 0 27784 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1649977179
transform -1 0 28612 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _139_
timestamp 1649977179
transform -1 0 27968 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp 1649977179
transform -1 0 28428 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _141_
timestamp 1649977179
transform -1 0 28612 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _142_
timestamp 1649977179
transform -1 0 29072 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _143_
timestamp 1649977179
transform -1 0 29348 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _144_
timestamp 1649977179
transform -1 0 29992 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _145_
timestamp 1649977179
transform -1 0 30084 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp 1649977179
transform -1 0 30176 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _147_
timestamp 1649977179
transform -1 0 30820 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 1649977179
transform -1 0 31464 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _149_
timestamp 1649977179
transform -1 0 31556 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _150_
timestamp 1649977179
transform -1 0 32384 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _151_
timestamp 1649977179
transform -1 0 32384 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _152_
timestamp 1649977179
transform -1 0 33028 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _153_
timestamp 1649977179
transform -1 0 33028 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1649977179
transform -1 0 33672 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _155_
timestamp 1649977179
transform -1 0 33580 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _156_
timestamp 1649977179
transform -1 0 34316 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _157_
timestamp 1649977179
transform -1 0 34224 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1649977179
transform -1 0 34960 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _159_
timestamp 1649977179
transform -1 0 36708 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1649977179
transform -1 0 36800 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _161_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 36524 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _162_
timestamp 1649977179
transform -1 0 37904 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _163_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 37996 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _164_
timestamp 1649977179
transform -1 0 36156 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _165_
timestamp 1649977179
transform 1 0 22816 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1649977179
transform 1 0 23000 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _167_
timestamp 1649977179
transform 1 0 12696 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _168_
timestamp 1649977179
transform 1 0 13524 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _169_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 37260 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _170_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 37444 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__dfxtp_4  _171_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 38180 0 1 35904
box -38 -48 1786 592
use sky130_fd_sc_hd__clkbuf_1  input1
timestamp 1649977179
transform -1 0 36064 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2
timestamp 1649977179
transform -1 0 35236 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input3 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 37720 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1649977179
transform -1 0 38180 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform 1 0 37904 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input6
timestamp 1649977179
transform 1 0 2392 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 1649977179
transform 1 0 3128 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 1649977179
transform 1 0 4600 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1649977179
transform 1 0 11960 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1649977179
transform -1 0 13064 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1649977179
transform -1 0 13616 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1649977179
transform -1 0 14444 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1649977179
transform -1 0 14904 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1649977179
transform -1 0 15548 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1649977179
transform -1 0 16192 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1649977179
transform -1 0 17388 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1649977179
transform -1 0 18124 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1649977179
transform 1 0 18492 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input19
timestamp 1649977179
transform -1 0 5888 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1649977179
transform -1 0 19596 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1649977179
transform -1 0 20332 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1649977179
transform -1 0 21068 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1649977179
transform -1 0 22080 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input24
timestamp 1649977179
transform 1 0 6072 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1649977179
transform 1 0 6808 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1649977179
transform 1 0 7544 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input27
timestamp 1649977179
transform 1 0 8280 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1649977179
transform 1 0 9016 0 1 35904
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1649977179
transform 1 0 9752 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 1649977179
transform 1 0 10120 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input31
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1649977179
transform 1 0 23000 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1649977179
transform 1 0 30820 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1649977179
transform 1 0 31096 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1649977179
transform 1 0 32108 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1649977179
transform 1 0 32752 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1649977179
transform 1 0 33396 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1649977179
transform 1 0 34684 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1649977179
transform 1 0 24380 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1649977179
transform 1 0 25024 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1649977179
transform 1 0 25668 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1649977179
transform 1 0 25944 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1649977179
transform -1 0 27232 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1649977179
transform 1 0 27600 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1649977179
transform 1 0 28244 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1649977179
transform 1 0 29532 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1649977179
transform 1 0 30176 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1649977179
transform 1 0 35328 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1649977179
transform 1 0 35972 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1649977179
transform 1 0 36248 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1649977179
transform -1 0 35880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1649977179
transform -1 0 2668 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1649977179
transform -1 0 3312 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1649977179
transform -1 0 4876 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1649977179
transform -1 0 12236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1649977179
transform -1 0 12972 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input57
timestamp 1649977179
transform -1 0 13616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input58
timestamp 1649977179
transform -1 0 14444 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input59
timestamp 1649977179
transform -1 0 14904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1649977179
transform -1 0 15548 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input61
timestamp 1649977179
transform -1 0 16192 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1649977179
transform -1 0 17388 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input63
timestamp 1649977179
transform -1 0 18124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input64
timestamp 1649977179
transform 1 0 18492 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input65
timestamp 1649977179
transform -1 0 5244 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input66
timestamp 1649977179
transform -1 0 19596 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input67
timestamp 1649977179
transform 1 0 20056 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input68
timestamp 1649977179
transform 1 0 20792 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input69
timestamp 1649977179
transform -1 0 22080 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input70
timestamp 1649977179
transform -1 0 5888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input71
timestamp 1649977179
transform -1 0 7084 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input72
timestamp 1649977179
transform -1 0 7820 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input73
timestamp 1649977179
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input74
timestamp 1649977179
transform -1 0 9292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input75
timestamp 1649977179
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input76
timestamp 1649977179
transform -1 0 10396 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input77
timestamp 1649977179
transform -1 0 11040 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input78
timestamp 1649977179
transform -1 0 23276 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input79
timestamp 1649977179
transform 1 0 30360 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input80
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input81
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input82
timestamp 1649977179
transform 1 0 33396 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input83
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input84
timestamp 1649977179
transform 1 0 34684 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1649977179
transform -1 0 24656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1649977179
transform -1 0 25300 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1649977179
transform -1 0 25944 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1649977179
transform -1 0 26220 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1649977179
transform -1 0 27232 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1649977179
transform -1 0 27876 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1649977179
transform -1 0 28520 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input92
timestamp 1649977179
transform -1 0 29164 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input93
timestamp 1649977179
transform -1 0 30544 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input94
timestamp 1649977179
transform 1 0 34776 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input95
timestamp 1649977179
transform 1 0 37260 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input96
timestamp 1649977179
transform 1 0 36248 0 1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input97
timestamp 1649977179
transform 1 0 36524 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output98 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 37812 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1649977179
transform 1 0 37812 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1649977179
transform 1 0 36432 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1649977179
transform 1 0 37812 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1649977179
transform 1 0 37812 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1649977179
transform 1 0 37812 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1649977179
transform 1 0 37812 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1649977179
transform 1 0 37812 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1649977179
transform 1 0 37812 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1649977179
transform 1 0 37812 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1649977179
transform 1 0 37812 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1649977179
transform 1 0 37812 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1649977179
transform 1 0 37812 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1649977179
transform 1 0 37812 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1649977179
transform 1 0 37812 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1649977179
transform 1 0 37812 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1649977179
transform 1 0 37812 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output115
timestamp 1649977179
transform 1 0 37812 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1649977179
transform 1 0 37812 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output117
timestamp 1649977179
transform 1 0 37812 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output118
timestamp 1649977179
transform 1 0 37812 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1649977179
transform 1 0 37812 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1649977179
transform 1 0 37812 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output121
timestamp 1649977179
transform 1 0 37812 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1649977179
transform 1 0 37812 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1649977179
transform 1 0 37812 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1649977179
transform 1 0 37812 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1649977179
transform 1 0 37812 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1649977179
transform 1 0 37812 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1649977179
transform 1 0 37812 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1649977179
transform 1 0 37812 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1649977179
transform 1 0 37812 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output130
timestamp 1649977179
transform 1 0 37812 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1649977179
transform 1 0 37812 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output132
timestamp 1649977179
transform 1 0 37812 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1649977179
transform 1 0 37812 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1649977179
transform 1 0 37812 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output135
timestamp 1649977179
transform 1 0 37812 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output136
timestamp 1649977179
transform 1 0 37812 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output137
timestamp 1649977179
transform 1 0 37812 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1649977179
transform 1 0 37812 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1649977179
transform 1 0 37812 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1649977179
transform 1 0 37812 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1649977179
transform 1 0 37812 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1649977179
transform 1 0 37812 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1649977179
transform 1 0 37076 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1649977179
transform 1 0 37812 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1649977179
transform 1 0 36800 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1649977179
transform -1 0 4232 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output147
timestamp 1649977179
transform 1 0 22264 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output148
timestamp 1649977179
transform -1 0 4232 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output149
timestamp 1649977179
transform -1 0 22632 0 1 2176
box -38 -48 406 592
<< labels >>
flabel metal3 s 39200 37272 40000 37392 0 FreeSans 480 0 0 0 i_clk
port 0 nsew signal input
flabel metal3 s 39200 36592 40000 36712 0 FreeSans 480 0 0 0 i_rst
port 1 nsew signal input
flabel metal2 s 37646 39200 37702 40000 0 FreeSans 224 90 0 0 i_wb0_cyc
port 2 nsew signal input
flabel metal2 s 37646 0 37702 800 0 FreeSans 224 90 0 0 i_wb1_cyc
port 3 nsew signal input
flabel metal3 s 39200 35912 40000 36032 0 FreeSans 480 0 0 0 o_sel_sig
port 4 nsew signal tristate
flabel metal3 s 39200 35232 40000 35352 0 FreeSans 480 0 0 0 o_wb_cyc
port 5 nsew signal tristate
flabel metal3 s 39200 2592 40000 2712 0 FreeSans 480 0 0 0 owb_4_burst
port 6 nsew signal tristate
flabel metal3 s 39200 3272 40000 3392 0 FreeSans 480 0 0 0 owb_8_burst
port 7 nsew signal tristate
flabel metal3 s 39200 3952 40000 4072 0 FreeSans 480 0 0 0 owb_ack
port 8 nsew signal input
flabel metal3 s 39200 4632 40000 4752 0 FreeSans 480 0 0 0 owb_adr[0]
port 9 nsew signal tristate
flabel metal3 s 39200 11432 40000 11552 0 FreeSans 480 0 0 0 owb_adr[10]
port 10 nsew signal tristate
flabel metal3 s 39200 12112 40000 12232 0 FreeSans 480 0 0 0 owb_adr[11]
port 11 nsew signal tristate
flabel metal3 s 39200 12792 40000 12912 0 FreeSans 480 0 0 0 owb_adr[12]
port 12 nsew signal tristate
flabel metal3 s 39200 13472 40000 13592 0 FreeSans 480 0 0 0 owb_adr[13]
port 13 nsew signal tristate
flabel metal3 s 39200 14152 40000 14272 0 FreeSans 480 0 0 0 owb_adr[14]
port 14 nsew signal tristate
flabel metal3 s 39200 14832 40000 14952 0 FreeSans 480 0 0 0 owb_adr[15]
port 15 nsew signal tristate
flabel metal3 s 39200 15512 40000 15632 0 FreeSans 480 0 0 0 owb_adr[16]
port 16 nsew signal tristate
flabel metal3 s 39200 16192 40000 16312 0 FreeSans 480 0 0 0 owb_adr[17]
port 17 nsew signal tristate
flabel metal3 s 39200 16872 40000 16992 0 FreeSans 480 0 0 0 owb_adr[18]
port 18 nsew signal tristate
flabel metal3 s 39200 17552 40000 17672 0 FreeSans 480 0 0 0 owb_adr[19]
port 19 nsew signal tristate
flabel metal3 s 39200 5312 40000 5432 0 FreeSans 480 0 0 0 owb_adr[1]
port 20 nsew signal tristate
flabel metal3 s 39200 18232 40000 18352 0 FreeSans 480 0 0 0 owb_adr[20]
port 21 nsew signal tristate
flabel metal3 s 39200 18912 40000 19032 0 FreeSans 480 0 0 0 owb_adr[21]
port 22 nsew signal tristate
flabel metal3 s 39200 19592 40000 19712 0 FreeSans 480 0 0 0 owb_adr[22]
port 23 nsew signal tristate
flabel metal3 s 39200 20272 40000 20392 0 FreeSans 480 0 0 0 owb_adr[23]
port 24 nsew signal tristate
flabel metal3 s 39200 5992 40000 6112 0 FreeSans 480 0 0 0 owb_adr[2]
port 25 nsew signal tristate
flabel metal3 s 39200 6672 40000 6792 0 FreeSans 480 0 0 0 owb_adr[3]
port 26 nsew signal tristate
flabel metal3 s 39200 7352 40000 7472 0 FreeSans 480 0 0 0 owb_adr[4]
port 27 nsew signal tristate
flabel metal3 s 39200 8032 40000 8152 0 FreeSans 480 0 0 0 owb_adr[5]
port 28 nsew signal tristate
flabel metal3 s 39200 8712 40000 8832 0 FreeSans 480 0 0 0 owb_adr[6]
port 29 nsew signal tristate
flabel metal3 s 39200 9392 40000 9512 0 FreeSans 480 0 0 0 owb_adr[7]
port 30 nsew signal tristate
flabel metal3 s 39200 10072 40000 10192 0 FreeSans 480 0 0 0 owb_adr[8]
port 31 nsew signal tristate
flabel metal3 s 39200 10752 40000 10872 0 FreeSans 480 0 0 0 owb_adr[9]
port 32 nsew signal tristate
flabel metal3 s 39200 20952 40000 21072 0 FreeSans 480 0 0 0 owb_err
port 33 nsew signal input
flabel metal3 s 39200 21632 40000 21752 0 FreeSans 480 0 0 0 owb_o_dat[0]
port 34 nsew signal tristate
flabel metal3 s 39200 28432 40000 28552 0 FreeSans 480 0 0 0 owb_o_dat[10]
port 35 nsew signal tristate
flabel metal3 s 39200 29112 40000 29232 0 FreeSans 480 0 0 0 owb_o_dat[11]
port 36 nsew signal tristate
flabel metal3 s 39200 29792 40000 29912 0 FreeSans 480 0 0 0 owb_o_dat[12]
port 37 nsew signal tristate
flabel metal3 s 39200 30472 40000 30592 0 FreeSans 480 0 0 0 owb_o_dat[13]
port 38 nsew signal tristate
flabel metal3 s 39200 31152 40000 31272 0 FreeSans 480 0 0 0 owb_o_dat[14]
port 39 nsew signal tristate
flabel metal3 s 39200 31832 40000 31952 0 FreeSans 480 0 0 0 owb_o_dat[15]
port 40 nsew signal tristate
flabel metal3 s 39200 22312 40000 22432 0 FreeSans 480 0 0 0 owb_o_dat[1]
port 41 nsew signal tristate
flabel metal3 s 39200 22992 40000 23112 0 FreeSans 480 0 0 0 owb_o_dat[2]
port 42 nsew signal tristate
flabel metal3 s 39200 23672 40000 23792 0 FreeSans 480 0 0 0 owb_o_dat[3]
port 43 nsew signal tristate
flabel metal3 s 39200 24352 40000 24472 0 FreeSans 480 0 0 0 owb_o_dat[4]
port 44 nsew signal tristate
flabel metal3 s 39200 25032 40000 25152 0 FreeSans 480 0 0 0 owb_o_dat[5]
port 45 nsew signal tristate
flabel metal3 s 39200 25712 40000 25832 0 FreeSans 480 0 0 0 owb_o_dat[6]
port 46 nsew signal tristate
flabel metal3 s 39200 26392 40000 26512 0 FreeSans 480 0 0 0 owb_o_dat[7]
port 47 nsew signal tristate
flabel metal3 s 39200 27072 40000 27192 0 FreeSans 480 0 0 0 owb_o_dat[8]
port 48 nsew signal tristate
flabel metal3 s 39200 27752 40000 27872 0 FreeSans 480 0 0 0 owb_o_dat[9]
port 49 nsew signal tristate
flabel metal3 s 39200 32512 40000 32632 0 FreeSans 480 0 0 0 owb_sel[0]
port 50 nsew signal tristate
flabel metal3 s 39200 33192 40000 33312 0 FreeSans 480 0 0 0 owb_sel[1]
port 51 nsew signal tristate
flabel metal3 s 39200 33872 40000 33992 0 FreeSans 480 0 0 0 owb_stb
port 52 nsew signal tristate
flabel metal3 s 39200 34552 40000 34672 0 FreeSans 480 0 0 0 owb_we
port 53 nsew signal tristate
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 54 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 54 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 55 nsew ground bidirectional
flabel metal2 s 2318 39200 2374 40000 0 FreeSans 224 90 0 0 wb0_4_burst
port 56 nsew signal input
flabel metal2 s 3054 39200 3110 40000 0 FreeSans 224 90 0 0 wb0_8_burst
port 57 nsew signal input
flabel metal2 s 3790 39200 3846 40000 0 FreeSans 224 90 0 0 wb0_ack
port 58 nsew signal tristate
flabel metal2 s 4526 39200 4582 40000 0 FreeSans 224 90 0 0 wb0_adr[0]
port 59 nsew signal input
flabel metal2 s 11886 39200 11942 40000 0 FreeSans 224 90 0 0 wb0_adr[10]
port 60 nsew signal input
flabel metal2 s 12622 39200 12678 40000 0 FreeSans 224 90 0 0 wb0_adr[11]
port 61 nsew signal input
flabel metal2 s 13358 39200 13414 40000 0 FreeSans 224 90 0 0 wb0_adr[12]
port 62 nsew signal input
flabel metal2 s 14094 39200 14150 40000 0 FreeSans 224 90 0 0 wb0_adr[13]
port 63 nsew signal input
flabel metal2 s 14830 39200 14886 40000 0 FreeSans 224 90 0 0 wb0_adr[14]
port 64 nsew signal input
flabel metal2 s 15566 39200 15622 40000 0 FreeSans 224 90 0 0 wb0_adr[15]
port 65 nsew signal input
flabel metal2 s 16302 39200 16358 40000 0 FreeSans 224 90 0 0 wb0_adr[16]
port 66 nsew signal input
flabel metal2 s 17038 39200 17094 40000 0 FreeSans 224 90 0 0 wb0_adr[17]
port 67 nsew signal input
flabel metal2 s 17774 39200 17830 40000 0 FreeSans 224 90 0 0 wb0_adr[18]
port 68 nsew signal input
flabel metal2 s 18510 39200 18566 40000 0 FreeSans 224 90 0 0 wb0_adr[19]
port 69 nsew signal input
flabel metal2 s 5262 39200 5318 40000 0 FreeSans 224 90 0 0 wb0_adr[1]
port 70 nsew signal input
flabel metal2 s 19246 39200 19302 40000 0 FreeSans 224 90 0 0 wb0_adr[20]
port 71 nsew signal input
flabel metal2 s 19982 39200 20038 40000 0 FreeSans 224 90 0 0 wb0_adr[21]
port 72 nsew signal input
flabel metal2 s 20718 39200 20774 40000 0 FreeSans 224 90 0 0 wb0_adr[22]
port 73 nsew signal input
flabel metal2 s 21454 39200 21510 40000 0 FreeSans 224 90 0 0 wb0_adr[23]
port 74 nsew signal input
flabel metal2 s 5998 39200 6054 40000 0 FreeSans 224 90 0 0 wb0_adr[2]
port 75 nsew signal input
flabel metal2 s 6734 39200 6790 40000 0 FreeSans 224 90 0 0 wb0_adr[3]
port 76 nsew signal input
flabel metal2 s 7470 39200 7526 40000 0 FreeSans 224 90 0 0 wb0_adr[4]
port 77 nsew signal input
flabel metal2 s 8206 39200 8262 40000 0 FreeSans 224 90 0 0 wb0_adr[5]
port 78 nsew signal input
flabel metal2 s 8942 39200 8998 40000 0 FreeSans 224 90 0 0 wb0_adr[6]
port 79 nsew signal input
flabel metal2 s 9678 39200 9734 40000 0 FreeSans 224 90 0 0 wb0_adr[7]
port 80 nsew signal input
flabel metal2 s 10414 39200 10470 40000 0 FreeSans 224 90 0 0 wb0_adr[8]
port 81 nsew signal input
flabel metal2 s 11150 39200 11206 40000 0 FreeSans 224 90 0 0 wb0_adr[9]
port 82 nsew signal input
flabel metal2 s 22190 39200 22246 40000 0 FreeSans 224 90 0 0 wb0_err
port 83 nsew signal tristate
flabel metal2 s 22926 39200 22982 40000 0 FreeSans 224 90 0 0 wb0_o_dat[0]
port 84 nsew signal input
flabel metal2 s 30286 39200 30342 40000 0 FreeSans 224 90 0 0 wb0_o_dat[10]
port 85 nsew signal input
flabel metal2 s 31022 39200 31078 40000 0 FreeSans 224 90 0 0 wb0_o_dat[11]
port 86 nsew signal input
flabel metal2 s 31758 39200 31814 40000 0 FreeSans 224 90 0 0 wb0_o_dat[12]
port 87 nsew signal input
flabel metal2 s 32494 39200 32550 40000 0 FreeSans 224 90 0 0 wb0_o_dat[13]
port 88 nsew signal input
flabel metal2 s 33230 39200 33286 40000 0 FreeSans 224 90 0 0 wb0_o_dat[14]
port 89 nsew signal input
flabel metal2 s 33966 39200 34022 40000 0 FreeSans 224 90 0 0 wb0_o_dat[15]
port 90 nsew signal input
flabel metal2 s 23662 39200 23718 40000 0 FreeSans 224 90 0 0 wb0_o_dat[1]
port 91 nsew signal input
flabel metal2 s 24398 39200 24454 40000 0 FreeSans 224 90 0 0 wb0_o_dat[2]
port 92 nsew signal input
flabel metal2 s 25134 39200 25190 40000 0 FreeSans 224 90 0 0 wb0_o_dat[3]
port 93 nsew signal input
flabel metal2 s 25870 39200 25926 40000 0 FreeSans 224 90 0 0 wb0_o_dat[4]
port 94 nsew signal input
flabel metal2 s 26606 39200 26662 40000 0 FreeSans 224 90 0 0 wb0_o_dat[5]
port 95 nsew signal input
flabel metal2 s 27342 39200 27398 40000 0 FreeSans 224 90 0 0 wb0_o_dat[6]
port 96 nsew signal input
flabel metal2 s 28078 39200 28134 40000 0 FreeSans 224 90 0 0 wb0_o_dat[7]
port 97 nsew signal input
flabel metal2 s 28814 39200 28870 40000 0 FreeSans 224 90 0 0 wb0_o_dat[8]
port 98 nsew signal input
flabel metal2 s 29550 39200 29606 40000 0 FreeSans 224 90 0 0 wb0_o_dat[9]
port 99 nsew signal input
flabel metal2 s 34702 39200 34758 40000 0 FreeSans 224 90 0 0 wb0_sel[0]
port 100 nsew signal input
flabel metal2 s 35438 39200 35494 40000 0 FreeSans 224 90 0 0 wb0_sel[1]
port 101 nsew signal input
flabel metal2 s 36174 39200 36230 40000 0 FreeSans 224 90 0 0 wb0_stb
port 102 nsew signal input
flabel metal2 s 36910 39200 36966 40000 0 FreeSans 224 90 0 0 wb0_we
port 103 nsew signal input
flabel metal2 s 2318 0 2374 800 0 FreeSans 224 90 0 0 wb1_4_burst
port 104 nsew signal input
flabel metal2 s 3054 0 3110 800 0 FreeSans 224 90 0 0 wb1_8_burst
port 105 nsew signal input
flabel metal2 s 3790 0 3846 800 0 FreeSans 224 90 0 0 wb1_ack
port 106 nsew signal tristate
flabel metal2 s 4526 0 4582 800 0 FreeSans 224 90 0 0 wb1_adr[0]
port 107 nsew signal input
flabel metal2 s 11886 0 11942 800 0 FreeSans 224 90 0 0 wb1_adr[10]
port 108 nsew signal input
flabel metal2 s 12622 0 12678 800 0 FreeSans 224 90 0 0 wb1_adr[11]
port 109 nsew signal input
flabel metal2 s 13358 0 13414 800 0 FreeSans 224 90 0 0 wb1_adr[12]
port 110 nsew signal input
flabel metal2 s 14094 0 14150 800 0 FreeSans 224 90 0 0 wb1_adr[13]
port 111 nsew signal input
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 wb1_adr[14]
port 112 nsew signal input
flabel metal2 s 15566 0 15622 800 0 FreeSans 224 90 0 0 wb1_adr[15]
port 113 nsew signal input
flabel metal2 s 16302 0 16358 800 0 FreeSans 224 90 0 0 wb1_adr[16]
port 114 nsew signal input
flabel metal2 s 17038 0 17094 800 0 FreeSans 224 90 0 0 wb1_adr[17]
port 115 nsew signal input
flabel metal2 s 17774 0 17830 800 0 FreeSans 224 90 0 0 wb1_adr[18]
port 116 nsew signal input
flabel metal2 s 18510 0 18566 800 0 FreeSans 224 90 0 0 wb1_adr[19]
port 117 nsew signal input
flabel metal2 s 5262 0 5318 800 0 FreeSans 224 90 0 0 wb1_adr[1]
port 118 nsew signal input
flabel metal2 s 19246 0 19302 800 0 FreeSans 224 90 0 0 wb1_adr[20]
port 119 nsew signal input
flabel metal2 s 19982 0 20038 800 0 FreeSans 224 90 0 0 wb1_adr[21]
port 120 nsew signal input
flabel metal2 s 20718 0 20774 800 0 FreeSans 224 90 0 0 wb1_adr[22]
port 121 nsew signal input
flabel metal2 s 21454 0 21510 800 0 FreeSans 224 90 0 0 wb1_adr[23]
port 122 nsew signal input
flabel metal2 s 5998 0 6054 800 0 FreeSans 224 90 0 0 wb1_adr[2]
port 123 nsew signal input
flabel metal2 s 6734 0 6790 800 0 FreeSans 224 90 0 0 wb1_adr[3]
port 124 nsew signal input
flabel metal2 s 7470 0 7526 800 0 FreeSans 224 90 0 0 wb1_adr[4]
port 125 nsew signal input
flabel metal2 s 8206 0 8262 800 0 FreeSans 224 90 0 0 wb1_adr[5]
port 126 nsew signal input
flabel metal2 s 8942 0 8998 800 0 FreeSans 224 90 0 0 wb1_adr[6]
port 127 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 wb1_adr[7]
port 128 nsew signal input
flabel metal2 s 10414 0 10470 800 0 FreeSans 224 90 0 0 wb1_adr[8]
port 129 nsew signal input
flabel metal2 s 11150 0 11206 800 0 FreeSans 224 90 0 0 wb1_adr[9]
port 130 nsew signal input
flabel metal2 s 22190 0 22246 800 0 FreeSans 224 90 0 0 wb1_err
port 131 nsew signal tristate
flabel metal2 s 22926 0 22982 800 0 FreeSans 224 90 0 0 wb1_o_dat[0]
port 132 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 wb1_o_dat[10]
port 133 nsew signal input
flabel metal2 s 31022 0 31078 800 0 FreeSans 224 90 0 0 wb1_o_dat[11]
port 134 nsew signal input
flabel metal2 s 31758 0 31814 800 0 FreeSans 224 90 0 0 wb1_o_dat[12]
port 135 nsew signal input
flabel metal2 s 32494 0 32550 800 0 FreeSans 224 90 0 0 wb1_o_dat[13]
port 136 nsew signal input
flabel metal2 s 33230 0 33286 800 0 FreeSans 224 90 0 0 wb1_o_dat[14]
port 137 nsew signal input
flabel metal2 s 33966 0 34022 800 0 FreeSans 224 90 0 0 wb1_o_dat[15]
port 138 nsew signal input
flabel metal2 s 23662 0 23718 800 0 FreeSans 224 90 0 0 wb1_o_dat[1]
port 139 nsew signal input
flabel metal2 s 24398 0 24454 800 0 FreeSans 224 90 0 0 wb1_o_dat[2]
port 140 nsew signal input
flabel metal2 s 25134 0 25190 800 0 FreeSans 224 90 0 0 wb1_o_dat[3]
port 141 nsew signal input
flabel metal2 s 25870 0 25926 800 0 FreeSans 224 90 0 0 wb1_o_dat[4]
port 142 nsew signal input
flabel metal2 s 26606 0 26662 800 0 FreeSans 224 90 0 0 wb1_o_dat[5]
port 143 nsew signal input
flabel metal2 s 27342 0 27398 800 0 FreeSans 224 90 0 0 wb1_o_dat[6]
port 144 nsew signal input
flabel metal2 s 28078 0 28134 800 0 FreeSans 224 90 0 0 wb1_o_dat[7]
port 145 nsew signal input
flabel metal2 s 28814 0 28870 800 0 FreeSans 224 90 0 0 wb1_o_dat[8]
port 146 nsew signal input
flabel metal2 s 29550 0 29606 800 0 FreeSans 224 90 0 0 wb1_o_dat[9]
port 147 nsew signal input
flabel metal2 s 34702 0 34758 800 0 FreeSans 224 90 0 0 wb1_sel[0]
port 148 nsew signal input
flabel metal2 s 35438 0 35494 800 0 FreeSans 224 90 0 0 wb1_sel[1]
port 149 nsew signal input
flabel metal2 s 36174 0 36230 800 0 FreeSans 224 90 0 0 wb1_stb
port 150 nsew signal input
flabel metal2 s 36910 0 36966 800 0 FreeSans 224 90 0 0 wb1_we
port 151 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
