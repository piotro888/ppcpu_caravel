magic
tech sky130B
magscale 1 2
timestamp 1662658114
<< obsli1 >>
rect 1104 2159 78844 77809
<< obsm1 >>
rect 14 1572 79290 78056
<< metal2 >>
rect 18 79200 74 80000
rect 1306 79200 1362 80000
rect 3238 79200 3294 80000
rect 4526 79200 4582 80000
rect 5814 79200 5870 80000
rect 7102 79200 7158 80000
rect 9034 79200 9090 80000
rect 10322 79200 10378 80000
rect 11610 79200 11666 80000
rect 12898 79200 12954 80000
rect 14830 79200 14886 80000
rect 16118 79200 16174 80000
rect 17406 79200 17462 80000
rect 18694 79200 18750 80000
rect 20626 79200 20682 80000
rect 21914 79200 21970 80000
rect 23202 79200 23258 80000
rect 24490 79200 24546 80000
rect 26422 79200 26478 80000
rect 27710 79200 27766 80000
rect 28998 79200 29054 80000
rect 30286 79200 30342 80000
rect 31574 79200 31630 80000
rect 33506 79200 33562 80000
rect 34794 79200 34850 80000
rect 36082 79200 36138 80000
rect 37370 79200 37426 80000
rect 39302 79200 39358 80000
rect 40590 79200 40646 80000
rect 41878 79200 41934 80000
rect 43166 79200 43222 80000
rect 45098 79200 45154 80000
rect 46386 79200 46442 80000
rect 47674 79200 47730 80000
rect 48962 79200 49018 80000
rect 50894 79200 50950 80000
rect 52182 79200 52238 80000
rect 53470 79200 53526 80000
rect 54758 79200 54814 80000
rect 56690 79200 56746 80000
rect 57978 79200 58034 80000
rect 59266 79200 59322 80000
rect 60554 79200 60610 80000
rect 62486 79200 62542 80000
rect 63774 79200 63830 80000
rect 65062 79200 65118 80000
rect 66350 79200 66406 80000
rect 67638 79200 67694 80000
rect 69570 79200 69626 80000
rect 70858 79200 70914 80000
rect 72146 79200 72202 80000
rect 73434 79200 73490 80000
rect 75366 79200 75422 80000
rect 76654 79200 76710 80000
rect 77942 79200 77998 80000
rect 79230 79200 79286 80000
rect 18 0 74 800
rect 1306 0 1362 800
rect 2594 0 2650 800
rect 3882 0 3938 800
rect 5170 0 5226 800
rect 7102 0 7158 800
rect 8390 0 8446 800
rect 9678 0 9734 800
rect 10966 0 11022 800
rect 12898 0 12954 800
rect 14186 0 14242 800
rect 15474 0 15530 800
rect 16762 0 16818 800
rect 18694 0 18750 800
rect 19982 0 20038 800
rect 21270 0 21326 800
rect 22558 0 22614 800
rect 24490 0 24546 800
rect 25778 0 25834 800
rect 27066 0 27122 800
rect 28354 0 28410 800
rect 30286 0 30342 800
rect 31574 0 31630 800
rect 32862 0 32918 800
rect 34150 0 34206 800
rect 35438 0 35494 800
rect 37370 0 37426 800
rect 38658 0 38714 800
rect 39946 0 40002 800
rect 41234 0 41290 800
rect 43166 0 43222 800
rect 44454 0 44510 800
rect 45742 0 45798 800
rect 47030 0 47086 800
rect 48962 0 49018 800
rect 50250 0 50306 800
rect 51538 0 51594 800
rect 52826 0 52882 800
rect 54758 0 54814 800
rect 56046 0 56102 800
rect 57334 0 57390 800
rect 58622 0 58678 800
rect 60554 0 60610 800
rect 61842 0 61898 800
rect 63130 0 63186 800
rect 64418 0 64474 800
rect 66350 0 66406 800
rect 67638 0 67694 800
rect 68926 0 68982 800
rect 70214 0 70270 800
rect 71502 0 71558 800
rect 73434 0 73490 800
rect 74722 0 74778 800
rect 76010 0 76066 800
rect 77298 0 77354 800
rect 79230 0 79286 800
<< obsm2 >>
rect 130 79144 1250 79234
rect 1418 79144 3182 79234
rect 3350 79144 4470 79234
rect 4638 79144 5758 79234
rect 5926 79144 7046 79234
rect 7214 79144 8978 79234
rect 9146 79144 10266 79234
rect 10434 79144 11554 79234
rect 11722 79144 12842 79234
rect 13010 79144 14774 79234
rect 14942 79144 16062 79234
rect 16230 79144 17350 79234
rect 17518 79144 18638 79234
rect 18806 79144 20570 79234
rect 20738 79144 21858 79234
rect 22026 79144 23146 79234
rect 23314 79144 24434 79234
rect 24602 79144 26366 79234
rect 26534 79144 27654 79234
rect 27822 79144 28942 79234
rect 29110 79144 30230 79234
rect 30398 79144 31518 79234
rect 31686 79144 33450 79234
rect 33618 79144 34738 79234
rect 34906 79144 36026 79234
rect 36194 79144 37314 79234
rect 37482 79144 39246 79234
rect 39414 79144 40534 79234
rect 40702 79144 41822 79234
rect 41990 79144 43110 79234
rect 43278 79144 45042 79234
rect 45210 79144 46330 79234
rect 46498 79144 47618 79234
rect 47786 79144 48906 79234
rect 49074 79144 50838 79234
rect 51006 79144 52126 79234
rect 52294 79144 53414 79234
rect 53582 79144 54702 79234
rect 54870 79144 56634 79234
rect 56802 79144 57922 79234
rect 58090 79144 59210 79234
rect 59378 79144 60498 79234
rect 60666 79144 62430 79234
rect 62598 79144 63718 79234
rect 63886 79144 65006 79234
rect 65174 79144 66294 79234
rect 66462 79144 67582 79234
rect 67750 79144 69514 79234
rect 69682 79144 70802 79234
rect 70970 79144 72090 79234
rect 72258 79144 73378 79234
rect 73546 79144 75310 79234
rect 75478 79144 76598 79234
rect 76766 79144 77886 79234
rect 78054 79144 79174 79234
rect 20 856 79284 79144
rect 130 31 1250 856
rect 1418 31 2538 856
rect 2706 31 3826 856
rect 3994 31 5114 856
rect 5282 31 7046 856
rect 7214 31 8334 856
rect 8502 31 9622 856
rect 9790 31 10910 856
rect 11078 31 12842 856
rect 13010 31 14130 856
rect 14298 31 15418 856
rect 15586 31 16706 856
rect 16874 31 18638 856
rect 18806 31 19926 856
rect 20094 31 21214 856
rect 21382 31 22502 856
rect 22670 31 24434 856
rect 24602 31 25722 856
rect 25890 31 27010 856
rect 27178 31 28298 856
rect 28466 31 30230 856
rect 30398 31 31518 856
rect 31686 31 32806 856
rect 32974 31 34094 856
rect 34262 31 35382 856
rect 35550 31 37314 856
rect 37482 31 38602 856
rect 38770 31 39890 856
rect 40058 31 41178 856
rect 41346 31 43110 856
rect 43278 31 44398 856
rect 44566 31 45686 856
rect 45854 31 46974 856
rect 47142 31 48906 856
rect 49074 31 50194 856
rect 50362 31 51482 856
rect 51650 31 52770 856
rect 52938 31 54702 856
rect 54870 31 55990 856
rect 56158 31 57278 856
rect 57446 31 58566 856
rect 58734 31 60498 856
rect 60666 31 61786 856
rect 61954 31 63074 856
rect 63242 31 64362 856
rect 64530 31 66294 856
rect 66462 31 67582 856
rect 67750 31 68870 856
rect 69038 31 70158 856
rect 70326 31 71446 856
rect 71614 31 73378 856
rect 73546 31 74666 856
rect 74834 31 75954 856
rect 76122 31 77242 856
rect 77410 31 79174 856
<< metal3 >>
rect 0 78888 800 79008
rect 79200 78888 80000 79008
rect 0 77528 800 77648
rect 79200 77528 80000 77648
rect 79200 76168 80000 76288
rect 0 75488 800 75608
rect 79200 74808 80000 74928
rect 0 74128 800 74248
rect 0 72768 800 72888
rect 79200 72768 80000 72888
rect 0 71408 800 71528
rect 79200 71408 80000 71528
rect 0 70048 800 70168
rect 79200 70048 80000 70168
rect 79200 68688 80000 68808
rect 0 68008 800 68128
rect 0 66648 800 66768
rect 79200 66648 80000 66768
rect 0 65288 800 65408
rect 79200 65288 80000 65408
rect 0 63928 800 64048
rect 79200 63928 80000 64048
rect 79200 62568 80000 62688
rect 0 61888 800 62008
rect 79200 61208 80000 61328
rect 0 60528 800 60648
rect 0 59168 800 59288
rect 79200 59168 80000 59288
rect 0 57808 800 57928
rect 79200 57808 80000 57928
rect 79200 56448 80000 56568
rect 0 55768 800 55888
rect 79200 55088 80000 55208
rect 0 54408 800 54528
rect 0 53048 800 53168
rect 79200 53048 80000 53168
rect 0 51688 800 51808
rect 79200 51688 80000 51808
rect 79200 50328 80000 50448
rect 0 49648 800 49768
rect 79200 48968 80000 49088
rect 0 48288 800 48408
rect 0 46928 800 47048
rect 79200 46928 80000 47048
rect 0 45568 800 45688
rect 79200 45568 80000 45688
rect 79200 44208 80000 44328
rect 0 43528 800 43648
rect 79200 42848 80000 42968
rect 0 42168 800 42288
rect 0 40808 800 40928
rect 79200 40808 80000 40928
rect 0 39448 800 39568
rect 79200 39448 80000 39568
rect 79200 38088 80000 38208
rect 0 37408 800 37528
rect 79200 36728 80000 36848
rect 0 36048 800 36168
rect 0 34688 800 34808
rect 79200 34688 80000 34808
rect 0 33328 800 33448
rect 79200 33328 80000 33448
rect 0 31968 800 32088
rect 79200 31968 80000 32088
rect 79200 30608 80000 30728
rect 0 29928 800 30048
rect 0 28568 800 28688
rect 79200 28568 80000 28688
rect 0 27208 800 27328
rect 79200 27208 80000 27328
rect 0 25848 800 25968
rect 79200 25848 80000 25968
rect 79200 24488 80000 24608
rect 0 23808 800 23928
rect 79200 23128 80000 23248
rect 0 22448 800 22568
rect 0 21088 800 21208
rect 79200 21088 80000 21208
rect 0 19728 800 19848
rect 79200 19728 80000 19848
rect 79200 18368 80000 18488
rect 0 17688 800 17808
rect 79200 17008 80000 17128
rect 0 16328 800 16448
rect 0 14968 800 15088
rect 79200 14968 80000 15088
rect 0 13608 800 13728
rect 79200 13608 80000 13728
rect 79200 12248 80000 12368
rect 0 11568 800 11688
rect 79200 10888 80000 11008
rect 0 10208 800 10328
rect 0 8848 800 8968
rect 79200 8848 80000 8968
rect 0 7488 800 7608
rect 79200 7488 80000 7608
rect 79200 6128 80000 6248
rect 0 5448 800 5568
rect 79200 4768 80000 4888
rect 0 4088 800 4208
rect 0 2728 800 2848
rect 79200 2728 80000 2848
rect 0 1368 800 1488
rect 79200 1368 80000 1488
rect 79200 8 80000 128
<< obsm3 >>
rect 880 78808 79120 78981
rect 800 77728 79200 78808
rect 880 77448 79120 77728
rect 800 76368 79200 77448
rect 800 76088 79120 76368
rect 800 75688 79200 76088
rect 880 75408 79200 75688
rect 800 75008 79200 75408
rect 800 74728 79120 75008
rect 800 74328 79200 74728
rect 880 74048 79200 74328
rect 800 72968 79200 74048
rect 880 72688 79120 72968
rect 800 71608 79200 72688
rect 880 71328 79120 71608
rect 800 70248 79200 71328
rect 880 69968 79120 70248
rect 800 68888 79200 69968
rect 800 68608 79120 68888
rect 800 68208 79200 68608
rect 880 67928 79200 68208
rect 800 66848 79200 67928
rect 880 66568 79120 66848
rect 800 65488 79200 66568
rect 880 65208 79120 65488
rect 800 64128 79200 65208
rect 880 63848 79120 64128
rect 800 62768 79200 63848
rect 800 62488 79120 62768
rect 800 62088 79200 62488
rect 880 61808 79200 62088
rect 800 61408 79200 61808
rect 800 61128 79120 61408
rect 800 60728 79200 61128
rect 880 60448 79200 60728
rect 800 59368 79200 60448
rect 880 59088 79120 59368
rect 800 58008 79200 59088
rect 880 57728 79120 58008
rect 800 56648 79200 57728
rect 800 56368 79120 56648
rect 800 55968 79200 56368
rect 880 55688 79200 55968
rect 800 55288 79200 55688
rect 800 55008 79120 55288
rect 800 54608 79200 55008
rect 880 54328 79200 54608
rect 800 53248 79200 54328
rect 880 52968 79120 53248
rect 800 51888 79200 52968
rect 880 51608 79120 51888
rect 800 50528 79200 51608
rect 800 50248 79120 50528
rect 800 49848 79200 50248
rect 880 49568 79200 49848
rect 800 49168 79200 49568
rect 800 48888 79120 49168
rect 800 48488 79200 48888
rect 880 48208 79200 48488
rect 800 47128 79200 48208
rect 880 46848 79120 47128
rect 800 45768 79200 46848
rect 880 45488 79120 45768
rect 800 44408 79200 45488
rect 800 44128 79120 44408
rect 800 43728 79200 44128
rect 880 43448 79200 43728
rect 800 43048 79200 43448
rect 800 42768 79120 43048
rect 800 42368 79200 42768
rect 880 42088 79200 42368
rect 800 41008 79200 42088
rect 880 40728 79120 41008
rect 800 39648 79200 40728
rect 880 39368 79120 39648
rect 800 38288 79200 39368
rect 800 38008 79120 38288
rect 800 37608 79200 38008
rect 880 37328 79200 37608
rect 800 36928 79200 37328
rect 800 36648 79120 36928
rect 800 36248 79200 36648
rect 880 35968 79200 36248
rect 800 34888 79200 35968
rect 880 34608 79120 34888
rect 800 33528 79200 34608
rect 880 33248 79120 33528
rect 800 32168 79200 33248
rect 880 31888 79120 32168
rect 800 30808 79200 31888
rect 800 30528 79120 30808
rect 800 30128 79200 30528
rect 880 29848 79200 30128
rect 800 28768 79200 29848
rect 880 28488 79120 28768
rect 800 27408 79200 28488
rect 880 27128 79120 27408
rect 800 26048 79200 27128
rect 880 25768 79120 26048
rect 800 24688 79200 25768
rect 800 24408 79120 24688
rect 800 24008 79200 24408
rect 880 23728 79200 24008
rect 800 23328 79200 23728
rect 800 23048 79120 23328
rect 800 22648 79200 23048
rect 880 22368 79200 22648
rect 800 21288 79200 22368
rect 880 21008 79120 21288
rect 800 19928 79200 21008
rect 880 19648 79120 19928
rect 800 18568 79200 19648
rect 800 18288 79120 18568
rect 800 17888 79200 18288
rect 880 17608 79200 17888
rect 800 17208 79200 17608
rect 800 16928 79120 17208
rect 800 16528 79200 16928
rect 880 16248 79200 16528
rect 800 15168 79200 16248
rect 880 14888 79120 15168
rect 800 13808 79200 14888
rect 880 13528 79120 13808
rect 800 12448 79200 13528
rect 800 12168 79120 12448
rect 800 11768 79200 12168
rect 880 11488 79200 11768
rect 800 11088 79200 11488
rect 800 10808 79120 11088
rect 800 10408 79200 10808
rect 880 10128 79200 10408
rect 800 9048 79200 10128
rect 880 8768 79120 9048
rect 800 7688 79200 8768
rect 880 7408 79120 7688
rect 800 6328 79200 7408
rect 800 6048 79120 6328
rect 800 5648 79200 6048
rect 880 5368 79200 5648
rect 800 4968 79200 5368
rect 800 4688 79120 4968
rect 800 4288 79200 4688
rect 880 4008 79200 4288
rect 800 2928 79200 4008
rect 880 2648 79120 2928
rect 800 1568 79200 2648
rect 880 1288 79120 1568
rect 800 208 79200 1288
rect 800 35 79120 208
<< metal4 >>
rect 4208 2128 4528 77840
rect 19568 2128 19888 77840
rect 34928 2128 35248 77840
rect 50288 2128 50608 77840
rect 65648 2128 65968 77840
<< obsm4 >>
rect 23243 2619 34848 77485
rect 35328 2619 50208 77485
rect 50688 2619 65568 77485
rect 66048 2619 67285 77485
<< labels >>
rlabel metal2 s 66350 0 66406 800 6 c_alu_carry_en
port 1 nsew signal input
rlabel metal2 s 40590 79200 40646 80000 6 c_alu_flags_ie
port 2 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 c_alu_mode[0]
port 3 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 c_alu_mode[1]
port 4 nsew signal input
rlabel metal2 s 60554 79200 60610 80000 6 c_alu_mode[2]
port 5 nsew signal input
rlabel metal2 s 44454 0 44510 800 6 c_alu_mode[3]
port 6 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 c_jump_cond_code[0]
port 7 nsew signal input
rlabel metal2 s 45098 79200 45154 80000 6 c_jump_cond_code[1]
port 8 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 c_jump_cond_code[2]
port 9 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 c_jump_cond_code[3]
port 10 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 c_jump_cond_code[4]
port 11 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 c_l_reg_sel[0]
port 12 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 c_l_reg_sel[1]
port 13 nsew signal input
rlabel metal3 s 79200 2728 80000 2848 6 c_l_reg_sel[2]
port 14 nsew signal input
rlabel metal3 s 79200 77528 80000 77648 6 c_mem_access
port 15 nsew signal input
rlabel metal2 s 77942 79200 77998 80000 6 c_mem_we
port 16 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 c_mem_width
port 17 nsew signal input
rlabel metal3 s 79200 12248 80000 12368 6 c_pc_ie
port 18 nsew signal input
rlabel metal3 s 79200 6128 80000 6248 6 c_pc_inc
port 19 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 c_r_bus_imm
port 20 nsew signal input
rlabel metal3 s 79200 24488 80000 24608 6 c_r_reg_sel[0]
port 21 nsew signal input
rlabel metal2 s 23202 79200 23258 80000 6 c_r_reg_sel[1]
port 22 nsew signal input
rlabel metal3 s 79200 72768 80000 72888 6 c_r_reg_sel[2]
port 23 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 c_rf_ie[0]
port 24 nsew signal input
rlabel metal2 s 61842 0 61898 800 6 c_rf_ie[1]
port 25 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 c_rf_ie[2]
port 26 nsew signal input
rlabel metal2 s 16118 79200 16174 80000 6 c_rf_ie[3]
port 27 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 c_rf_ie[4]
port 28 nsew signal input
rlabel metal3 s 79200 30608 80000 30728 6 c_rf_ie[5]
port 29 nsew signal input
rlabel metal2 s 9034 79200 9090 80000 6 c_rf_ie[6]
port 30 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 c_rf_ie[7]
port 31 nsew signal input
rlabel metal3 s 79200 44208 80000 44328 6 c_sreg_irt
port 32 nsew signal input
rlabel metal3 s 79200 48968 80000 49088 6 c_sreg_jal_over
port 33 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 c_sreg_load
port 34 nsew signal input
rlabel metal2 s 37370 79200 37426 80000 6 c_sreg_store
port 35 nsew signal input
rlabel metal2 s 77298 0 77354 800 6 c_sys
port 36 nsew signal input
rlabel metal2 s 69570 79200 69626 80000 6 c_used_operands[0]
port 37 nsew signal input
rlabel metal2 s 4526 79200 4582 80000 6 c_used_operands[1]
port 38 nsew signal input
rlabel metal2 s 27710 79200 27766 80000 6 dbg_pc[0]
port 39 nsew signal output
rlabel metal3 s 0 77528 800 77648 6 dbg_pc[10]
port 40 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 dbg_pc[11]
port 41 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 dbg_pc[12]
port 42 nsew signal output
rlabel metal2 s 38658 0 38714 800 6 dbg_pc[13]
port 43 nsew signal output
rlabel metal2 s 14830 79200 14886 80000 6 dbg_pc[14]
port 44 nsew signal output
rlabel metal2 s 79230 0 79286 800 6 dbg_pc[15]
port 45 nsew signal output
rlabel metal3 s 79200 28568 80000 28688 6 dbg_pc[1]
port 46 nsew signal output
rlabel metal2 s 70858 79200 70914 80000 6 dbg_pc[2]
port 47 nsew signal output
rlabel metal3 s 79200 51688 80000 51808 6 dbg_pc[3]
port 48 nsew signal output
rlabel metal3 s 0 70048 800 70168 6 dbg_pc[4]
port 49 nsew signal output
rlabel metal2 s 25778 0 25834 800 6 dbg_pc[5]
port 50 nsew signal output
rlabel metal2 s 67638 79200 67694 80000 6 dbg_pc[6]
port 51 nsew signal output
rlabel metal2 s 1306 79200 1362 80000 6 dbg_pc[7]
port 52 nsew signal output
rlabel metal2 s 24490 0 24546 800 6 dbg_pc[8]
port 53 nsew signal output
rlabel metal2 s 24490 79200 24546 80000 6 dbg_pc[9]
port 54 nsew signal output
rlabel metal3 s 79200 74808 80000 74928 6 dbg_r0[0]
port 55 nsew signal output
rlabel metal3 s 0 48288 800 48408 6 dbg_r0[10]
port 56 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 dbg_r0[11]
port 57 nsew signal output
rlabel metal3 s 79200 46928 80000 47048 6 dbg_r0[12]
port 58 nsew signal output
rlabel metal3 s 79200 36728 80000 36848 6 dbg_r0[13]
port 59 nsew signal output
rlabel metal3 s 0 72768 800 72888 6 dbg_r0[14]
port 60 nsew signal output
rlabel metal3 s 79200 25848 80000 25968 6 dbg_r0[15]
port 61 nsew signal output
rlabel metal3 s 0 22448 800 22568 6 dbg_r0[1]
port 62 nsew signal output
rlabel metal3 s 79200 66648 80000 66768 6 dbg_r0[2]
port 63 nsew signal output
rlabel metal2 s 57978 79200 58034 80000 6 dbg_r0[3]
port 64 nsew signal output
rlabel metal3 s 0 60528 800 60648 6 dbg_r0[4]
port 65 nsew signal output
rlabel metal2 s 59266 79200 59322 80000 6 dbg_r0[5]
port 66 nsew signal output
rlabel metal3 s 0 23808 800 23928 6 dbg_r0[6]
port 67 nsew signal output
rlabel metal2 s 48962 79200 49018 80000 6 dbg_r0[7]
port 68 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 dbg_r0[8]
port 69 nsew signal output
rlabel metal3 s 0 1368 800 1488 6 dbg_r0[9]
port 70 nsew signal output
rlabel metal3 s 79200 1368 80000 1488 6 i_clk
port 71 nsew signal input
rlabel metal3 s 79200 34688 80000 34808 6 i_flush
port 72 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 i_imm[0]
port 73 nsew signal input
rlabel metal2 s 26422 79200 26478 80000 6 i_imm[10]
port 74 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 i_imm[11]
port 75 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 i_imm[12]
port 76 nsew signal input
rlabel metal3 s 79200 71408 80000 71528 6 i_imm[13]
port 77 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 i_imm[14]
port 78 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 i_imm[15]
port 79 nsew signal input
rlabel metal3 s 0 54408 800 54528 6 i_imm[1]
port 80 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 i_imm[2]
port 81 nsew signal input
rlabel metal2 s 31574 79200 31630 80000 6 i_imm[3]
port 82 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 i_imm[4]
port 83 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 i_imm[5]
port 84 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 i_imm[6]
port 85 nsew signal input
rlabel metal2 s 53470 79200 53526 80000 6 i_imm[7]
port 86 nsew signal input
rlabel metal2 s 67638 0 67694 800 6 i_imm[8]
port 87 nsew signal input
rlabel metal3 s 79200 53048 80000 53168 6 i_imm[9]
port 88 nsew signal input
rlabel metal2 s 39302 79200 39358 80000 6 i_irq
port 89 nsew signal input
rlabel metal3 s 79200 45568 80000 45688 6 i_jmp_predict
port 90 nsew signal input
rlabel metal3 s 0 51688 800 51808 6 i_mem_exception
port 91 nsew signal input
rlabel metal2 s 79230 79200 79286 80000 6 i_next_ready
port 92 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 i_reg_data[0]
port 93 nsew signal input
rlabel metal2 s 50894 79200 50950 80000 6 i_reg_data[10]
port 94 nsew signal input
rlabel metal2 s 62486 79200 62542 80000 6 i_reg_data[11]
port 95 nsew signal input
rlabel metal3 s 79200 23128 80000 23248 6 i_reg_data[12]
port 96 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 i_reg_data[13]
port 97 nsew signal input
rlabel metal2 s 10322 79200 10378 80000 6 i_reg_data[14]
port 98 nsew signal input
rlabel metal2 s 21914 79200 21970 80000 6 i_reg_data[15]
port 99 nsew signal input
rlabel metal3 s 0 36048 800 36168 6 i_reg_data[1]
port 100 nsew signal input
rlabel metal2 s 46386 79200 46442 80000 6 i_reg_data[2]
port 101 nsew signal input
rlabel metal2 s 76010 0 76066 800 6 i_reg_data[3]
port 102 nsew signal input
rlabel metal3 s 0 17688 800 17808 6 i_reg_data[4]
port 103 nsew signal input
rlabel metal3 s 79200 4768 80000 4888 6 i_reg_data[5]
port 104 nsew signal input
rlabel metal2 s 17406 79200 17462 80000 6 i_reg_data[6]
port 105 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 i_reg_data[7]
port 106 nsew signal input
rlabel metal3 s 79200 63928 80000 64048 6 i_reg_data[8]
port 107 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 i_reg_data[9]
port 108 nsew signal input
rlabel metal3 s 79200 13608 80000 13728 6 i_reg_ie[0]
port 109 nsew signal input
rlabel metal3 s 79200 68688 80000 68808 6 i_reg_ie[1]
port 110 nsew signal input
rlabel metal3 s 79200 65288 80000 65408 6 i_reg_ie[2]
port 111 nsew signal input
rlabel metal2 s 28998 79200 29054 80000 6 i_reg_ie[3]
port 112 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 i_reg_ie[4]
port 113 nsew signal input
rlabel metal2 s 73434 0 73490 800 6 i_reg_ie[5]
port 114 nsew signal input
rlabel metal3 s 79200 50328 80000 50448 6 i_reg_ie[6]
port 115 nsew signal input
rlabel metal3 s 79200 62568 80000 62688 6 i_reg_ie[7]
port 116 nsew signal input
rlabel metal2 s 73434 79200 73490 80000 6 i_rst
port 117 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 i_submit
port 118 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 o_addr[0]
port 119 nsew signal output
rlabel metal3 s 79200 18368 80000 18488 6 o_addr[10]
port 120 nsew signal output
rlabel metal2 s 43166 79200 43222 80000 6 o_addr[11]
port 121 nsew signal output
rlabel metal2 s 35438 0 35494 800 6 o_addr[12]
port 122 nsew signal output
rlabel metal3 s 79200 10888 80000 11008 6 o_addr[13]
port 123 nsew signal output
rlabel metal3 s 0 59168 800 59288 6 o_addr[14]
port 124 nsew signal output
rlabel metal2 s 54758 0 54814 800 6 o_addr[15]
port 125 nsew signal output
rlabel metal2 s 11610 79200 11666 80000 6 o_addr[1]
port 126 nsew signal output
rlabel metal3 s 79200 42848 80000 42968 6 o_addr[2]
port 127 nsew signal output
rlabel metal2 s 32862 0 32918 800 6 o_addr[3]
port 128 nsew signal output
rlabel metal2 s 36082 79200 36138 80000 6 o_addr[4]
port 129 nsew signal output
rlabel metal3 s 0 2728 800 2848 6 o_addr[5]
port 130 nsew signal output
rlabel metal2 s 65062 79200 65118 80000 6 o_addr[6]
port 131 nsew signal output
rlabel metal2 s 31574 0 31630 800 6 o_addr[7]
port 132 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 o_addr[8]
port 133 nsew signal output
rlabel metal2 s 76654 79200 76710 80000 6 o_addr[9]
port 134 nsew signal output
rlabel metal3 s 79200 14968 80000 15088 6 o_c_data_page
port 135 nsew signal output
rlabel metal3 s 79200 39448 80000 39568 6 o_c_instr_page
port 136 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 o_data[0]
port 137 nsew signal output
rlabel metal3 s 79200 57808 80000 57928 6 o_data[10]
port 138 nsew signal output
rlabel metal3 s 79200 7488 80000 7608 6 o_data[11]
port 139 nsew signal output
rlabel metal2 s 47030 0 47086 800 6 o_data[12]
port 140 nsew signal output
rlabel metal3 s 0 53048 800 53168 6 o_data[13]
port 141 nsew signal output
rlabel metal2 s 18 79200 74 80000 6 o_data[14]
port 142 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 o_data[15]
port 143 nsew signal output
rlabel metal2 s 18694 79200 18750 80000 6 o_data[1]
port 144 nsew signal output
rlabel metal2 s 63130 0 63186 800 6 o_data[2]
port 145 nsew signal output
rlabel metal3 s 0 49648 800 49768 6 o_data[3]
port 146 nsew signal output
rlabel metal2 s 66350 79200 66406 80000 6 o_data[4]
port 147 nsew signal output
rlabel metal2 s 3238 79200 3294 80000 6 o_data[5]
port 148 nsew signal output
rlabel metal2 s 20626 79200 20682 80000 6 o_data[6]
port 149 nsew signal output
rlabel metal2 s 33506 79200 33562 80000 6 o_data[7]
port 150 nsew signal output
rlabel metal2 s 30286 79200 30342 80000 6 o_data[8]
port 151 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 o_data[9]
port 152 nsew signal output
rlabel metal2 s 12898 0 12954 800 6 o_exec_pc[0]
port 153 nsew signal output
rlabel metal3 s 79200 19728 80000 19848 6 o_exec_pc[10]
port 154 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 o_exec_pc[11]
port 155 nsew signal output
rlabel metal3 s 79200 76168 80000 76288 6 o_exec_pc[12]
port 156 nsew signal output
rlabel metal3 s 0 37408 800 37528 6 o_exec_pc[13]
port 157 nsew signal output
rlabel metal2 s 41878 79200 41934 80000 6 o_exec_pc[14]
port 158 nsew signal output
rlabel metal2 s 9678 0 9734 800 6 o_exec_pc[15]
port 159 nsew signal output
rlabel metal3 s 79200 27208 80000 27328 6 o_exec_pc[1]
port 160 nsew signal output
rlabel metal3 s 79200 59168 80000 59288 6 o_exec_pc[2]
port 161 nsew signal output
rlabel metal2 s 7102 79200 7158 80000 6 o_exec_pc[3]
port 162 nsew signal output
rlabel metal3 s 79200 40808 80000 40928 6 o_exec_pc[4]
port 163 nsew signal output
rlabel metal3 s 0 71408 800 71528 6 o_exec_pc[5]
port 164 nsew signal output
rlabel metal3 s 0 16328 800 16448 6 o_exec_pc[6]
port 165 nsew signal output
rlabel metal3 s 79200 70048 80000 70168 6 o_exec_pc[7]
port 166 nsew signal output
rlabel metal2 s 47674 79200 47730 80000 6 o_exec_pc[8]
port 167 nsew signal output
rlabel metal2 s 21270 0 21326 800 6 o_exec_pc[9]
port 168 nsew signal output
rlabel metal3 s 79200 31968 80000 32088 6 o_flush
port 169 nsew signal output
rlabel metal3 s 0 5448 800 5568 6 o_icache_flush
port 170 nsew signal output
rlabel metal3 s 79200 8848 80000 8968 6 o_mem_access
port 171 nsew signal output
rlabel metal3 s 0 75488 800 75608 6 o_mem_we
port 172 nsew signal output
rlabel metal2 s 71502 0 71558 800 6 o_mem_width
port 173 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 o_pc_update
port 174 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 o_ready
port 175 nsew signal output
rlabel metal3 s 79200 21088 80000 21208 6 o_reg_ie[0]
port 176 nsew signal output
rlabel metal3 s 79200 78888 80000 79008 6 o_reg_ie[1]
port 177 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 o_reg_ie[2]
port 178 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 o_reg_ie[3]
port 179 nsew signal output
rlabel metal3 s 0 31968 800 32088 6 o_reg_ie[4]
port 180 nsew signal output
rlabel metal3 s 79200 33328 80000 33448 6 o_reg_ie[5]
port 181 nsew signal output
rlabel metal2 s 1306 0 1362 800 6 o_reg_ie[6]
port 182 nsew signal output
rlabel metal3 s 79200 61208 80000 61328 6 o_reg_ie[7]
port 183 nsew signal output
rlabel metal2 s 75366 79200 75422 80000 6 o_submit
port 184 nsew signal output
rlabel metal3 s 79200 8 80000 128 6 sr_bus_addr[0]
port 185 nsew signal output
rlabel metal2 s 72146 79200 72202 80000 6 sr_bus_addr[10]
port 186 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 sr_bus_addr[11]
port 187 nsew signal output
rlabel metal3 s 0 46928 800 47048 6 sr_bus_addr[12]
port 188 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 sr_bus_addr[13]
port 189 nsew signal output
rlabel metal2 s 18 0 74 800 6 sr_bus_addr[14]
port 190 nsew signal output
rlabel metal2 s 57334 0 57390 800 6 sr_bus_addr[15]
port 191 nsew signal output
rlabel metal3 s 0 55768 800 55888 6 sr_bus_addr[1]
port 192 nsew signal output
rlabel metal2 s 5814 79200 5870 80000 6 sr_bus_addr[2]
port 193 nsew signal output
rlabel metal3 s 0 28568 800 28688 6 sr_bus_addr[3]
port 194 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 sr_bus_addr[4]
port 195 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 sr_bus_addr[5]
port 196 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 sr_bus_addr[6]
port 197 nsew signal output
rlabel metal2 s 52182 79200 52238 80000 6 sr_bus_addr[7]
port 198 nsew signal output
rlabel metal2 s 34794 79200 34850 80000 6 sr_bus_addr[8]
port 199 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 sr_bus_addr[9]
port 200 nsew signal output
rlabel metal2 s 63774 79200 63830 80000 6 sr_bus_data_o[0]
port 201 nsew signal output
rlabel metal3 s 79200 17008 80000 17128 6 sr_bus_data_o[10]
port 202 nsew signal output
rlabel metal3 s 0 63928 800 64048 6 sr_bus_data_o[11]
port 203 nsew signal output
rlabel metal3 s 79200 56448 80000 56568 6 sr_bus_data_o[12]
port 204 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 sr_bus_data_o[13]
port 205 nsew signal output
rlabel metal2 s 28354 0 28410 800 6 sr_bus_data_o[14]
port 206 nsew signal output
rlabel metal3 s 0 13608 800 13728 6 sr_bus_data_o[15]
port 207 nsew signal output
rlabel metal3 s 79200 55088 80000 55208 6 sr_bus_data_o[1]
port 208 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 sr_bus_data_o[2]
port 209 nsew signal output
rlabel metal2 s 56690 79200 56746 80000 6 sr_bus_data_o[3]
port 210 nsew signal output
rlabel metal2 s 54758 79200 54814 80000 6 sr_bus_data_o[4]
port 211 nsew signal output
rlabel metal3 s 0 78888 800 79008 6 sr_bus_data_o[5]
port 212 nsew signal output
rlabel metal2 s 12898 79200 12954 80000 6 sr_bus_data_o[6]
port 213 nsew signal output
rlabel metal2 s 56046 0 56102 800 6 sr_bus_data_o[7]
port 214 nsew signal output
rlabel metal3 s 0 19728 800 19848 6 sr_bus_data_o[8]
port 215 nsew signal output
rlabel metal3 s 0 68008 800 68128 6 sr_bus_data_o[9]
port 216 nsew signal output
rlabel metal3 s 79200 38088 80000 38208 6 sr_bus_we
port 217 nsew signal output
rlabel metal4 s 4208 2128 4528 77840 6 vccd1
port 218 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 77840 6 vccd1
port 218 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 77840 6 vccd1
port 218 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 77840 6 vssd1
port 219 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 77840 6 vssd1
port 219 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 80000 80000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 11769936
string GDS_FILE /home/piotro/ppcpu_caravel/openlane/execute/runs/22_09_08_19_20/results/signoff/execute.magic.gds
string GDS_START 1279502
<< end >>

