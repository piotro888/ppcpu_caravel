magic
tech sky130B
magscale 1 2
timestamp 1663070791
<< nwell >>
rect 1066 37253 38862 37574
rect 1066 36165 38862 36731
rect 1066 35077 38862 35643
rect 1066 33989 38862 34555
rect 1066 32901 38862 33467
rect 1066 31813 38862 32379
rect 1066 30725 38862 31291
rect 1066 29637 38862 30203
rect 1066 28549 38862 29115
rect 1066 27461 38862 28027
rect 1066 26373 38862 26939
rect 1066 25285 38862 25851
rect 1066 24197 38862 24763
rect 1066 23109 38862 23675
rect 1066 22021 38862 22587
rect 1066 20933 38862 21499
rect 1066 19845 38862 20411
rect 1066 18757 38862 19323
rect 1066 17669 38862 18235
rect 1066 16581 38862 17147
rect 1066 15493 38862 16059
rect 1066 14405 38862 14971
rect 1066 13317 38862 13883
rect 1066 12229 38862 12795
rect 1066 11141 38862 11707
rect 1066 10053 38862 10619
rect 1066 8965 38862 9531
rect 1066 7877 38862 8443
rect 1066 6789 38862 7355
rect 1066 5701 38862 6267
rect 1066 4613 38862 5179
rect 1066 3525 38862 4091
rect 1066 2437 38862 3003
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 1104 1368 38824 37732
<< metal2 >>
rect 1766 39200 1822 40000
rect 2318 39200 2374 40000
rect 2870 39200 2926 40000
rect 3422 39200 3478 40000
rect 3974 39200 4030 40000
rect 4526 39200 4582 40000
rect 5078 39200 5134 40000
rect 5630 39200 5686 40000
rect 6182 39200 6238 40000
rect 6734 39200 6790 40000
rect 7286 39200 7342 40000
rect 7838 39200 7894 40000
rect 8390 39200 8446 40000
rect 8942 39200 8998 40000
rect 9494 39200 9550 40000
rect 10046 39200 10102 40000
rect 10598 39200 10654 40000
rect 11150 39200 11206 40000
rect 11702 39200 11758 40000
rect 12254 39200 12310 40000
rect 12806 39200 12862 40000
rect 13358 39200 13414 40000
rect 13910 39200 13966 40000
rect 14462 39200 14518 40000
rect 15014 39200 15070 40000
rect 15566 39200 15622 40000
rect 16118 39200 16174 40000
rect 16670 39200 16726 40000
rect 17222 39200 17278 40000
rect 17774 39200 17830 40000
rect 18326 39200 18382 40000
rect 18878 39200 18934 40000
rect 19430 39200 19486 40000
rect 19982 39200 20038 40000
rect 20534 39200 20590 40000
rect 21086 39200 21142 40000
rect 21638 39200 21694 40000
rect 22190 39200 22246 40000
rect 22742 39200 22798 40000
rect 23294 39200 23350 40000
rect 23846 39200 23902 40000
rect 24398 39200 24454 40000
rect 24950 39200 25006 40000
rect 25502 39200 25558 40000
rect 26054 39200 26110 40000
rect 26606 39200 26662 40000
rect 27158 39200 27214 40000
rect 27710 39200 27766 40000
rect 28262 39200 28318 40000
rect 28814 39200 28870 40000
rect 29366 39200 29422 40000
rect 29918 39200 29974 40000
rect 30470 39200 30526 40000
rect 31022 39200 31078 40000
rect 31574 39200 31630 40000
rect 32126 39200 32182 40000
rect 32678 39200 32734 40000
rect 33230 39200 33286 40000
rect 33782 39200 33838 40000
rect 34334 39200 34390 40000
rect 34886 39200 34942 40000
rect 35438 39200 35494 40000
rect 35990 39200 36046 40000
rect 36542 39200 36598 40000
rect 37094 39200 37150 40000
rect 37646 39200 37702 40000
rect 38198 39200 38254 40000
rect 1766 0 1822 800
rect 2318 0 2374 800
rect 2870 0 2926 800
rect 3422 0 3478 800
rect 3974 0 4030 800
rect 4526 0 4582 800
rect 5078 0 5134 800
rect 5630 0 5686 800
rect 6182 0 6238 800
rect 6734 0 6790 800
rect 7286 0 7342 800
rect 7838 0 7894 800
rect 8390 0 8446 800
rect 8942 0 8998 800
rect 9494 0 9550 800
rect 10046 0 10102 800
rect 10598 0 10654 800
rect 11150 0 11206 800
rect 11702 0 11758 800
rect 12254 0 12310 800
rect 12806 0 12862 800
rect 13358 0 13414 800
rect 13910 0 13966 800
rect 14462 0 14518 800
rect 15014 0 15070 800
rect 15566 0 15622 800
rect 16118 0 16174 800
rect 16670 0 16726 800
rect 17222 0 17278 800
rect 17774 0 17830 800
rect 18326 0 18382 800
rect 18878 0 18934 800
rect 19430 0 19486 800
rect 19982 0 20038 800
rect 20534 0 20590 800
rect 21086 0 21142 800
rect 21638 0 21694 800
rect 22190 0 22246 800
rect 22742 0 22798 800
rect 23294 0 23350 800
rect 23846 0 23902 800
rect 24398 0 24454 800
rect 24950 0 25006 800
rect 25502 0 25558 800
rect 26054 0 26110 800
rect 26606 0 26662 800
rect 27158 0 27214 800
rect 27710 0 27766 800
rect 28262 0 28318 800
rect 28814 0 28870 800
rect 29366 0 29422 800
rect 29918 0 29974 800
rect 30470 0 30526 800
rect 31022 0 31078 800
rect 31574 0 31630 800
rect 32126 0 32182 800
rect 32678 0 32734 800
rect 33230 0 33286 800
rect 33782 0 33838 800
rect 34334 0 34390 800
rect 34886 0 34942 800
rect 35438 0 35494 800
rect 35990 0 36046 800
rect 36542 0 36598 800
rect 37094 0 37150 800
rect 37646 0 37702 800
rect 38198 0 38254 800
<< obsm2 >>
rect 1878 39144 2262 39250
rect 2430 39144 2814 39250
rect 2982 39144 3366 39250
rect 3534 39144 3918 39250
rect 4086 39144 4470 39250
rect 4638 39144 5022 39250
rect 5190 39144 5574 39250
rect 5742 39144 6126 39250
rect 6294 39144 6678 39250
rect 6846 39144 7230 39250
rect 7398 39144 7782 39250
rect 7950 39144 8334 39250
rect 8502 39144 8886 39250
rect 9054 39144 9438 39250
rect 9606 39144 9990 39250
rect 10158 39144 10542 39250
rect 10710 39144 11094 39250
rect 11262 39144 11646 39250
rect 11814 39144 12198 39250
rect 12366 39144 12750 39250
rect 12918 39144 13302 39250
rect 13470 39144 13854 39250
rect 14022 39144 14406 39250
rect 14574 39144 14958 39250
rect 15126 39144 15510 39250
rect 15678 39144 16062 39250
rect 16230 39144 16614 39250
rect 16782 39144 17166 39250
rect 17334 39144 17718 39250
rect 17886 39144 18270 39250
rect 18438 39144 18822 39250
rect 18990 39144 19374 39250
rect 19542 39144 19926 39250
rect 20094 39144 20478 39250
rect 20646 39144 21030 39250
rect 21198 39144 21582 39250
rect 21750 39144 22134 39250
rect 22302 39144 22686 39250
rect 22854 39144 23238 39250
rect 23406 39144 23790 39250
rect 23958 39144 24342 39250
rect 24510 39144 24894 39250
rect 25062 39144 25446 39250
rect 25614 39144 25998 39250
rect 26166 39144 26550 39250
rect 26718 39144 27102 39250
rect 27270 39144 27654 39250
rect 27822 39144 28206 39250
rect 28374 39144 28758 39250
rect 28926 39144 29310 39250
rect 29478 39144 29862 39250
rect 30030 39144 30414 39250
rect 30582 39144 30966 39250
rect 31134 39144 31518 39250
rect 31686 39144 32070 39250
rect 32238 39144 32622 39250
rect 32790 39144 33174 39250
rect 33342 39144 33726 39250
rect 33894 39144 34278 39250
rect 34446 39144 34830 39250
rect 34998 39144 35382 39250
rect 35550 39144 35934 39250
rect 36102 39144 36486 39250
rect 36654 39144 37038 39250
rect 37206 39144 37590 39250
rect 37758 39144 38142 39250
rect 38310 39144 38346 39250
rect 1768 856 38346 39144
rect 1878 734 2262 856
rect 2430 734 2814 856
rect 2982 734 3366 856
rect 3534 734 3918 856
rect 4086 734 4470 856
rect 4638 734 5022 856
rect 5190 734 5574 856
rect 5742 734 6126 856
rect 6294 734 6678 856
rect 6846 734 7230 856
rect 7398 734 7782 856
rect 7950 734 8334 856
rect 8502 734 8886 856
rect 9054 734 9438 856
rect 9606 734 9990 856
rect 10158 734 10542 856
rect 10710 734 11094 856
rect 11262 734 11646 856
rect 11814 734 12198 856
rect 12366 734 12750 856
rect 12918 734 13302 856
rect 13470 734 13854 856
rect 14022 734 14406 856
rect 14574 734 14958 856
rect 15126 734 15510 856
rect 15678 734 16062 856
rect 16230 734 16614 856
rect 16782 734 17166 856
rect 17334 734 17718 856
rect 17886 734 18270 856
rect 18438 734 18822 856
rect 18990 734 19374 856
rect 19542 734 19926 856
rect 20094 734 20478 856
rect 20646 734 21030 856
rect 21198 734 21582 856
rect 21750 734 22134 856
rect 22302 734 22686 856
rect 22854 734 23238 856
rect 23406 734 23790 856
rect 23958 734 24342 856
rect 24510 734 24894 856
rect 25062 734 25446 856
rect 25614 734 25998 856
rect 26166 734 26550 856
rect 26718 734 27102 856
rect 27270 734 27654 856
rect 27822 734 28206 856
rect 28374 734 28758 856
rect 28926 734 29310 856
rect 29478 734 29862 856
rect 30030 734 30414 856
rect 30582 734 30966 856
rect 31134 734 31518 856
rect 31686 734 32070 856
rect 32238 734 32622 856
rect 32790 734 33174 856
rect 33342 734 33726 856
rect 33894 734 34278 856
rect 34446 734 34830 856
rect 34998 734 35382 856
rect 35550 734 35934 856
rect 36102 734 36486 856
rect 36654 734 37038 856
rect 37206 734 37590 856
rect 37758 734 38142 856
rect 38310 734 38346 856
<< obsm3 >>
rect 4210 1667 38351 37569
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< obsm4 >>
rect 18643 2048 19488 36549
rect 19968 2048 34848 36549
rect 35328 2048 36557 36549
rect 18643 1667 36557 2048
<< labels >>
rlabel metal2 s 38198 0 38254 800 6 clk_m
port 1 nsew signal input
rlabel metal2 s 38198 39200 38254 40000 6 clk_s
port 2 nsew signal input
rlabel metal2 s 1766 0 1822 800 6 m_rst
port 3 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 m_wb_4_burst
port 4 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 m_wb_8_burst
port 5 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 m_wb_ack
port 6 nsew signal output
rlabel metal2 s 3974 0 4030 800 6 m_wb_adr[0]
port 7 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 m_wb_adr[10]
port 8 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 m_wb_adr[11]
port 9 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 m_wb_adr[12]
port 10 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 m_wb_adr[13]
port 11 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 m_wb_adr[14]
port 12 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 m_wb_adr[15]
port 13 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 m_wb_adr[16]
port 14 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 m_wb_adr[17]
port 15 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 m_wb_adr[18]
port 16 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 m_wb_adr[19]
port 17 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 m_wb_adr[1]
port 18 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 m_wb_adr[20]
port 19 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 m_wb_adr[21]
port 20 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 m_wb_adr[22]
port 21 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 m_wb_adr[23]
port 22 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 m_wb_adr[2]
port 23 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 m_wb_adr[3]
port 24 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 m_wb_adr[4]
port 25 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 m_wb_adr[5]
port 26 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 m_wb_adr[6]
port 27 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 m_wb_adr[7]
port 28 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 m_wb_adr[8]
port 29 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 m_wb_adr[9]
port 30 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 m_wb_cyc
port 31 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 m_wb_err
port 32 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 m_wb_i_dat[0]
port 33 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 m_wb_i_dat[10]
port 34 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 m_wb_i_dat[11]
port 35 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 m_wb_i_dat[12]
port 36 nsew signal output
rlabel metal2 s 25502 0 25558 800 6 m_wb_i_dat[13]
port 37 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 m_wb_i_dat[14]
port 38 nsew signal output
rlabel metal2 s 26606 0 26662 800 6 m_wb_i_dat[15]
port 39 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 m_wb_i_dat[1]
port 40 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 m_wb_i_dat[2]
port 41 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 m_wb_i_dat[3]
port 42 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 m_wb_i_dat[4]
port 43 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 m_wb_i_dat[5]
port 44 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 m_wb_i_dat[6]
port 45 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 m_wb_i_dat[7]
port 46 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 m_wb_i_dat[8]
port 47 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 m_wb_i_dat[9]
port 48 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 m_wb_o_dat[0]
port 49 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 m_wb_o_dat[10]
port 50 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 m_wb_o_dat[11]
port 51 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 m_wb_o_dat[12]
port 52 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 m_wb_o_dat[13]
port 53 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 m_wb_o_dat[14]
port 54 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 m_wb_o_dat[15]
port 55 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 m_wb_o_dat[1]
port 56 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 m_wb_o_dat[2]
port 57 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 m_wb_o_dat[3]
port 58 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 m_wb_o_dat[4]
port 59 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 m_wb_o_dat[5]
port 60 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 m_wb_o_dat[6]
port 61 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 m_wb_o_dat[7]
port 62 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 m_wb_o_dat[8]
port 63 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 m_wb_o_dat[9]
port 64 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 m_wb_sel[0]
port 65 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 m_wb_sel[1]
port 66 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 m_wb_stb
port 67 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 m_wb_we
port 68 nsew signal input
rlabel metal2 s 1766 39200 1822 40000 6 s_rst
port 69 nsew signal input
rlabel metal2 s 2318 39200 2374 40000 6 s_wb_4_burst
port 70 nsew signal output
rlabel metal2 s 2870 39200 2926 40000 6 s_wb_8_burst
port 71 nsew signal output
rlabel metal2 s 3422 39200 3478 40000 6 s_wb_ack
port 72 nsew signal input
rlabel metal2 s 3974 39200 4030 40000 6 s_wb_adr[0]
port 73 nsew signal output
rlabel metal2 s 9494 39200 9550 40000 6 s_wb_adr[10]
port 74 nsew signal output
rlabel metal2 s 10046 39200 10102 40000 6 s_wb_adr[11]
port 75 nsew signal output
rlabel metal2 s 10598 39200 10654 40000 6 s_wb_adr[12]
port 76 nsew signal output
rlabel metal2 s 11150 39200 11206 40000 6 s_wb_adr[13]
port 77 nsew signal output
rlabel metal2 s 11702 39200 11758 40000 6 s_wb_adr[14]
port 78 nsew signal output
rlabel metal2 s 12254 39200 12310 40000 6 s_wb_adr[15]
port 79 nsew signal output
rlabel metal2 s 12806 39200 12862 40000 6 s_wb_adr[16]
port 80 nsew signal output
rlabel metal2 s 13358 39200 13414 40000 6 s_wb_adr[17]
port 81 nsew signal output
rlabel metal2 s 13910 39200 13966 40000 6 s_wb_adr[18]
port 82 nsew signal output
rlabel metal2 s 14462 39200 14518 40000 6 s_wb_adr[19]
port 83 nsew signal output
rlabel metal2 s 4526 39200 4582 40000 6 s_wb_adr[1]
port 84 nsew signal output
rlabel metal2 s 15014 39200 15070 40000 6 s_wb_adr[20]
port 85 nsew signal output
rlabel metal2 s 15566 39200 15622 40000 6 s_wb_adr[21]
port 86 nsew signal output
rlabel metal2 s 16118 39200 16174 40000 6 s_wb_adr[22]
port 87 nsew signal output
rlabel metal2 s 16670 39200 16726 40000 6 s_wb_adr[23]
port 88 nsew signal output
rlabel metal2 s 5078 39200 5134 40000 6 s_wb_adr[2]
port 89 nsew signal output
rlabel metal2 s 5630 39200 5686 40000 6 s_wb_adr[3]
port 90 nsew signal output
rlabel metal2 s 6182 39200 6238 40000 6 s_wb_adr[4]
port 91 nsew signal output
rlabel metal2 s 6734 39200 6790 40000 6 s_wb_adr[5]
port 92 nsew signal output
rlabel metal2 s 7286 39200 7342 40000 6 s_wb_adr[6]
port 93 nsew signal output
rlabel metal2 s 7838 39200 7894 40000 6 s_wb_adr[7]
port 94 nsew signal output
rlabel metal2 s 8390 39200 8446 40000 6 s_wb_adr[8]
port 95 nsew signal output
rlabel metal2 s 8942 39200 8998 40000 6 s_wb_adr[9]
port 96 nsew signal output
rlabel metal2 s 17222 39200 17278 40000 6 s_wb_cyc
port 97 nsew signal output
rlabel metal2 s 17774 39200 17830 40000 6 s_wb_err
port 98 nsew signal input
rlabel metal2 s 18326 39200 18382 40000 6 s_wb_i_dat[0]
port 99 nsew signal input
rlabel metal2 s 23846 39200 23902 40000 6 s_wb_i_dat[10]
port 100 nsew signal input
rlabel metal2 s 24398 39200 24454 40000 6 s_wb_i_dat[11]
port 101 nsew signal input
rlabel metal2 s 24950 39200 25006 40000 6 s_wb_i_dat[12]
port 102 nsew signal input
rlabel metal2 s 25502 39200 25558 40000 6 s_wb_i_dat[13]
port 103 nsew signal input
rlabel metal2 s 26054 39200 26110 40000 6 s_wb_i_dat[14]
port 104 nsew signal input
rlabel metal2 s 26606 39200 26662 40000 6 s_wb_i_dat[15]
port 105 nsew signal input
rlabel metal2 s 18878 39200 18934 40000 6 s_wb_i_dat[1]
port 106 nsew signal input
rlabel metal2 s 19430 39200 19486 40000 6 s_wb_i_dat[2]
port 107 nsew signal input
rlabel metal2 s 19982 39200 20038 40000 6 s_wb_i_dat[3]
port 108 nsew signal input
rlabel metal2 s 20534 39200 20590 40000 6 s_wb_i_dat[4]
port 109 nsew signal input
rlabel metal2 s 21086 39200 21142 40000 6 s_wb_i_dat[5]
port 110 nsew signal input
rlabel metal2 s 21638 39200 21694 40000 6 s_wb_i_dat[6]
port 111 nsew signal input
rlabel metal2 s 22190 39200 22246 40000 6 s_wb_i_dat[7]
port 112 nsew signal input
rlabel metal2 s 22742 39200 22798 40000 6 s_wb_i_dat[8]
port 113 nsew signal input
rlabel metal2 s 23294 39200 23350 40000 6 s_wb_i_dat[9]
port 114 nsew signal input
rlabel metal2 s 27158 39200 27214 40000 6 s_wb_o_dat[0]
port 115 nsew signal output
rlabel metal2 s 32678 39200 32734 40000 6 s_wb_o_dat[10]
port 116 nsew signal output
rlabel metal2 s 33230 39200 33286 40000 6 s_wb_o_dat[11]
port 117 nsew signal output
rlabel metal2 s 33782 39200 33838 40000 6 s_wb_o_dat[12]
port 118 nsew signal output
rlabel metal2 s 34334 39200 34390 40000 6 s_wb_o_dat[13]
port 119 nsew signal output
rlabel metal2 s 34886 39200 34942 40000 6 s_wb_o_dat[14]
port 120 nsew signal output
rlabel metal2 s 35438 39200 35494 40000 6 s_wb_o_dat[15]
port 121 nsew signal output
rlabel metal2 s 27710 39200 27766 40000 6 s_wb_o_dat[1]
port 122 nsew signal output
rlabel metal2 s 28262 39200 28318 40000 6 s_wb_o_dat[2]
port 123 nsew signal output
rlabel metal2 s 28814 39200 28870 40000 6 s_wb_o_dat[3]
port 124 nsew signal output
rlabel metal2 s 29366 39200 29422 40000 6 s_wb_o_dat[4]
port 125 nsew signal output
rlabel metal2 s 29918 39200 29974 40000 6 s_wb_o_dat[5]
port 126 nsew signal output
rlabel metal2 s 30470 39200 30526 40000 6 s_wb_o_dat[6]
port 127 nsew signal output
rlabel metal2 s 31022 39200 31078 40000 6 s_wb_o_dat[7]
port 128 nsew signal output
rlabel metal2 s 31574 39200 31630 40000 6 s_wb_o_dat[8]
port 129 nsew signal output
rlabel metal2 s 32126 39200 32182 40000 6 s_wb_o_dat[9]
port 130 nsew signal output
rlabel metal2 s 35990 39200 36046 40000 6 s_wb_sel[0]
port 131 nsew signal output
rlabel metal2 s 36542 39200 36598 40000 6 s_wb_sel[1]
port 132 nsew signal output
rlabel metal2 s 37094 39200 37150 40000 6 s_wb_stb
port 133 nsew signal output
rlabel metal2 s 37646 39200 37702 40000 6 s_wb_we
port 134 nsew signal output
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 135 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 135 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 136 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 2470728
string GDS_FILE /home/piotro/ppcpu_caravel/openlane/wb_cross_clk/runs/22_09_13_14_04/results/signoff/wb_cross_clk.magic.gds
string GDS_START 280276
<< end >>

