VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO int_ram
  CLASS BLOCK ;
  FOREIGN int_ram ;
  ORIGIN 0.000 0.000 ;
  SIZE 550.000 BY 550.000 ;
  PIN i_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 42.200 550.000 42.800 ;
    END
  END i_addr[0]
  PIN i_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 80.960 550.000 81.560 ;
    END
  END i_addr[1]
  PIN i_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 119.720 550.000 120.320 ;
    END
  END i_addr[2]
  PIN i_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 158.480 550.000 159.080 ;
    END
  END i_addr[3]
  PIN i_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 197.240 550.000 197.840 ;
    END
  END i_addr[4]
  PIN i_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 236.000 550.000 236.600 ;
    END
  END i_addr[5]
  PIN i_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 274.760 550.000 275.360 ;
    END
  END i_addr[6]
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 16.360 550.000 16.960 ;
    END
  END i_clk
  PIN i_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 55.120 550.000 55.720 ;
    END
  END i_data[0]
  PIN i_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 391.040 550.000 391.640 ;
    END
  END i_data[10]
  PIN i_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 416.880 550.000 417.480 ;
    END
  END i_data[11]
  PIN i_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 442.720 550.000 443.320 ;
    END
  END i_data[12]
  PIN i_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 468.560 550.000 469.160 ;
    END
  END i_data[13]
  PIN i_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 494.400 550.000 495.000 ;
    END
  END i_data[14]
  PIN i_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 520.240 550.000 520.840 ;
    END
  END i_data[15]
  PIN i_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 93.880 550.000 94.480 ;
    END
  END i_data[1]
  PIN i_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 132.640 550.000 133.240 ;
    END
  END i_data[2]
  PIN i_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 171.400 550.000 172.000 ;
    END
  END i_data[3]
  PIN i_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 210.160 550.000 210.760 ;
    END
  END i_data[4]
  PIN i_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 248.920 550.000 249.520 ;
    END
  END i_data[5]
  PIN i_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 287.680 550.000 288.280 ;
    END
  END i_data[6]
  PIN i_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 313.520 550.000 314.120 ;
    END
  END i_data[7]
  PIN i_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 339.360 550.000 339.960 ;
    END
  END i_data[8]
  PIN i_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 365.200 550.000 365.800 ;
    END
  END i_data[9]
  PIN i_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 29.280 550.000 29.880 ;
    END
  END i_we
  PIN o_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 68.040 550.000 68.640 ;
    END
  END o_data[0]
  PIN o_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 403.960 550.000 404.560 ;
    END
  END o_data[10]
  PIN o_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 429.800 550.000 430.400 ;
    END
  END o_data[11]
  PIN o_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 455.640 550.000 456.240 ;
    END
  END o_data[12]
  PIN o_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 481.480 550.000 482.080 ;
    END
  END o_data[13]
  PIN o_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 507.320 550.000 507.920 ;
    END
  END o_data[14]
  PIN o_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 533.160 550.000 533.760 ;
    END
  END o_data[15]
  PIN o_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 106.800 550.000 107.400 ;
    END
  END o_data[1]
  PIN o_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 145.560 550.000 146.160 ;
    END
  END o_data[2]
  PIN o_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 184.320 550.000 184.920 ;
    END
  END o_data[3]
  PIN o_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 223.080 550.000 223.680 ;
    END
  END o_data[4]
  PIN o_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 261.840 550.000 262.440 ;
    END
  END o_data[5]
  PIN o_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 300.600 550.000 301.200 ;
    END
  END o_data[6]
  PIN o_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 326.440 550.000 327.040 ;
    END
  END o_data[7]
  PIN o_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 352.280 550.000 352.880 ;
    END
  END o_data[8]
  PIN o_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 546.000 378.120 550.000 378.720 ;
    END
  END o_data[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 538.800 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 538.800 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 538.800 ;
    END
  END vssd1
  OBS
      LAYER nwell ;
        RECT 5.330 534.425 544.370 537.255 ;
        RECT 5.330 528.985 544.370 531.815 ;
        RECT 5.330 523.545 544.370 526.375 ;
        RECT 5.330 518.105 544.370 520.935 ;
        RECT 5.330 512.665 544.370 515.495 ;
        RECT 5.330 507.225 544.370 510.055 ;
        RECT 5.330 501.785 544.370 504.615 ;
        RECT 5.330 496.345 544.370 499.175 ;
        RECT 5.330 490.905 544.370 493.735 ;
        RECT 5.330 485.465 544.370 488.295 ;
        RECT 5.330 480.025 544.370 482.855 ;
        RECT 5.330 474.585 544.370 477.415 ;
        RECT 5.330 469.145 544.370 471.975 ;
        RECT 5.330 463.705 544.370 466.535 ;
        RECT 5.330 458.265 544.370 461.095 ;
        RECT 5.330 452.825 544.370 455.655 ;
        RECT 5.330 447.385 544.370 450.215 ;
        RECT 5.330 441.945 544.370 444.775 ;
        RECT 5.330 436.505 544.370 439.335 ;
        RECT 5.330 431.065 544.370 433.895 ;
        RECT 5.330 425.625 544.370 428.455 ;
        RECT 5.330 420.185 544.370 423.015 ;
        RECT 5.330 414.745 544.370 417.575 ;
        RECT 5.330 409.305 544.370 412.135 ;
        RECT 5.330 403.865 544.370 406.695 ;
        RECT 5.330 398.425 544.370 401.255 ;
        RECT 5.330 392.985 544.370 395.815 ;
        RECT 5.330 387.545 544.370 390.375 ;
        RECT 5.330 382.105 544.370 384.935 ;
        RECT 5.330 376.665 544.370 379.495 ;
        RECT 5.330 371.225 544.370 374.055 ;
        RECT 5.330 365.785 544.370 368.615 ;
        RECT 5.330 360.345 544.370 363.175 ;
        RECT 5.330 354.905 544.370 357.735 ;
        RECT 5.330 349.465 544.370 352.295 ;
        RECT 5.330 344.025 544.370 346.855 ;
        RECT 5.330 338.585 544.370 341.415 ;
        RECT 5.330 333.145 544.370 335.975 ;
        RECT 5.330 327.705 544.370 330.535 ;
        RECT 5.330 322.265 544.370 325.095 ;
        RECT 5.330 316.825 544.370 319.655 ;
        RECT 5.330 311.385 544.370 314.215 ;
        RECT 5.330 305.945 544.370 308.775 ;
        RECT 5.330 300.505 544.370 303.335 ;
        RECT 5.330 295.065 544.370 297.895 ;
        RECT 5.330 289.625 544.370 292.455 ;
        RECT 5.330 284.185 544.370 287.015 ;
        RECT 5.330 278.745 544.370 281.575 ;
        RECT 5.330 273.305 544.370 276.135 ;
        RECT 5.330 267.865 544.370 270.695 ;
        RECT 5.330 262.425 544.370 265.255 ;
        RECT 5.330 256.985 544.370 259.815 ;
        RECT 5.330 251.545 544.370 254.375 ;
        RECT 5.330 246.105 544.370 248.935 ;
        RECT 5.330 240.665 544.370 243.495 ;
        RECT 5.330 235.225 544.370 238.055 ;
        RECT 5.330 229.785 544.370 232.615 ;
        RECT 5.330 224.345 544.370 227.175 ;
        RECT 5.330 218.905 544.370 221.735 ;
        RECT 5.330 213.465 544.370 216.295 ;
        RECT 5.330 208.025 544.370 210.855 ;
        RECT 5.330 202.585 544.370 205.415 ;
        RECT 5.330 197.145 544.370 199.975 ;
        RECT 5.330 191.705 544.370 194.535 ;
        RECT 5.330 186.265 544.370 189.095 ;
        RECT 5.330 180.825 544.370 183.655 ;
        RECT 5.330 175.385 544.370 178.215 ;
        RECT 5.330 169.945 544.370 172.775 ;
        RECT 5.330 164.505 544.370 167.335 ;
        RECT 5.330 159.065 544.370 161.895 ;
        RECT 5.330 153.625 544.370 156.455 ;
        RECT 5.330 148.185 544.370 151.015 ;
        RECT 5.330 142.745 544.370 145.575 ;
        RECT 5.330 137.305 544.370 140.135 ;
        RECT 5.330 131.865 544.370 134.695 ;
        RECT 5.330 126.425 544.370 129.255 ;
        RECT 5.330 120.985 544.370 123.815 ;
        RECT 5.330 115.545 544.370 118.375 ;
        RECT 5.330 110.105 544.370 112.935 ;
        RECT 5.330 104.665 544.370 107.495 ;
        RECT 5.330 99.225 544.370 102.055 ;
        RECT 5.330 93.785 544.370 96.615 ;
        RECT 5.330 88.345 544.370 91.175 ;
        RECT 5.330 82.905 544.370 85.735 ;
        RECT 5.330 77.465 544.370 80.295 ;
        RECT 5.330 72.025 544.370 74.855 ;
        RECT 5.330 66.585 544.370 69.415 ;
        RECT 5.330 61.145 544.370 63.975 ;
        RECT 5.330 55.705 544.370 58.535 ;
        RECT 5.330 50.265 544.370 53.095 ;
        RECT 5.330 44.825 544.370 47.655 ;
        RECT 5.330 39.385 544.370 42.215 ;
        RECT 5.330 33.945 544.370 36.775 ;
        RECT 5.330 28.505 544.370 31.335 ;
        RECT 5.330 23.065 544.370 25.895 ;
        RECT 5.330 17.625 544.370 20.455 ;
        RECT 5.330 12.185 544.370 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 544.180 538.645 ;
      LAYER met1 ;
        RECT 5.520 9.220 545.030 538.800 ;
      LAYER met2 ;
        RECT 7.920 9.190 545.000 538.745 ;
      LAYER met3 ;
        RECT 14.785 534.160 546.000 538.725 ;
        RECT 14.785 532.760 545.600 534.160 ;
        RECT 14.785 521.240 546.000 532.760 ;
        RECT 14.785 519.840 545.600 521.240 ;
        RECT 14.785 508.320 546.000 519.840 ;
        RECT 14.785 506.920 545.600 508.320 ;
        RECT 14.785 495.400 546.000 506.920 ;
        RECT 14.785 494.000 545.600 495.400 ;
        RECT 14.785 482.480 546.000 494.000 ;
        RECT 14.785 481.080 545.600 482.480 ;
        RECT 14.785 469.560 546.000 481.080 ;
        RECT 14.785 468.160 545.600 469.560 ;
        RECT 14.785 456.640 546.000 468.160 ;
        RECT 14.785 455.240 545.600 456.640 ;
        RECT 14.785 443.720 546.000 455.240 ;
        RECT 14.785 442.320 545.600 443.720 ;
        RECT 14.785 430.800 546.000 442.320 ;
        RECT 14.785 429.400 545.600 430.800 ;
        RECT 14.785 417.880 546.000 429.400 ;
        RECT 14.785 416.480 545.600 417.880 ;
        RECT 14.785 404.960 546.000 416.480 ;
        RECT 14.785 403.560 545.600 404.960 ;
        RECT 14.785 392.040 546.000 403.560 ;
        RECT 14.785 390.640 545.600 392.040 ;
        RECT 14.785 379.120 546.000 390.640 ;
        RECT 14.785 377.720 545.600 379.120 ;
        RECT 14.785 366.200 546.000 377.720 ;
        RECT 14.785 364.800 545.600 366.200 ;
        RECT 14.785 353.280 546.000 364.800 ;
        RECT 14.785 351.880 545.600 353.280 ;
        RECT 14.785 340.360 546.000 351.880 ;
        RECT 14.785 338.960 545.600 340.360 ;
        RECT 14.785 327.440 546.000 338.960 ;
        RECT 14.785 326.040 545.600 327.440 ;
        RECT 14.785 314.520 546.000 326.040 ;
        RECT 14.785 313.120 545.600 314.520 ;
        RECT 14.785 301.600 546.000 313.120 ;
        RECT 14.785 300.200 545.600 301.600 ;
        RECT 14.785 288.680 546.000 300.200 ;
        RECT 14.785 287.280 545.600 288.680 ;
        RECT 14.785 275.760 546.000 287.280 ;
        RECT 14.785 274.360 545.600 275.760 ;
        RECT 14.785 262.840 546.000 274.360 ;
        RECT 14.785 261.440 545.600 262.840 ;
        RECT 14.785 249.920 546.000 261.440 ;
        RECT 14.785 248.520 545.600 249.920 ;
        RECT 14.785 237.000 546.000 248.520 ;
        RECT 14.785 235.600 545.600 237.000 ;
        RECT 14.785 224.080 546.000 235.600 ;
        RECT 14.785 222.680 545.600 224.080 ;
        RECT 14.785 211.160 546.000 222.680 ;
        RECT 14.785 209.760 545.600 211.160 ;
        RECT 14.785 198.240 546.000 209.760 ;
        RECT 14.785 196.840 545.600 198.240 ;
        RECT 14.785 185.320 546.000 196.840 ;
        RECT 14.785 183.920 545.600 185.320 ;
        RECT 14.785 172.400 546.000 183.920 ;
        RECT 14.785 171.000 545.600 172.400 ;
        RECT 14.785 159.480 546.000 171.000 ;
        RECT 14.785 158.080 545.600 159.480 ;
        RECT 14.785 146.560 546.000 158.080 ;
        RECT 14.785 145.160 545.600 146.560 ;
        RECT 14.785 133.640 546.000 145.160 ;
        RECT 14.785 132.240 545.600 133.640 ;
        RECT 14.785 120.720 546.000 132.240 ;
        RECT 14.785 119.320 545.600 120.720 ;
        RECT 14.785 107.800 546.000 119.320 ;
        RECT 14.785 106.400 545.600 107.800 ;
        RECT 14.785 94.880 546.000 106.400 ;
        RECT 14.785 93.480 545.600 94.880 ;
        RECT 14.785 81.960 546.000 93.480 ;
        RECT 14.785 80.560 545.600 81.960 ;
        RECT 14.785 69.040 546.000 80.560 ;
        RECT 14.785 67.640 545.600 69.040 ;
        RECT 14.785 56.120 546.000 67.640 ;
        RECT 14.785 54.720 545.600 56.120 ;
        RECT 14.785 43.200 546.000 54.720 ;
        RECT 14.785 41.800 545.600 43.200 ;
        RECT 14.785 30.280 546.000 41.800 ;
        RECT 14.785 28.880 545.600 30.280 ;
        RECT 14.785 17.360 546.000 28.880 ;
        RECT 14.785 15.960 545.600 17.360 ;
        RECT 14.785 10.715 546.000 15.960 ;
      LAYER met4 ;
        RECT 67.455 13.095 97.440 534.985 ;
        RECT 99.840 13.095 174.240 534.985 ;
        RECT 176.640 13.095 251.040 534.985 ;
        RECT 253.440 13.095 327.840 534.985 ;
        RECT 330.240 13.095 404.640 534.985 ;
        RECT 407.040 13.095 481.440 534.985 ;
        RECT 483.840 13.095 537.905 534.985 ;
  END
END int_ram
END LIBRARY

