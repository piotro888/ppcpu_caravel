magic
tech sky130B
magscale 1 2
timestamp 1662930718
<< viali >>
rect 30573 37417 30607 37451
rect 14749 37281 14783 37315
rect 14565 37213 14599 37247
rect 31217 37213 31251 37247
rect 31033 37077 31067 37111
rect 14289 36873 14323 36907
rect 6377 35649 6411 35683
rect 6644 35649 6678 35683
rect 8769 35649 8803 35683
rect 9036 35649 9070 35683
rect 7757 35445 7791 35479
rect 10149 35445 10183 35479
rect 17233 35037 17267 35071
rect 16966 34969 17000 35003
rect 15853 34901 15887 34935
rect 18061 34697 18095 34731
rect 16948 34561 16982 34595
rect 16681 34493 16715 34527
rect 15761 34153 15795 34187
rect 17141 33949 17175 33983
rect 16874 33881 16908 33915
rect 16681 33609 16715 33643
rect 15025 33473 15059 33507
rect 16865 33473 16899 33507
rect 14749 33405 14783 33439
rect 14933 33405 14967 33439
rect 17141 33405 17175 33439
rect 15393 33337 15427 33371
rect 16037 33269 16071 33303
rect 17049 33269 17083 33303
rect 17601 33269 17635 33303
rect 15577 33065 15611 33099
rect 14197 32929 14231 32963
rect 12909 32861 12943 32895
rect 16221 32861 16255 32895
rect 12664 32793 12698 32827
rect 16466 32793 16500 32827
rect 11529 32725 11563 32759
rect 14381 32725 14415 32759
rect 14473 32725 14507 32759
rect 14841 32725 14875 32759
rect 17601 32725 17635 32759
rect 14657 32385 14691 32419
rect 16681 32385 16715 32419
rect 15393 32249 15427 32283
rect 14841 32181 14875 32215
rect 16865 32181 16899 32215
rect 14473 31977 14507 32011
rect 15025 31977 15059 32011
rect 17233 31977 17267 32011
rect 17141 31841 17175 31875
rect 20177 31841 20211 31875
rect 9597 31773 9631 31807
rect 9853 31773 9887 31807
rect 15025 31773 15059 31807
rect 15209 31773 15243 31807
rect 15301 31773 15335 31807
rect 15761 31773 15795 31807
rect 17325 31773 17359 31807
rect 17417 31773 17451 31807
rect 17969 31773 18003 31807
rect 18061 31773 18095 31807
rect 18613 31773 18647 31807
rect 20049 31773 20083 31807
rect 20269 31773 20303 31807
rect 19533 31705 19567 31739
rect 20177 31705 20211 31739
rect 20453 31705 20487 31739
rect 10977 31637 11011 31671
rect 20913 31637 20947 31671
rect 16773 31433 16807 31467
rect 17969 31433 18003 31467
rect 19625 31433 19659 31467
rect 18245 31365 18279 31399
rect 1676 31297 1710 31331
rect 3249 31297 3283 31331
rect 8300 31297 8334 31331
rect 16957 31297 16991 31331
rect 17233 31297 17267 31331
rect 1409 31229 1443 31263
rect 8033 31229 8067 31263
rect 18061 31229 18095 31263
rect 18153 31229 18187 31263
rect 18337 31229 18371 31263
rect 18521 31229 18555 31263
rect 2789 31093 2823 31127
rect 9413 31093 9447 31127
rect 17141 31093 17175 31127
rect 19073 31093 19107 31127
rect 20085 30889 20119 30923
rect 14105 30753 14139 30787
rect 37841 30753 37875 30787
rect 9413 30685 9447 30719
rect 20361 30685 20395 30719
rect 20458 30685 20492 30719
rect 38117 30685 38151 30719
rect 14350 30617 14384 30651
rect 17877 30617 17911 30651
rect 20085 30617 20119 30651
rect 20269 30617 20303 30651
rect 21097 30617 21131 30651
rect 10701 30549 10735 30583
rect 15485 30549 15519 30583
rect 18337 30549 18371 30583
rect 9321 30345 9355 30379
rect 38117 30345 38151 30379
rect 16926 30277 16960 30311
rect 16681 30209 16715 30243
rect 18797 30209 18831 30243
rect 19073 30209 19107 30243
rect 18521 30141 18555 30175
rect 19349 30141 19383 30175
rect 18613 30073 18647 30107
rect 18061 30005 18095 30039
rect 19809 30005 19843 30039
rect 16681 29801 16715 29835
rect 18061 29733 18095 29767
rect 19441 29665 19475 29699
rect 19533 29665 19567 29699
rect 15301 29597 15335 29631
rect 15393 29597 15427 29631
rect 19349 29597 19383 29631
rect 19809 29597 19843 29631
rect 15209 29529 15243 29563
rect 15669 29529 15703 29563
rect 16129 29529 16163 29563
rect 19625 29529 19659 29563
rect 11253 29461 11287 29495
rect 15577 29461 15611 29495
rect 18613 29461 18647 29495
rect 19257 29461 19291 29495
rect 20361 29461 20395 29495
rect 8861 29257 8895 29291
rect 16957 29257 16991 29291
rect 7748 29189 7782 29223
rect 11897 29189 11931 29223
rect 12541 29189 12575 29223
rect 16037 29189 16071 29223
rect 17141 29189 17175 29223
rect 19809 29189 19843 29223
rect 16861 29155 16895 29189
rect 10977 29121 11011 29155
rect 11713 29121 11747 29155
rect 11989 29121 12023 29155
rect 13257 29121 13291 29155
rect 17233 29121 17267 29155
rect 19349 29121 19383 29155
rect 7481 29053 7515 29087
rect 13001 29053 13035 29087
rect 15485 29053 15519 29087
rect 17049 29053 17083 29087
rect 19073 29053 19107 29087
rect 11529 28985 11563 29019
rect 14381 28985 14415 29019
rect 19165 28985 19199 29019
rect 19257 28985 19291 29019
rect 12817 28713 12851 28747
rect 15853 28713 15887 28747
rect 18613 28713 18647 28747
rect 19257 28713 19291 28747
rect 7021 28509 7055 28543
rect 10425 28509 10459 28543
rect 12633 28509 12667 28543
rect 17233 28509 17267 28543
rect 19533 28509 19567 28543
rect 12173 28441 12207 28475
rect 16966 28441 17000 28475
rect 19257 28441 19291 28475
rect 5549 28373 5583 28407
rect 9873 28373 9907 28407
rect 19441 28373 19475 28407
rect 20269 28373 20303 28407
rect 3893 28169 3927 28203
rect 13645 28169 13679 28203
rect 18153 28169 18187 28203
rect 18245 28169 18279 28203
rect 21097 28169 21131 28203
rect 12510 28101 12544 28135
rect 14565 28101 14599 28135
rect 20545 28101 20579 28135
rect 2513 28033 2547 28067
rect 2780 28033 2814 28067
rect 9321 28033 9355 28067
rect 9781 28033 9815 28067
rect 10701 28033 10735 28067
rect 11805 28033 11839 28067
rect 14289 28033 14323 28067
rect 14657 28033 14691 28067
rect 15301 28033 15335 28067
rect 18061 28033 18095 28067
rect 18889 28033 18923 28067
rect 19901 28033 19935 28067
rect 19993 28033 20027 28067
rect 9873 27965 9907 27999
rect 10609 27965 10643 27999
rect 10793 27965 10827 27999
rect 10885 27965 10919 27999
rect 12265 27965 12299 27999
rect 14473 27965 14507 27999
rect 18429 27965 18463 27999
rect 18981 27965 19015 27999
rect 19533 27965 19567 27999
rect 19717 27965 19751 27999
rect 19809 27965 19843 27999
rect 10425 27897 10459 27931
rect 14289 27897 14323 27931
rect 17509 27897 17543 27931
rect 11713 27829 11747 27863
rect 15485 27829 15519 27863
rect 18337 27829 18371 27863
rect 20085 27829 20119 27863
rect 2789 27625 2823 27659
rect 18521 27625 18555 27659
rect 10517 27557 10551 27591
rect 11805 27557 11839 27591
rect 17325 27557 17359 27591
rect 18337 27557 18371 27591
rect 20913 27557 20947 27591
rect 21649 27557 21683 27591
rect 1409 27489 1443 27523
rect 9597 27489 9631 27523
rect 11253 27489 11287 27523
rect 20085 27489 20119 27523
rect 7665 27421 7699 27455
rect 9321 27421 9355 27455
rect 11437 27421 11471 27455
rect 13001 27421 13035 27455
rect 15945 27421 15979 27455
rect 19901 27421 19935 27455
rect 20177 27421 20211 27455
rect 1676 27353 1710 27387
rect 12909 27353 12943 27387
rect 16190 27353 16224 27387
rect 18489 27353 18523 27387
rect 18705 27353 18739 27387
rect 19717 27353 19751 27387
rect 20637 27353 20671 27387
rect 7481 27285 7515 27319
rect 8953 27285 8987 27319
rect 9413 27285 9447 27319
rect 11345 27285 11379 27319
rect 12265 27285 12299 27319
rect 14197 27285 14231 27319
rect 15209 27285 15243 27319
rect 17877 27285 17911 27319
rect 21097 27285 21131 27319
rect 9689 27081 9723 27115
rect 12357 27081 12391 27115
rect 14105 27081 14139 27115
rect 15761 27081 15795 27115
rect 18889 27081 18923 27115
rect 19073 27081 19107 27115
rect 19625 27081 19659 27115
rect 7932 27013 7966 27047
rect 11697 27013 11731 27047
rect 11897 27013 11931 27047
rect 18521 27013 18555 27047
rect 20821 27013 20855 27047
rect 22569 27013 22603 27047
rect 7665 26945 7699 26979
rect 9873 26945 9907 26979
rect 9965 26945 9999 26979
rect 10149 26945 10183 26979
rect 10333 26945 10367 26979
rect 12541 26945 12575 26979
rect 14013 26945 14047 26979
rect 14197 26945 14231 26979
rect 14933 26945 14967 26979
rect 15577 26945 15611 26979
rect 16681 26945 16715 26979
rect 16937 26945 16971 26979
rect 19809 26945 19843 26979
rect 22109 26945 22143 26979
rect 18705 26877 18739 26911
rect 18797 26877 18831 26911
rect 19165 26877 19199 26911
rect 19890 26877 19924 26911
rect 19993 26877 20027 26911
rect 20085 26877 20119 26911
rect 21833 26877 21867 26911
rect 9045 26809 9079 26843
rect 10057 26809 10091 26843
rect 15117 26809 15151 26843
rect 18061 26809 18095 26843
rect 21097 26809 21131 26843
rect 22017 26809 22051 26843
rect 11529 26741 11563 26775
rect 11713 26741 11747 26775
rect 13093 26741 13127 26775
rect 21281 26741 21315 26775
rect 21925 26741 21959 26775
rect 2789 26537 2823 26571
rect 8953 26537 8987 26571
rect 9873 26537 9907 26571
rect 11897 26537 11931 26571
rect 19533 26537 19567 26571
rect 20361 26537 20395 26571
rect 5365 26469 5399 26503
rect 15025 26469 15059 26503
rect 16129 26469 16163 26503
rect 18521 26469 18555 26503
rect 19717 26469 19751 26503
rect 1409 26401 1443 26435
rect 4077 26401 4111 26435
rect 11437 26401 11471 26435
rect 12909 26401 12943 26435
rect 14473 26401 14507 26435
rect 18061 26401 18095 26435
rect 21741 26401 21775 26435
rect 3801 26333 3835 26367
rect 9229 26333 9263 26367
rect 9689 26333 9723 26367
rect 12081 26333 12115 26367
rect 12265 26333 12299 26367
rect 12357 26333 12391 26367
rect 14841 26333 14875 26367
rect 20269 26333 20303 26367
rect 21373 26333 21407 26367
rect 21649 26333 21683 26367
rect 21925 26333 21959 26367
rect 22109 26333 22143 26367
rect 22661 26333 22695 26367
rect 19579 26299 19613 26333
rect 1676 26265 1710 26299
rect 8953 26265 8987 26299
rect 9137 26265 9171 26299
rect 10333 26265 10367 26299
rect 14749 26265 14783 26299
rect 17417 26265 17451 26299
rect 17969 26265 18003 26299
rect 19349 26265 19383 26299
rect 13553 26197 13587 26231
rect 14657 26197 14691 26231
rect 18061 26197 18095 26231
rect 22845 26197 22879 26231
rect 7849 25993 7883 26027
rect 13001 25993 13035 26027
rect 19073 25993 19107 26027
rect 20729 25993 20763 26027
rect 22201 25993 22235 26027
rect 8554 25925 8588 25959
rect 21189 25925 21223 25959
rect 7665 25857 7699 25891
rect 11621 25857 11655 25891
rect 11888 25857 11922 25891
rect 13824 25857 13858 25891
rect 13921 25857 13955 25891
rect 14013 25857 14047 25891
rect 14197 25857 14231 25891
rect 14749 25857 14783 25891
rect 15016 25857 15050 25891
rect 16865 25857 16899 25891
rect 17049 25857 17083 25891
rect 17785 25857 17819 25891
rect 21925 25857 21959 25891
rect 22109 25857 22143 25891
rect 8309 25789 8343 25823
rect 20085 25721 20119 25755
rect 9689 25653 9723 25687
rect 14197 25653 14231 25687
rect 16129 25653 16163 25687
rect 17049 25653 17083 25687
rect 22385 25653 22419 25687
rect 9413 25449 9447 25483
rect 11437 25449 11471 25483
rect 13093 25449 13127 25483
rect 14289 25449 14323 25483
rect 17877 25449 17911 25483
rect 21741 25449 21775 25483
rect 9321 25381 9355 25415
rect 20453 25381 20487 25415
rect 21005 25381 21039 25415
rect 9505 25313 9539 25347
rect 10425 25313 10459 25347
rect 10609 25313 10643 25347
rect 16313 25313 16347 25347
rect 19533 25313 19567 25347
rect 19901 25313 19935 25347
rect 9229 25245 9263 25279
rect 10701 25245 10735 25279
rect 11621 25245 11655 25279
rect 11713 25245 11747 25279
rect 13001 25245 13035 25279
rect 13277 25245 13311 25279
rect 15485 25245 15519 25279
rect 16037 25245 16071 25279
rect 16405 25245 16439 25279
rect 16957 25245 16991 25279
rect 17325 25245 17359 25279
rect 18017 25245 18051 25279
rect 18245 25245 18279 25279
rect 18383 25245 18417 25279
rect 18521 25245 18555 25279
rect 19625 25245 19659 25279
rect 19993 25245 20027 25279
rect 20729 25245 20763 25279
rect 10425 25177 10459 25211
rect 11437 25177 11471 25211
rect 12541 25177 12575 25211
rect 13185 25177 13219 25211
rect 18153 25177 18187 25211
rect 20821 25177 20855 25211
rect 19349 25109 19383 25143
rect 19717 25109 19751 25143
rect 20637 25109 20671 25143
rect 9597 24905 9631 24939
rect 12357 24905 12391 24939
rect 18061 24905 18095 24939
rect 24225 24905 24259 24939
rect 13921 24837 13955 24871
rect 19533 24837 19567 24871
rect 20177 24837 20211 24871
rect 13691 24803 13725 24837
rect 11713 24769 11747 24803
rect 12265 24769 12299 24803
rect 12541 24769 12575 24803
rect 16681 24769 16715 24803
rect 16948 24769 16982 24803
rect 19441 24769 19475 24803
rect 19717 24769 19751 24803
rect 20361 24769 20395 24803
rect 20913 24769 20947 24803
rect 23673 24769 23707 24803
rect 23764 24769 23798 24803
rect 24225 24769 24259 24803
rect 24409 24769 24443 24803
rect 21097 24701 21131 24735
rect 22937 24701 22971 24735
rect 23489 24701 23523 24735
rect 13553 24633 13587 24667
rect 19717 24633 19751 24667
rect 12725 24565 12759 24599
rect 13737 24565 13771 24599
rect 14381 24565 14415 24599
rect 18981 24565 19015 24599
rect 22017 24565 22051 24599
rect 23581 24565 23615 24599
rect 13553 24361 13587 24395
rect 14105 24361 14139 24395
rect 16957 24361 16991 24395
rect 18245 24361 18279 24395
rect 18429 24361 18463 24395
rect 20085 24361 20119 24395
rect 20821 24361 20855 24395
rect 23397 24361 23431 24395
rect 12449 24293 12483 24327
rect 20177 24293 20211 24327
rect 21557 24293 21591 24327
rect 22385 24293 22419 24327
rect 22569 24293 22603 24327
rect 23489 24293 23523 24327
rect 14289 24225 14323 24259
rect 15209 24225 15243 24259
rect 19993 24225 20027 24259
rect 22109 24225 22143 24259
rect 23397 24225 23431 24259
rect 12909 24157 12943 24191
rect 13093 24157 13127 24191
rect 13185 24157 13219 24191
rect 13323 24157 13357 24191
rect 14381 24157 14415 24191
rect 14473 24157 14507 24191
rect 14565 24157 14599 24191
rect 16865 24157 16899 24191
rect 17141 24157 17175 24191
rect 20269 24157 20303 24191
rect 23581 24157 23615 24191
rect 18613 24089 18647 24123
rect 23213 24089 23247 24123
rect 18413 24021 18447 24055
rect 19349 24021 19383 24055
rect 24409 24021 24443 24055
rect 13277 23817 13311 23851
rect 15209 23817 15243 23851
rect 16773 23817 16807 23851
rect 17785 23817 17819 23851
rect 19533 23817 19567 23851
rect 20545 23817 20579 23851
rect 21925 23817 21959 23851
rect 18245 23749 18279 23783
rect 13001 23681 13035 23715
rect 13185 23681 13219 23715
rect 13277 23681 13311 23715
rect 13737 23681 13771 23715
rect 13921 23681 13955 23715
rect 15025 23681 15059 23715
rect 16957 23681 16991 23715
rect 17601 23681 17635 23715
rect 17785 23681 17819 23715
rect 21281 23681 21315 23715
rect 22017 23681 22051 23715
rect 22293 23681 22327 23715
rect 22569 23681 22603 23715
rect 23305 23681 23339 23715
rect 23397 23681 23431 23715
rect 23673 23681 23707 23715
rect 24133 23681 24167 23715
rect 24317 23681 24351 23715
rect 14841 23613 14875 23647
rect 21833 23613 21867 23647
rect 12541 23545 12575 23579
rect 14013 23545 14047 23579
rect 23581 23545 23615 23579
rect 24317 23545 24351 23579
rect 15761 23477 15795 23511
rect 23121 23477 23155 23511
rect 24593 23477 24627 23511
rect 12725 23273 12759 23307
rect 15117 23273 15151 23307
rect 15761 23273 15795 23307
rect 16773 23273 16807 23307
rect 17969 23273 18003 23307
rect 19349 23273 19383 23307
rect 20545 23273 20579 23307
rect 21649 23273 21683 23307
rect 23213 23273 23247 23307
rect 13369 23205 13403 23239
rect 15301 23205 15335 23239
rect 17325 23205 17359 23239
rect 17785 23205 17819 23239
rect 22201 23205 22235 23239
rect 23029 23205 23063 23239
rect 23673 23205 23707 23239
rect 15945 23137 15979 23171
rect 16129 23137 16163 23171
rect 22753 23137 22787 23171
rect 16037 23069 16071 23103
rect 16221 23069 16255 23103
rect 16957 23069 16991 23103
rect 19257 23069 19291 23103
rect 20545 23069 20579 23103
rect 20723 23069 20757 23103
rect 21557 23069 21591 23103
rect 24409 23069 24443 23103
rect 14933 23001 14967 23035
rect 17049 23001 17083 23035
rect 17953 23001 17987 23035
rect 18153 23001 18187 23035
rect 15133 22933 15167 22967
rect 17141 22933 17175 22967
rect 18705 22933 18739 22967
rect 19717 22933 19751 22967
rect 14841 22729 14875 22763
rect 15485 22729 15519 22763
rect 15761 22729 15795 22763
rect 17141 22729 17175 22763
rect 17417 22729 17451 22763
rect 17877 22729 17911 22763
rect 22017 22729 22051 22763
rect 23857 22729 23891 22763
rect 14841 22593 14875 22627
rect 15025 22593 15059 22627
rect 15485 22593 15519 22627
rect 15649 22593 15683 22627
rect 15853 22593 15887 22627
rect 17049 22593 17083 22627
rect 17263 22593 17297 22627
rect 18061 22593 18095 22627
rect 18245 22593 18279 22627
rect 18337 22593 18371 22627
rect 19993 22593 20027 22627
rect 20269 22593 20303 22627
rect 21097 22593 21131 22627
rect 21281 22593 21315 22627
rect 21833 22593 21867 22627
rect 22109 22593 22143 22627
rect 22293 22593 22327 22627
rect 17417 22525 17451 22559
rect 18153 22525 18187 22559
rect 18889 22525 18923 22559
rect 22753 22525 22787 22559
rect 19257 22457 19291 22491
rect 19349 22457 19383 22491
rect 19809 22389 19843 22423
rect 20177 22389 20211 22423
rect 21189 22389 21223 22423
rect 23305 22389 23339 22423
rect 16681 22185 16715 22219
rect 17877 22185 17911 22219
rect 17969 22117 18003 22151
rect 22753 22049 22787 22083
rect 17509 21981 17543 22015
rect 18061 21981 18095 22015
rect 18705 21981 18739 22015
rect 19901 21981 19935 22015
rect 20545 21981 20579 22015
rect 20913 21981 20947 22015
rect 21649 21981 21683 22015
rect 21879 21981 21913 22015
rect 22017 21981 22051 22015
rect 22661 21981 22695 22015
rect 22845 21981 22879 22015
rect 23305 21981 23339 22015
rect 19809 21913 19843 21947
rect 23397 21913 23431 21947
rect 17601 21845 17635 21879
rect 21741 21845 21775 21879
rect 18245 21641 18279 21675
rect 18797 21641 18831 21675
rect 19809 21641 19843 21675
rect 20729 21641 20763 21675
rect 23765 21641 23799 21675
rect 19717 21505 19751 21539
rect 20085 21505 20119 21539
rect 20269 21505 20303 21539
rect 20913 21505 20947 21539
rect 21097 21505 21131 21539
rect 21189 21505 21223 21539
rect 22109 21505 22143 21539
rect 22661 21505 22695 21539
rect 22937 21505 22971 21539
rect 21833 21437 21867 21471
rect 22385 21437 22419 21471
rect 20085 21369 20119 21403
rect 21557 21097 21591 21131
rect 22201 21097 22235 21131
rect 19441 21029 19475 21063
rect 20545 21029 20579 21063
rect 19579 20961 19613 20995
rect 18705 20893 18739 20927
rect 19349 20893 19383 20927
rect 19717 20893 19751 20927
rect 21465 20893 21499 20927
rect 22109 20893 22143 20927
rect 22293 20893 22327 20927
rect 22753 20825 22787 20859
rect 19165 20553 19199 20587
rect 20453 20553 20487 20587
rect 21833 20553 21867 20587
rect 22385 20553 22419 20587
rect 1593 18377 1627 18411
rect 1409 18241 1443 18275
rect 2053 18241 2087 18275
rect 37289 12801 37323 12835
rect 37841 12801 37875 12835
rect 38025 12597 38059 12631
rect 38117 12325 38151 12359
rect 37933 12189 37967 12223
rect 1409 2805 1443 2839
rect 34897 2805 34931 2839
rect 16865 2601 16899 2635
rect 1409 2465 1443 2499
rect 1685 2465 1719 2499
rect 35081 2465 35115 2499
rect 17049 2397 17083 2431
rect 17509 2397 17543 2431
rect 35265 2329 35299 2363
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 30561 37451 30619 37457
rect 30561 37417 30573 37451
rect 30607 37448 30619 37451
rect 30926 37448 30932 37460
rect 30607 37420 30932 37448
rect 30607 37417 30619 37420
rect 30561 37411 30619 37417
rect 30926 37408 30932 37420
rect 30984 37408 30990 37460
rect 14737 37315 14795 37321
rect 14737 37281 14749 37315
rect 14783 37312 14795 37315
rect 17770 37312 17776 37324
rect 14783 37284 17776 37312
rect 14783 37281 14795 37284
rect 14737 37275 14795 37281
rect 17770 37272 17776 37284
rect 17828 37272 17834 37324
rect 13538 37204 13544 37256
rect 13596 37244 13602 37256
rect 14274 37244 14280 37256
rect 13596 37216 14280 37244
rect 13596 37204 13602 37216
rect 14274 37204 14280 37216
rect 14332 37244 14338 37256
rect 14553 37247 14611 37253
rect 14553 37244 14565 37247
rect 14332 37216 14565 37244
rect 14332 37204 14338 37216
rect 14553 37213 14565 37216
rect 14599 37213 14611 37247
rect 14553 37207 14611 37213
rect 30926 37204 30932 37256
rect 30984 37244 30990 37256
rect 31205 37247 31263 37253
rect 31205 37244 31217 37247
rect 30984 37216 31217 37244
rect 30984 37204 30990 37216
rect 31205 37213 31217 37216
rect 31251 37213 31263 37247
rect 31205 37207 31263 37213
rect 31018 37108 31024 37120
rect 30979 37080 31024 37108
rect 31018 37068 31024 37080
rect 31076 37068 31082 37120
rect 1104 37018 38824 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 38824 37018
rect 1104 36944 38824 36966
rect 14274 36904 14280 36916
rect 14235 36876 14280 36904
rect 14274 36864 14280 36876
rect 14332 36864 14338 36916
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 3418 35980 3424 36032
rect 3476 36020 3482 36032
rect 9398 36020 9404 36032
rect 3476 35992 9404 36020
rect 3476 35980 3482 35992
rect 9398 35980 9404 35992
rect 9456 35980 9462 36032
rect 1104 35930 38824 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 38824 35930
rect 1104 35856 38824 35878
rect 8294 35748 8300 35760
rect 6380 35720 8300 35748
rect 6380 35689 6408 35720
rect 8294 35708 8300 35720
rect 8352 35708 8358 35760
rect 6638 35689 6644 35692
rect 6365 35683 6423 35689
rect 6365 35649 6377 35683
rect 6411 35649 6423 35683
rect 6365 35643 6423 35649
rect 6632 35643 6644 35689
rect 6696 35680 6702 35692
rect 8312 35680 8340 35708
rect 8757 35683 8815 35689
rect 8757 35680 8769 35683
rect 6696 35652 6732 35680
rect 8312 35652 8769 35680
rect 6638 35640 6644 35643
rect 6696 35640 6702 35652
rect 8757 35649 8769 35652
rect 8803 35649 8815 35683
rect 8757 35643 8815 35649
rect 9024 35683 9082 35689
rect 9024 35649 9036 35683
rect 9070 35680 9082 35683
rect 17218 35680 17224 35692
rect 9070 35652 17224 35680
rect 9070 35649 9082 35652
rect 9024 35643 9082 35649
rect 17218 35640 17224 35652
rect 17276 35640 17282 35692
rect 18782 35544 18788 35556
rect 10060 35516 18788 35544
rect 7745 35479 7803 35485
rect 7745 35445 7757 35479
rect 7791 35476 7803 35479
rect 10060 35476 10088 35516
rect 18782 35504 18788 35516
rect 18840 35504 18846 35556
rect 7791 35448 10088 35476
rect 10137 35479 10195 35485
rect 7791 35445 7803 35448
rect 7745 35439 7803 35445
rect 10137 35445 10149 35479
rect 10183 35476 10195 35479
rect 17678 35476 17684 35488
rect 10183 35448 17684 35476
rect 10183 35445 10195 35448
rect 10137 35439 10195 35445
rect 17678 35436 17684 35448
rect 17736 35436 17742 35488
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 17126 35028 17132 35080
rect 17184 35068 17190 35080
rect 17221 35071 17279 35077
rect 17221 35068 17233 35071
rect 17184 35040 17233 35068
rect 17184 35028 17190 35040
rect 17221 35037 17233 35040
rect 17267 35037 17279 35071
rect 17221 35031 17279 35037
rect 16758 34960 16764 35012
rect 16816 35000 16822 35012
rect 16954 35003 17012 35009
rect 16954 35000 16966 35003
rect 16816 34972 16966 35000
rect 16816 34960 16822 34972
rect 16954 34969 16966 34972
rect 17000 34969 17012 35003
rect 16954 34963 17012 34969
rect 15841 34935 15899 34941
rect 15841 34901 15853 34935
rect 15887 34932 15899 34935
rect 17126 34932 17132 34944
rect 15887 34904 17132 34932
rect 15887 34901 15899 34904
rect 15841 34895 15899 34901
rect 17126 34892 17132 34904
rect 17184 34892 17190 34944
rect 1104 34842 38824 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 38824 34842
rect 1104 34768 38824 34790
rect 18049 34731 18107 34737
rect 18049 34697 18061 34731
rect 18095 34728 18107 34731
rect 18874 34728 18880 34740
rect 18095 34700 18880 34728
rect 18095 34697 18107 34700
rect 18049 34691 18107 34697
rect 18874 34688 18880 34700
rect 18932 34688 18938 34740
rect 16942 34601 16948 34604
rect 16936 34555 16948 34601
rect 17000 34592 17006 34604
rect 17000 34564 17036 34592
rect 16942 34552 16948 34555
rect 17000 34552 17006 34564
rect 16669 34527 16727 34533
rect 16669 34493 16681 34527
rect 16715 34493 16727 34527
rect 16669 34487 16727 34493
rect 16684 34388 16712 34487
rect 17034 34388 17040 34400
rect 16684 34360 17040 34388
rect 17034 34348 17040 34360
rect 17092 34348 17098 34400
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 15749 34187 15807 34193
rect 15749 34153 15761 34187
rect 15795 34184 15807 34187
rect 17310 34184 17316 34196
rect 15795 34156 17316 34184
rect 15795 34153 15807 34156
rect 15749 34147 15807 34153
rect 17310 34144 17316 34156
rect 17368 34144 17374 34196
rect 17034 33940 17040 33992
rect 17092 33980 17098 33992
rect 17129 33983 17187 33989
rect 17129 33980 17141 33983
rect 17092 33952 17141 33980
rect 17092 33940 17098 33952
rect 17129 33949 17141 33952
rect 17175 33949 17187 33983
rect 17129 33943 17187 33949
rect 16666 33872 16672 33924
rect 16724 33912 16730 33924
rect 16862 33915 16920 33921
rect 16862 33912 16874 33915
rect 16724 33884 16874 33912
rect 16724 33872 16730 33884
rect 16862 33881 16874 33884
rect 16908 33881 16920 33915
rect 16862 33875 16920 33881
rect 15838 33804 15844 33856
rect 15896 33844 15902 33856
rect 31018 33844 31024 33856
rect 15896 33816 31024 33844
rect 15896 33804 15902 33816
rect 31018 33804 31024 33816
rect 31076 33804 31082 33856
rect 1104 33754 38824 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 38824 33754
rect 1104 33680 38824 33702
rect 16666 33640 16672 33652
rect 16627 33612 16672 33640
rect 16666 33600 16672 33612
rect 16724 33600 16730 33652
rect 15013 33507 15071 33513
rect 15013 33473 15025 33507
rect 15059 33504 15071 33507
rect 16482 33504 16488 33516
rect 15059 33476 16488 33504
rect 15059 33473 15071 33476
rect 15013 33467 15071 33473
rect 16482 33464 16488 33476
rect 16540 33464 16546 33516
rect 16853 33507 16911 33513
rect 16853 33473 16865 33507
rect 16899 33504 16911 33507
rect 18138 33504 18144 33516
rect 16899 33476 18144 33504
rect 16899 33473 16911 33476
rect 16853 33467 16911 33473
rect 18138 33464 18144 33476
rect 18196 33464 18202 33516
rect 14182 33396 14188 33448
rect 14240 33436 14246 33448
rect 14737 33439 14795 33445
rect 14737 33436 14749 33439
rect 14240 33408 14749 33436
rect 14240 33396 14246 33408
rect 14737 33405 14749 33408
rect 14783 33405 14795 33439
rect 14737 33399 14795 33405
rect 14921 33439 14979 33445
rect 14921 33405 14933 33439
rect 14967 33436 14979 33439
rect 15838 33436 15844 33448
rect 14967 33408 15844 33436
rect 14967 33405 14979 33408
rect 14921 33399 14979 33405
rect 15838 33396 15844 33408
rect 15896 33396 15902 33448
rect 16022 33396 16028 33448
rect 16080 33436 16086 33448
rect 17129 33439 17187 33445
rect 17129 33436 17141 33439
rect 16080 33408 17141 33436
rect 16080 33396 16086 33408
rect 17129 33405 17141 33408
rect 17175 33436 17187 33439
rect 17954 33436 17960 33448
rect 17175 33408 17960 33436
rect 17175 33405 17187 33408
rect 17129 33399 17187 33405
rect 17954 33396 17960 33408
rect 18012 33396 18018 33448
rect 15381 33371 15439 33377
rect 15381 33337 15393 33371
rect 15427 33368 15439 33371
rect 16666 33368 16672 33380
rect 15427 33340 16672 33368
rect 15427 33337 15439 33340
rect 15381 33331 15439 33337
rect 16666 33328 16672 33340
rect 16724 33328 16730 33380
rect 15102 33260 15108 33312
rect 15160 33300 15166 33312
rect 16022 33300 16028 33312
rect 15160 33272 16028 33300
rect 15160 33260 15166 33272
rect 16022 33260 16028 33272
rect 16080 33260 16086 33312
rect 17037 33303 17095 33309
rect 17037 33269 17049 33303
rect 17083 33300 17095 33303
rect 17310 33300 17316 33312
rect 17083 33272 17316 33300
rect 17083 33269 17095 33272
rect 17037 33263 17095 33269
rect 17310 33260 17316 33272
rect 17368 33300 17374 33312
rect 17589 33303 17647 33309
rect 17589 33300 17601 33303
rect 17368 33272 17601 33300
rect 17368 33260 17374 33272
rect 17589 33269 17601 33272
rect 17635 33269 17647 33303
rect 17589 33263 17647 33269
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 15565 33099 15623 33105
rect 15565 33065 15577 33099
rect 15611 33096 15623 33099
rect 15838 33096 15844 33108
rect 15611 33068 15844 33096
rect 15611 33065 15623 33068
rect 15565 33059 15623 33065
rect 15838 33056 15844 33068
rect 15896 33056 15902 33108
rect 14182 32960 14188 32972
rect 14143 32932 14188 32960
rect 14182 32920 14188 32932
rect 14240 32920 14246 32972
rect 12897 32895 12955 32901
rect 12897 32861 12909 32895
rect 12943 32892 12955 32895
rect 13814 32892 13820 32904
rect 12943 32864 13820 32892
rect 12943 32861 12955 32864
rect 12897 32855 12955 32861
rect 13814 32852 13820 32864
rect 13872 32892 13878 32904
rect 16209 32895 16267 32901
rect 16209 32892 16221 32895
rect 13872 32864 16221 32892
rect 13872 32852 13878 32864
rect 16209 32861 16221 32864
rect 16255 32892 16267 32895
rect 17034 32892 17040 32904
rect 16255 32864 17040 32892
rect 16255 32861 16267 32864
rect 16209 32855 16267 32861
rect 17034 32852 17040 32864
rect 17092 32852 17098 32904
rect 12652 32827 12710 32833
rect 12652 32793 12664 32827
rect 12698 32824 12710 32827
rect 15010 32824 15016 32836
rect 12698 32796 15016 32824
rect 12698 32793 12710 32796
rect 12652 32787 12710 32793
rect 15010 32784 15016 32796
rect 15068 32784 15074 32836
rect 15930 32784 15936 32836
rect 15988 32824 15994 32836
rect 16454 32827 16512 32833
rect 16454 32824 16466 32827
rect 15988 32796 16466 32824
rect 15988 32784 15994 32796
rect 16454 32793 16466 32796
rect 16500 32793 16512 32827
rect 16454 32787 16512 32793
rect 11514 32756 11520 32768
rect 11475 32728 11520 32756
rect 11514 32716 11520 32728
rect 11572 32716 11578 32768
rect 14366 32756 14372 32768
rect 14327 32728 14372 32756
rect 14366 32716 14372 32728
rect 14424 32716 14430 32768
rect 14458 32716 14464 32768
rect 14516 32756 14522 32768
rect 14516 32728 14561 32756
rect 14516 32716 14522 32728
rect 14642 32716 14648 32768
rect 14700 32756 14706 32768
rect 14829 32759 14887 32765
rect 14829 32756 14841 32759
rect 14700 32728 14841 32756
rect 14700 32716 14706 32728
rect 14829 32725 14841 32728
rect 14875 32725 14887 32759
rect 17586 32756 17592 32768
rect 17547 32728 17592 32756
rect 14829 32719 14887 32725
rect 17586 32716 17592 32728
rect 17644 32716 17650 32768
rect 1104 32666 38824 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 38824 32666
rect 1104 32592 38824 32614
rect 14642 32416 14648 32428
rect 14603 32388 14648 32416
rect 14642 32376 14648 32388
rect 14700 32376 14706 32428
rect 16666 32416 16672 32428
rect 16627 32388 16672 32416
rect 16666 32376 16672 32388
rect 16724 32376 16730 32428
rect 15746 32308 15752 32360
rect 15804 32348 15810 32360
rect 18230 32348 18236 32360
rect 15804 32320 18236 32348
rect 15804 32308 15810 32320
rect 18230 32308 18236 32320
rect 18288 32308 18294 32360
rect 14366 32240 14372 32292
rect 14424 32280 14430 32292
rect 15381 32283 15439 32289
rect 15381 32280 15393 32283
rect 14424 32252 15393 32280
rect 14424 32240 14430 32252
rect 15381 32249 15393 32252
rect 15427 32280 15439 32283
rect 15427 32252 26234 32280
rect 15427 32249 15439 32252
rect 15381 32243 15439 32249
rect 14829 32215 14887 32221
rect 14829 32181 14841 32215
rect 14875 32212 14887 32215
rect 14918 32212 14924 32224
rect 14875 32184 14924 32212
rect 14875 32181 14887 32184
rect 14829 32175 14887 32181
rect 14918 32172 14924 32184
rect 14976 32172 14982 32224
rect 16850 32212 16856 32224
rect 16811 32184 16856 32212
rect 16850 32172 16856 32184
rect 16908 32172 16914 32224
rect 17678 32172 17684 32224
rect 17736 32212 17742 32224
rect 21634 32212 21640 32224
rect 17736 32184 21640 32212
rect 17736 32172 17742 32184
rect 21634 32172 21640 32184
rect 21692 32172 21698 32224
rect 26206 32212 26234 32252
rect 37826 32212 37832 32224
rect 26206 32184 37832 32212
rect 37826 32172 37832 32184
rect 37884 32172 37890 32224
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 11514 31968 11520 32020
rect 11572 32008 11578 32020
rect 14461 32011 14519 32017
rect 14461 32008 14473 32011
rect 11572 31980 14473 32008
rect 11572 31968 11578 31980
rect 14461 31977 14473 31980
rect 14507 31977 14519 32011
rect 15010 32008 15016 32020
rect 14971 31980 15016 32008
rect 14461 31971 14519 31977
rect 9585 31807 9643 31813
rect 9585 31773 9597 31807
rect 9631 31773 9643 31807
rect 9585 31767 9643 31773
rect 8294 31696 8300 31748
rect 8352 31736 8358 31748
rect 9600 31736 9628 31767
rect 9674 31764 9680 31816
rect 9732 31804 9738 31816
rect 9841 31807 9899 31813
rect 9841 31804 9853 31807
rect 9732 31776 9853 31804
rect 9732 31764 9738 31776
rect 9841 31773 9853 31776
rect 9887 31773 9899 31807
rect 14476 31804 14504 31971
rect 15010 31968 15016 31980
rect 15068 31968 15074 32020
rect 17218 32008 17224 32020
rect 17179 31980 17224 32008
rect 17218 31968 17224 31980
rect 17276 31968 17282 32020
rect 17310 31968 17316 32020
rect 17368 32008 17374 32020
rect 19426 32008 19432 32020
rect 17368 31980 19432 32008
rect 17368 31968 17374 31980
rect 19426 31968 19432 31980
rect 19484 31968 19490 32020
rect 17954 31900 17960 31952
rect 18012 31940 18018 31952
rect 19518 31940 19524 31952
rect 18012 31912 19524 31940
rect 18012 31900 18018 31912
rect 19518 31900 19524 31912
rect 19576 31900 19582 31952
rect 15562 31872 15568 31884
rect 15212 31844 15568 31872
rect 15013 31807 15071 31813
rect 15013 31804 15025 31807
rect 14476 31776 15025 31804
rect 9841 31767 9899 31773
rect 15013 31773 15025 31776
rect 15059 31804 15071 31807
rect 15102 31804 15108 31816
rect 15059 31776 15108 31804
rect 15059 31773 15071 31776
rect 15013 31767 15071 31773
rect 15102 31764 15108 31776
rect 15160 31764 15166 31816
rect 15212 31813 15240 31844
rect 15562 31832 15568 31844
rect 15620 31872 15626 31884
rect 17129 31875 17187 31881
rect 15620 31844 16528 31872
rect 15620 31832 15626 31844
rect 15197 31807 15255 31813
rect 15197 31773 15209 31807
rect 15243 31773 15255 31807
rect 15197 31767 15255 31773
rect 15289 31807 15347 31813
rect 15289 31773 15301 31807
rect 15335 31804 15347 31807
rect 15746 31804 15752 31816
rect 15335 31776 15752 31804
rect 15335 31773 15347 31776
rect 15289 31767 15347 31773
rect 15746 31764 15752 31776
rect 15804 31764 15810 31816
rect 8352 31708 9628 31736
rect 15120 31736 15148 31764
rect 16298 31736 16304 31748
rect 15120 31708 16304 31736
rect 8352 31696 8358 31708
rect 16298 31696 16304 31708
rect 16356 31696 16362 31748
rect 10962 31668 10968 31680
rect 10923 31640 10968 31668
rect 10962 31628 10968 31640
rect 11020 31628 11026 31680
rect 16500 31668 16528 31844
rect 17129 31841 17141 31875
rect 17175 31872 17187 31875
rect 17218 31872 17224 31884
rect 17175 31844 17224 31872
rect 17175 31841 17187 31844
rect 17129 31835 17187 31841
rect 17218 31832 17224 31844
rect 17276 31832 17282 31884
rect 17678 31832 17684 31884
rect 17736 31872 17742 31884
rect 17736 31844 18092 31872
rect 17736 31832 17742 31844
rect 18064 31813 18092 31844
rect 18138 31832 18144 31884
rect 18196 31872 18202 31884
rect 20165 31875 20223 31881
rect 20165 31872 20177 31875
rect 18196 31844 20177 31872
rect 18196 31832 18202 31844
rect 20165 31841 20177 31844
rect 20211 31841 20223 31875
rect 20165 31835 20223 31841
rect 17313 31807 17371 31813
rect 17313 31773 17325 31807
rect 17359 31773 17371 31807
rect 17313 31767 17371 31773
rect 17405 31807 17463 31813
rect 17405 31773 17417 31807
rect 17451 31804 17463 31807
rect 17957 31807 18015 31813
rect 17957 31804 17969 31807
rect 17451 31776 17969 31804
rect 17451 31773 17463 31776
rect 17405 31767 17463 31773
rect 17957 31773 17969 31776
rect 18003 31773 18015 31807
rect 17957 31767 18015 31773
rect 18049 31807 18107 31813
rect 18049 31773 18061 31807
rect 18095 31804 18107 31807
rect 18601 31807 18659 31813
rect 18601 31804 18613 31807
rect 18095 31776 18613 31804
rect 18095 31773 18107 31776
rect 18049 31767 18107 31773
rect 18601 31773 18613 31776
rect 18647 31773 18659 31807
rect 18601 31767 18659 31773
rect 17328 31736 17356 31767
rect 19426 31764 19432 31816
rect 19484 31804 19490 31816
rect 20037 31807 20095 31813
rect 20037 31804 20049 31807
rect 19484 31776 20049 31804
rect 19484 31764 19490 31776
rect 20037 31773 20049 31776
rect 20083 31773 20095 31807
rect 20037 31767 20095 31773
rect 20254 31764 20260 31816
rect 20312 31804 20318 31816
rect 20312 31776 20357 31804
rect 20312 31764 20318 31776
rect 19334 31736 19340 31748
rect 17328 31708 19340 31736
rect 19334 31696 19340 31708
rect 19392 31696 19398 31748
rect 19518 31696 19524 31748
rect 19576 31736 19582 31748
rect 20165 31739 20223 31745
rect 20165 31736 20177 31739
rect 19576 31708 20177 31736
rect 19576 31696 19582 31708
rect 20165 31705 20177 31708
rect 20211 31705 20223 31739
rect 20165 31699 20223 31705
rect 20441 31739 20499 31745
rect 20441 31705 20453 31739
rect 20487 31705 20499 31739
rect 20441 31699 20499 31705
rect 18506 31668 18512 31680
rect 16500 31640 18512 31668
rect 18506 31628 18512 31640
rect 18564 31628 18570 31680
rect 20456 31668 20484 31699
rect 20622 31668 20628 31680
rect 20456 31640 20628 31668
rect 20622 31628 20628 31640
rect 20680 31668 20686 31680
rect 20901 31671 20959 31677
rect 20901 31668 20913 31671
rect 20680 31640 20913 31668
rect 20680 31628 20686 31640
rect 20901 31637 20913 31640
rect 20947 31637 20959 31671
rect 20901 31631 20959 31637
rect 1104 31578 38824 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 38824 31578
rect 1104 31504 38824 31526
rect 8294 31464 8300 31476
rect 8036 31436 8300 31464
rect 1670 31337 1676 31340
rect 1664 31328 1676 31337
rect 1631 31300 1676 31328
rect 1664 31291 1676 31300
rect 1728 31328 1734 31340
rect 3237 31331 3295 31337
rect 3237 31328 3249 31331
rect 1728 31300 3249 31328
rect 1670 31288 1676 31291
rect 1728 31288 1734 31300
rect 3237 31297 3249 31300
rect 3283 31297 3295 31331
rect 3237 31291 3295 31297
rect 1394 31260 1400 31272
rect 1355 31232 1400 31260
rect 1394 31220 1400 31232
rect 1452 31220 1458 31272
rect 7466 31220 7472 31272
rect 7524 31260 7530 31272
rect 8036 31269 8064 31436
rect 8294 31424 8300 31436
rect 8352 31424 8358 31476
rect 16758 31464 16764 31476
rect 16719 31436 16764 31464
rect 16758 31424 16764 31436
rect 16816 31424 16822 31476
rect 17218 31424 17224 31476
rect 17276 31464 17282 31476
rect 17957 31467 18015 31473
rect 17957 31464 17969 31467
rect 17276 31436 17969 31464
rect 17276 31424 17282 31436
rect 17957 31433 17969 31436
rect 18003 31433 18015 31467
rect 17957 31427 18015 31433
rect 19426 31424 19432 31476
rect 19484 31464 19490 31476
rect 19613 31467 19671 31473
rect 19613 31464 19625 31467
rect 19484 31436 19625 31464
rect 19484 31424 19490 31436
rect 19613 31433 19625 31436
rect 19659 31433 19671 31467
rect 19613 31427 19671 31433
rect 18233 31399 18291 31405
rect 18233 31365 18245 31399
rect 18279 31396 18291 31399
rect 18322 31396 18328 31408
rect 18279 31368 18328 31396
rect 18279 31365 18291 31368
rect 18233 31359 18291 31365
rect 18322 31356 18328 31368
rect 18380 31356 18386 31408
rect 8294 31337 8300 31340
rect 8288 31328 8300 31337
rect 8255 31300 8300 31328
rect 8288 31291 8300 31300
rect 8294 31288 8300 31291
rect 8352 31288 8358 31340
rect 16942 31328 16948 31340
rect 16903 31300 16948 31328
rect 16942 31288 16948 31300
rect 17000 31288 17006 31340
rect 17126 31288 17132 31340
rect 17184 31328 17190 31340
rect 17221 31331 17279 31337
rect 17221 31328 17233 31331
rect 17184 31300 17233 31328
rect 17184 31288 17190 31300
rect 17221 31297 17233 31300
rect 17267 31297 17279 31331
rect 17221 31291 17279 31297
rect 8021 31263 8079 31269
rect 8021 31260 8033 31263
rect 7524 31232 8033 31260
rect 7524 31220 7530 31232
rect 8021 31229 8033 31232
rect 8067 31229 8079 31263
rect 8021 31223 8079 31229
rect 17770 31220 17776 31272
rect 17828 31260 17834 31272
rect 18046 31260 18052 31272
rect 17828 31232 18052 31260
rect 17828 31220 17834 31232
rect 18046 31220 18052 31232
rect 18104 31220 18110 31272
rect 18141 31263 18199 31269
rect 18141 31229 18153 31263
rect 18187 31229 18199 31263
rect 18141 31223 18199 31229
rect 16482 31152 16488 31204
rect 16540 31192 16546 31204
rect 18156 31192 18184 31223
rect 18230 31220 18236 31272
rect 18288 31260 18294 31272
rect 18325 31263 18383 31269
rect 18325 31260 18337 31263
rect 18288 31232 18337 31260
rect 18288 31220 18294 31232
rect 18325 31229 18337 31232
rect 18371 31229 18383 31263
rect 18325 31223 18383 31229
rect 16540 31164 18184 31192
rect 18340 31192 18368 31223
rect 18506 31220 18512 31272
rect 18564 31260 18570 31272
rect 20070 31260 20076 31272
rect 18564 31232 20076 31260
rect 18564 31220 18570 31232
rect 20070 31220 20076 31232
rect 20128 31220 20134 31272
rect 18340 31164 19104 31192
rect 16540 31152 16546 31164
rect 2774 31084 2780 31136
rect 2832 31124 2838 31136
rect 9401 31127 9459 31133
rect 2832 31096 2877 31124
rect 2832 31084 2838 31096
rect 9401 31093 9413 31127
rect 9447 31124 9459 31127
rect 9766 31124 9772 31136
rect 9447 31096 9772 31124
rect 9447 31093 9459 31096
rect 9401 31087 9459 31093
rect 9766 31084 9772 31096
rect 9824 31084 9830 31136
rect 17129 31127 17187 31133
rect 17129 31093 17141 31127
rect 17175 31124 17187 31127
rect 17954 31124 17960 31136
rect 17175 31096 17960 31124
rect 17175 31093 17187 31096
rect 17129 31087 17187 31093
rect 17954 31084 17960 31096
rect 18012 31084 18018 31136
rect 19076 31133 19104 31164
rect 19061 31127 19119 31133
rect 19061 31093 19073 31127
rect 19107 31124 19119 31127
rect 20254 31124 20260 31136
rect 19107 31096 20260 31124
rect 19107 31093 19119 31096
rect 19061 31087 19119 31093
rect 20254 31084 20260 31096
rect 20312 31124 20318 31136
rect 20622 31124 20628 31136
rect 20312 31096 20628 31124
rect 20312 31084 20318 31096
rect 20622 31084 20628 31096
rect 20680 31084 20686 31136
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 16942 30880 16948 30932
rect 17000 30920 17006 30932
rect 20073 30923 20131 30929
rect 20073 30920 20085 30923
rect 17000 30892 20085 30920
rect 17000 30880 17006 30892
rect 20073 30889 20085 30892
rect 20119 30889 20131 30923
rect 20073 30883 20131 30889
rect 13814 30744 13820 30796
rect 13872 30784 13878 30796
rect 14093 30787 14151 30793
rect 14093 30784 14105 30787
rect 13872 30756 14105 30784
rect 13872 30744 13878 30756
rect 14093 30753 14105 30756
rect 14139 30753 14151 30787
rect 37826 30784 37832 30796
rect 37787 30756 37832 30784
rect 14093 30747 14151 30753
rect 9398 30716 9404 30728
rect 9359 30688 9404 30716
rect 9398 30676 9404 30688
rect 9456 30676 9462 30728
rect 14108 30716 14136 30747
rect 37826 30744 37832 30756
rect 37884 30744 37890 30796
rect 16666 30716 16672 30728
rect 14108 30688 16672 30716
rect 16666 30676 16672 30688
rect 16724 30676 16730 30728
rect 17126 30676 17132 30728
rect 17184 30716 17190 30728
rect 17770 30716 17776 30728
rect 17184 30688 17776 30716
rect 17184 30676 17190 30688
rect 17770 30676 17776 30688
rect 17828 30716 17834 30728
rect 20349 30719 20407 30725
rect 20349 30716 20361 30719
rect 17828 30688 20361 30716
rect 17828 30676 17834 30688
rect 20349 30685 20361 30688
rect 20395 30685 20407 30719
rect 20349 30679 20407 30685
rect 20438 30676 20444 30728
rect 20496 30725 20502 30728
rect 20496 30716 20504 30725
rect 38102 30716 38108 30728
rect 20496 30688 20541 30716
rect 38063 30688 38108 30716
rect 20496 30679 20504 30688
rect 20496 30676 20502 30679
rect 38102 30676 38108 30688
rect 38160 30676 38166 30728
rect 11422 30608 11428 30660
rect 11480 30648 11486 30660
rect 14338 30651 14396 30657
rect 14338 30648 14350 30651
rect 11480 30620 14350 30648
rect 11480 30608 11486 30620
rect 14338 30617 14350 30620
rect 14384 30617 14396 30651
rect 14338 30611 14396 30617
rect 17865 30651 17923 30657
rect 17865 30617 17877 30651
rect 17911 30648 17923 30651
rect 18046 30648 18052 30660
rect 17911 30620 18052 30648
rect 17911 30617 17923 30620
rect 17865 30611 17923 30617
rect 18046 30608 18052 30620
rect 18104 30648 18110 30660
rect 18506 30648 18512 30660
rect 18104 30620 18512 30648
rect 18104 30608 18110 30620
rect 18506 30608 18512 30620
rect 18564 30608 18570 30660
rect 20070 30648 20076 30660
rect 20031 30620 20076 30648
rect 20070 30608 20076 30620
rect 20128 30608 20134 30660
rect 20254 30648 20260 30660
rect 20215 30620 20260 30648
rect 20254 30608 20260 30620
rect 20312 30648 20318 30660
rect 21085 30651 21143 30657
rect 21085 30648 21097 30651
rect 20312 30620 21097 30648
rect 20312 30608 20318 30620
rect 21085 30617 21097 30620
rect 21131 30617 21143 30651
rect 21085 30611 21143 30617
rect 10686 30580 10692 30592
rect 10647 30552 10692 30580
rect 10686 30540 10692 30552
rect 10744 30540 10750 30592
rect 15378 30540 15384 30592
rect 15436 30580 15442 30592
rect 15473 30583 15531 30589
rect 15473 30580 15485 30583
rect 15436 30552 15485 30580
rect 15436 30540 15442 30552
rect 15473 30549 15485 30552
rect 15519 30549 15531 30583
rect 18322 30580 18328 30592
rect 18283 30552 18328 30580
rect 15473 30543 15531 30549
rect 18322 30540 18328 30552
rect 18380 30540 18386 30592
rect 1104 30490 38824 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 38824 30490
rect 1104 30416 38824 30438
rect 9309 30379 9367 30385
rect 9309 30345 9321 30379
rect 9355 30376 9367 30379
rect 9398 30376 9404 30388
rect 9355 30348 9404 30376
rect 9355 30345 9367 30348
rect 9309 30339 9367 30345
rect 9398 30336 9404 30348
rect 9456 30336 9462 30388
rect 14458 30336 14464 30388
rect 14516 30376 14522 30388
rect 14918 30376 14924 30388
rect 14516 30348 14924 30376
rect 14516 30336 14522 30348
rect 14918 30336 14924 30348
rect 14976 30376 14982 30388
rect 38102 30376 38108 30388
rect 14976 30348 19472 30376
rect 38063 30348 38108 30376
rect 14976 30336 14982 30348
rect 19444 30320 19472 30348
rect 38102 30336 38108 30348
rect 38160 30336 38166 30388
rect 16574 30268 16580 30320
rect 16632 30308 16638 30320
rect 16914 30311 16972 30317
rect 16914 30308 16926 30311
rect 16632 30280 16926 30308
rect 16632 30268 16638 30280
rect 16914 30277 16926 30280
rect 16960 30277 16972 30311
rect 19334 30308 19340 30320
rect 16914 30271 16972 30277
rect 18800 30280 19340 30308
rect 16666 30240 16672 30252
rect 16627 30212 16672 30240
rect 16666 30200 16672 30212
rect 16724 30200 16730 30252
rect 18800 30249 18828 30280
rect 19334 30268 19340 30280
rect 19392 30268 19398 30320
rect 19426 30268 19432 30320
rect 19484 30268 19490 30320
rect 19610 30268 19616 30320
rect 19668 30308 19674 30320
rect 19978 30308 19984 30320
rect 19668 30280 19984 30308
rect 19668 30268 19674 30280
rect 19978 30268 19984 30280
rect 20036 30308 20042 30320
rect 20438 30308 20444 30320
rect 20036 30280 20444 30308
rect 20036 30268 20042 30280
rect 20438 30268 20444 30280
rect 20496 30268 20502 30320
rect 18785 30243 18843 30249
rect 18785 30209 18797 30243
rect 18831 30209 18843 30243
rect 18785 30203 18843 30209
rect 19061 30243 19119 30249
rect 19061 30209 19073 30243
rect 19107 30240 19119 30243
rect 20070 30240 20076 30252
rect 19107 30212 20076 30240
rect 19107 30209 19119 30212
rect 19061 30203 19119 30209
rect 20070 30200 20076 30212
rect 20128 30200 20134 30252
rect 17954 30132 17960 30184
rect 18012 30172 18018 30184
rect 18509 30175 18567 30181
rect 18509 30172 18521 30175
rect 18012 30144 18521 30172
rect 18012 30132 18018 30144
rect 18509 30141 18521 30144
rect 18555 30172 18567 30175
rect 19337 30175 19395 30181
rect 18555 30144 18736 30172
rect 18555 30141 18567 30144
rect 18509 30135 18567 30141
rect 18601 30107 18659 30113
rect 18601 30104 18613 30107
rect 17604 30076 18613 30104
rect 6638 29996 6644 30048
rect 6696 30036 6702 30048
rect 17604 30036 17632 30076
rect 18601 30073 18613 30076
rect 18647 30073 18659 30107
rect 18708 30104 18736 30144
rect 19337 30141 19349 30175
rect 19383 30172 19395 30175
rect 20254 30172 20260 30184
rect 19383 30144 20260 30172
rect 19383 30141 19395 30144
rect 19337 30135 19395 30141
rect 19610 30104 19616 30116
rect 18708 30076 19616 30104
rect 18601 30067 18659 30073
rect 19610 30064 19616 30076
rect 19668 30064 19674 30116
rect 19812 30048 19840 30144
rect 20254 30132 20260 30144
rect 20312 30132 20318 30184
rect 6696 30008 17632 30036
rect 18049 30039 18107 30045
rect 6696 29996 6702 30008
rect 18049 30005 18061 30039
rect 18095 30036 18107 30039
rect 18966 30036 18972 30048
rect 18095 30008 18972 30036
rect 18095 30005 18107 30008
rect 18049 29999 18107 30005
rect 18966 29996 18972 30008
rect 19024 29996 19030 30048
rect 19794 30036 19800 30048
rect 19755 30008 19800 30036
rect 19794 29996 19800 30008
rect 19852 29996 19858 30048
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 12526 29792 12532 29844
rect 12584 29832 12590 29844
rect 13814 29832 13820 29844
rect 12584 29804 13820 29832
rect 12584 29792 12590 29804
rect 13814 29792 13820 29804
rect 13872 29832 13878 29844
rect 15746 29832 15752 29844
rect 13872 29804 15752 29832
rect 13872 29792 13878 29804
rect 15746 29792 15752 29804
rect 15804 29792 15810 29844
rect 16298 29792 16304 29844
rect 16356 29832 16362 29844
rect 16669 29835 16727 29841
rect 16669 29832 16681 29835
rect 16356 29804 16681 29832
rect 16356 29792 16362 29804
rect 16669 29801 16681 29804
rect 16715 29832 16727 29835
rect 17126 29832 17132 29844
rect 16715 29804 17132 29832
rect 16715 29801 16727 29804
rect 16669 29795 16727 29801
rect 17126 29792 17132 29804
rect 17184 29792 17190 29844
rect 11882 29724 11888 29776
rect 11940 29764 11946 29776
rect 18049 29767 18107 29773
rect 18049 29764 18061 29767
rect 11940 29736 18061 29764
rect 11940 29724 11946 29736
rect 18049 29733 18061 29736
rect 18095 29764 18107 29767
rect 18322 29764 18328 29776
rect 18095 29736 18328 29764
rect 18095 29733 18107 29736
rect 18049 29727 18107 29733
rect 18322 29724 18328 29736
rect 18380 29764 18386 29776
rect 18380 29736 19564 29764
rect 18380 29724 18386 29736
rect 18598 29696 18604 29708
rect 15212 29668 18604 29696
rect 12434 29588 12440 29640
rect 12492 29628 12498 29640
rect 15212 29628 15240 29668
rect 18598 29656 18604 29668
rect 18656 29656 18662 29708
rect 19426 29696 19432 29708
rect 19387 29668 19432 29696
rect 19426 29656 19432 29668
rect 19484 29656 19490 29708
rect 19536 29705 19564 29736
rect 19521 29699 19579 29705
rect 19521 29665 19533 29699
rect 19567 29665 19579 29699
rect 19521 29659 19579 29665
rect 12492 29600 15240 29628
rect 15289 29631 15347 29637
rect 12492 29588 12498 29600
rect 15289 29597 15301 29631
rect 15335 29597 15347 29631
rect 15289 29591 15347 29597
rect 15381 29631 15439 29637
rect 15381 29597 15393 29631
rect 15427 29628 15439 29631
rect 16942 29628 16948 29640
rect 15427 29600 16948 29628
rect 15427 29597 15439 29600
rect 15381 29591 15439 29597
rect 8846 29520 8852 29572
rect 8904 29560 8910 29572
rect 14734 29560 14740 29572
rect 8904 29532 14740 29560
rect 8904 29520 8910 29532
rect 14734 29520 14740 29532
rect 14792 29520 14798 29572
rect 15194 29560 15200 29572
rect 15155 29532 15200 29560
rect 15194 29520 15200 29532
rect 15252 29520 15258 29572
rect 11241 29495 11299 29501
rect 11241 29461 11253 29495
rect 11287 29492 11299 29495
rect 11882 29492 11888 29504
rect 11287 29464 11888 29492
rect 11287 29461 11299 29464
rect 11241 29455 11299 29461
rect 11882 29452 11888 29464
rect 11940 29452 11946 29504
rect 15102 29452 15108 29504
rect 15160 29492 15166 29504
rect 15304 29492 15332 29591
rect 16942 29588 16948 29600
rect 17000 29588 17006 29640
rect 19337 29631 19395 29637
rect 19337 29628 19349 29631
rect 18616 29600 19349 29628
rect 15657 29563 15715 29569
rect 15657 29529 15669 29563
rect 15703 29560 15715 29563
rect 15746 29560 15752 29572
rect 15703 29532 15752 29560
rect 15703 29529 15715 29532
rect 15657 29523 15715 29529
rect 15746 29520 15752 29532
rect 15804 29560 15810 29572
rect 16117 29563 16175 29569
rect 16117 29560 16129 29563
rect 15804 29532 16129 29560
rect 15804 29520 15810 29532
rect 16117 29529 16129 29532
rect 16163 29529 16175 29563
rect 16117 29523 16175 29529
rect 15562 29492 15568 29504
rect 15160 29464 15332 29492
rect 15523 29464 15568 29492
rect 15160 29452 15166 29464
rect 15562 29452 15568 29464
rect 15620 29452 15626 29504
rect 16022 29452 16028 29504
rect 16080 29492 16086 29504
rect 17218 29492 17224 29504
rect 16080 29464 17224 29492
rect 16080 29452 16086 29464
rect 17218 29452 17224 29464
rect 17276 29452 17282 29504
rect 18506 29452 18512 29504
rect 18564 29492 18570 29504
rect 18616 29501 18644 29600
rect 19337 29597 19349 29600
rect 19383 29597 19395 29631
rect 19337 29591 19395 29597
rect 19797 29631 19855 29637
rect 19797 29597 19809 29631
rect 19843 29628 19855 29631
rect 20070 29628 20076 29640
rect 19843 29600 20076 29628
rect 19843 29597 19855 29600
rect 19797 29591 19855 29597
rect 20070 29588 20076 29600
rect 20128 29628 20134 29640
rect 20254 29628 20260 29640
rect 20128 29600 20260 29628
rect 20128 29588 20134 29600
rect 20254 29588 20260 29600
rect 20312 29588 20318 29640
rect 19613 29563 19671 29569
rect 19613 29529 19625 29563
rect 19659 29529 19671 29563
rect 19613 29523 19671 29529
rect 18601 29495 18659 29501
rect 18601 29492 18613 29495
rect 18564 29464 18613 29492
rect 18564 29452 18570 29464
rect 18601 29461 18613 29464
rect 18647 29461 18659 29495
rect 18601 29455 18659 29461
rect 19058 29452 19064 29504
rect 19116 29492 19122 29504
rect 19245 29495 19303 29501
rect 19245 29492 19257 29495
rect 19116 29464 19257 29492
rect 19116 29452 19122 29464
rect 19245 29461 19257 29464
rect 19291 29461 19303 29495
rect 19628 29492 19656 29523
rect 19794 29492 19800 29504
rect 19628 29464 19800 29492
rect 19245 29455 19303 29461
rect 19794 29452 19800 29464
rect 19852 29492 19858 29504
rect 20349 29495 20407 29501
rect 20349 29492 20361 29495
rect 19852 29464 20361 29492
rect 19852 29452 19858 29464
rect 20349 29461 20361 29464
rect 20395 29492 20407 29495
rect 20438 29492 20444 29504
rect 20395 29464 20444 29492
rect 20395 29461 20407 29464
rect 20349 29455 20407 29461
rect 20438 29452 20444 29464
rect 20496 29452 20502 29504
rect 1104 29402 38824 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 38824 29402
rect 1104 29328 38824 29350
rect 8846 29288 8852 29300
rect 8807 29260 8852 29288
rect 8846 29248 8852 29260
rect 8904 29248 8910 29300
rect 15194 29288 15200 29300
rect 10060 29260 15200 29288
rect 7736 29223 7794 29229
rect 7736 29189 7748 29223
rect 7782 29220 7794 29223
rect 10060 29220 10088 29260
rect 15194 29248 15200 29260
rect 15252 29248 15258 29300
rect 16942 29248 16948 29300
rect 17000 29288 17006 29300
rect 17218 29288 17224 29300
rect 17000 29260 17045 29288
rect 17144 29260 17224 29288
rect 17000 29248 17006 29260
rect 7782 29192 10088 29220
rect 11885 29223 11943 29229
rect 7782 29189 7794 29192
rect 7736 29183 7794 29189
rect 11885 29189 11897 29223
rect 11931 29220 11943 29223
rect 12526 29220 12532 29232
rect 11931 29192 12532 29220
rect 11931 29189 11943 29192
rect 11885 29183 11943 29189
rect 12526 29180 12532 29192
rect 12584 29180 12590 29232
rect 12618 29180 12624 29232
rect 12676 29220 12682 29232
rect 16022 29220 16028 29232
rect 12676 29192 14412 29220
rect 12676 29180 12682 29192
rect 10962 29152 10968 29164
rect 10875 29124 10968 29152
rect 10962 29112 10968 29124
rect 11020 29152 11026 29164
rect 11698 29152 11704 29164
rect 11020 29124 11704 29152
rect 11020 29112 11026 29124
rect 11698 29112 11704 29124
rect 11756 29112 11762 29164
rect 11977 29155 12035 29161
rect 11977 29152 11989 29155
rect 11900 29124 11989 29152
rect 11900 29096 11928 29124
rect 11977 29121 11989 29124
rect 12023 29121 12035 29155
rect 11977 29115 12035 29121
rect 12802 29112 12808 29164
rect 12860 29152 12866 29164
rect 13245 29155 13303 29161
rect 13245 29152 13257 29155
rect 12860 29124 13257 29152
rect 12860 29112 12866 29124
rect 13245 29121 13257 29124
rect 13291 29121 13303 29155
rect 13245 29115 13303 29121
rect 7466 29084 7472 29096
rect 7427 29056 7472 29084
rect 7466 29044 7472 29056
rect 7524 29044 7530 29096
rect 11882 29044 11888 29096
rect 11940 29044 11946 29096
rect 12250 29044 12256 29096
rect 12308 29084 12314 29096
rect 12989 29087 13047 29093
rect 12989 29084 13001 29087
rect 12308 29056 13001 29084
rect 12308 29044 12314 29056
rect 12989 29053 13001 29056
rect 13035 29053 13047 29087
rect 12989 29047 13047 29053
rect 11514 29016 11520 29028
rect 11475 28988 11520 29016
rect 11514 28976 11520 28988
rect 11572 28976 11578 29028
rect 14384 29025 14412 29192
rect 15212 29192 16028 29220
rect 15212 29164 15240 29192
rect 16022 29180 16028 29192
rect 16080 29180 16086 29232
rect 17144 29229 17172 29260
rect 17218 29248 17224 29260
rect 17276 29248 17282 29300
rect 17402 29248 17408 29300
rect 17460 29288 17466 29300
rect 20070 29288 20076 29300
rect 17460 29260 20076 29288
rect 17460 29248 17466 29260
rect 20070 29248 20076 29260
rect 20128 29248 20134 29300
rect 17129 29223 17187 29229
rect 16849 29189 16907 29195
rect 16849 29186 16861 29189
rect 15194 29112 15200 29164
rect 15252 29112 15258 29164
rect 16684 29158 16861 29186
rect 16684 29152 16712 29158
rect 15488 29124 16712 29152
rect 16849 29155 16861 29158
rect 16895 29155 16907 29189
rect 17129 29189 17141 29223
rect 17175 29189 17187 29223
rect 17129 29183 17187 29189
rect 19242 29180 19248 29232
rect 19300 29220 19306 29232
rect 19797 29223 19855 29229
rect 19797 29220 19809 29223
rect 19300 29192 19809 29220
rect 19300 29180 19306 29192
rect 19797 29189 19809 29192
rect 19843 29189 19855 29223
rect 19797 29183 19855 29189
rect 16849 29149 16907 29155
rect 14734 29044 14740 29096
rect 14792 29084 14798 29096
rect 15488 29093 15516 29124
rect 17218 29112 17224 29164
rect 17276 29152 17282 29164
rect 17276 29124 17321 29152
rect 17276 29112 17282 29124
rect 18414 29112 18420 29164
rect 18472 29152 18478 29164
rect 18874 29152 18880 29164
rect 18472 29124 18880 29152
rect 18472 29112 18478 29124
rect 18874 29112 18880 29124
rect 18932 29112 18938 29164
rect 19337 29155 19395 29161
rect 19337 29121 19349 29155
rect 19383 29152 19395 29155
rect 21174 29152 21180 29164
rect 19383 29124 21180 29152
rect 19383 29121 19395 29124
rect 19337 29115 19395 29121
rect 21174 29112 21180 29124
rect 21232 29112 21238 29164
rect 15473 29087 15531 29093
rect 15473 29084 15485 29087
rect 14792 29056 15485 29084
rect 14792 29044 14798 29056
rect 15473 29053 15485 29056
rect 15519 29053 15531 29087
rect 17037 29087 17095 29093
rect 15473 29047 15531 29053
rect 16776 29048 16957 29076
rect 14369 29019 14427 29025
rect 14369 28985 14381 29019
rect 14415 29016 14427 29019
rect 16776 29016 16804 29048
rect 14415 28988 16804 29016
rect 16929 29016 16957 29048
rect 17037 29053 17049 29087
rect 17083 29084 17095 29087
rect 17126 29084 17132 29096
rect 17083 29056 17132 29084
rect 17083 29053 17095 29056
rect 17037 29047 17095 29053
rect 17126 29044 17132 29056
rect 17184 29084 17190 29096
rect 17402 29084 17408 29096
rect 17184 29056 17408 29084
rect 17184 29044 17190 29056
rect 17402 29044 17408 29056
rect 17460 29044 17466 29096
rect 19058 29084 19064 29096
rect 19019 29056 19064 29084
rect 19058 29044 19064 29056
rect 19116 29044 19122 29096
rect 18874 29016 18880 29028
rect 16929 28988 18880 29016
rect 14415 28985 14427 28988
rect 14369 28979 14427 28985
rect 18874 28976 18880 28988
rect 18932 28976 18938 29028
rect 19150 29016 19156 29028
rect 19111 28988 19156 29016
rect 19150 28976 19156 28988
rect 19208 28976 19214 29028
rect 19245 29019 19303 29025
rect 19245 28985 19257 29019
rect 19291 29016 19303 29019
rect 19426 29016 19432 29028
rect 19291 28988 19432 29016
rect 19291 28985 19303 28988
rect 19245 28979 19303 28985
rect 19426 28976 19432 28988
rect 19484 28976 19490 29028
rect 13354 28908 13360 28960
rect 13412 28948 13418 28960
rect 20530 28948 20536 28960
rect 13412 28920 20536 28948
rect 13412 28908 13418 28920
rect 20530 28908 20536 28920
rect 20588 28908 20594 28960
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 12802 28744 12808 28756
rect 12763 28716 12808 28744
rect 12802 28704 12808 28716
rect 12860 28704 12866 28756
rect 15841 28747 15899 28753
rect 15841 28713 15853 28747
rect 15887 28744 15899 28747
rect 16482 28744 16488 28756
rect 15887 28716 16488 28744
rect 15887 28713 15899 28716
rect 15841 28707 15899 28713
rect 16482 28704 16488 28716
rect 16540 28704 16546 28756
rect 18598 28744 18604 28756
rect 18559 28716 18604 28744
rect 18598 28704 18604 28716
rect 18656 28704 18662 28756
rect 19245 28747 19303 28753
rect 19245 28713 19257 28747
rect 19291 28744 19303 28747
rect 19334 28744 19340 28756
rect 19291 28716 19340 28744
rect 19291 28713 19303 28716
rect 19245 28707 19303 28713
rect 19334 28704 19340 28716
rect 19392 28704 19398 28756
rect 11882 28636 11888 28688
rect 11940 28676 11946 28688
rect 12434 28676 12440 28688
rect 11940 28648 12440 28676
rect 11940 28636 11946 28648
rect 12434 28636 12440 28648
rect 12492 28636 12498 28688
rect 7009 28543 7067 28549
rect 7009 28509 7021 28543
rect 7055 28540 7067 28543
rect 10413 28543 10471 28549
rect 10413 28540 10425 28543
rect 7055 28512 10425 28540
rect 7055 28509 7067 28512
rect 7009 28503 7067 28509
rect 10413 28509 10425 28512
rect 10459 28540 10471 28543
rect 10686 28540 10692 28552
rect 10459 28512 10692 28540
rect 10459 28509 10471 28512
rect 10413 28503 10471 28509
rect 10686 28500 10692 28512
rect 10744 28500 10750 28552
rect 11790 28500 11796 28552
rect 11848 28540 11854 28552
rect 12621 28543 12679 28549
rect 12621 28540 12633 28543
rect 11848 28512 12633 28540
rect 11848 28500 11854 28512
rect 12621 28509 12633 28512
rect 12667 28509 12679 28543
rect 12621 28503 12679 28509
rect 16666 28500 16672 28552
rect 16724 28540 16730 28552
rect 17221 28543 17279 28549
rect 17221 28540 17233 28543
rect 16724 28512 17233 28540
rect 16724 28500 16730 28512
rect 17221 28509 17233 28512
rect 17267 28509 17279 28543
rect 17221 28503 17279 28509
rect 19426 28500 19432 28552
rect 19484 28540 19490 28552
rect 19521 28543 19579 28549
rect 19521 28540 19533 28543
rect 19484 28512 19533 28540
rect 19484 28500 19490 28512
rect 19521 28509 19533 28512
rect 19567 28509 19579 28543
rect 19521 28503 19579 28509
rect 12161 28475 12219 28481
rect 12161 28441 12173 28475
rect 12207 28472 12219 28475
rect 12250 28472 12256 28484
rect 12207 28444 12256 28472
rect 12207 28441 12219 28444
rect 12161 28435 12219 28441
rect 12250 28432 12256 28444
rect 12308 28432 12314 28484
rect 16850 28432 16856 28484
rect 16908 28472 16914 28484
rect 16954 28475 17012 28481
rect 16954 28472 16966 28475
rect 16908 28444 16966 28472
rect 16908 28432 16914 28444
rect 16954 28441 16966 28444
rect 17000 28441 17012 28475
rect 16954 28435 17012 28441
rect 18782 28432 18788 28484
rect 18840 28472 18846 28484
rect 19242 28472 19248 28484
rect 18840 28444 19248 28472
rect 18840 28432 18846 28444
rect 19242 28432 19248 28444
rect 19300 28432 19306 28484
rect 2498 28364 2504 28416
rect 2556 28404 2562 28416
rect 5537 28407 5595 28413
rect 5537 28404 5549 28407
rect 2556 28376 5549 28404
rect 2556 28364 2562 28376
rect 5537 28373 5549 28376
rect 5583 28404 5595 28407
rect 7466 28404 7472 28416
rect 5583 28376 7472 28404
rect 5583 28373 5595 28376
rect 5537 28367 5595 28373
rect 7466 28364 7472 28376
rect 7524 28364 7530 28416
rect 9858 28404 9864 28416
rect 9819 28376 9864 28404
rect 9858 28364 9864 28376
rect 9916 28364 9922 28416
rect 9950 28364 9956 28416
rect 10008 28404 10014 28416
rect 18506 28404 18512 28416
rect 10008 28376 18512 28404
rect 10008 28364 10014 28376
rect 18506 28364 18512 28376
rect 18564 28364 18570 28416
rect 18690 28364 18696 28416
rect 18748 28404 18754 28416
rect 19429 28407 19487 28413
rect 19429 28404 19441 28407
rect 18748 28376 19441 28404
rect 18748 28364 18754 28376
rect 19429 28373 19441 28376
rect 19475 28373 19487 28407
rect 19429 28367 19487 28373
rect 20257 28407 20315 28413
rect 20257 28373 20269 28407
rect 20303 28404 20315 28407
rect 20438 28404 20444 28416
rect 20303 28376 20444 28404
rect 20303 28373 20315 28376
rect 20257 28367 20315 28373
rect 20438 28364 20444 28376
rect 20496 28364 20502 28416
rect 1104 28314 38824 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 38824 28314
rect 1104 28240 38824 28262
rect 3881 28203 3939 28209
rect 3881 28169 3893 28203
rect 3927 28200 3939 28203
rect 13354 28200 13360 28212
rect 3927 28172 13360 28200
rect 3927 28169 3939 28172
rect 3881 28163 3939 28169
rect 13354 28160 13360 28172
rect 13412 28160 13418 28212
rect 13630 28200 13636 28212
rect 13591 28172 13636 28200
rect 13630 28160 13636 28172
rect 13688 28160 13694 28212
rect 17862 28200 17868 28212
rect 14476 28172 17868 28200
rect 10042 28092 10048 28144
rect 10100 28132 10106 28144
rect 12498 28135 12556 28141
rect 12498 28132 12510 28135
rect 10100 28104 12510 28132
rect 10100 28092 10106 28104
rect 12498 28101 12510 28104
rect 12544 28101 12556 28135
rect 12498 28095 12556 28101
rect 12618 28092 12624 28144
rect 12676 28092 12682 28144
rect 1394 28024 1400 28076
rect 1452 28064 1458 28076
rect 2498 28064 2504 28076
rect 1452 28036 2504 28064
rect 1452 28024 1458 28036
rect 2498 28024 2504 28036
rect 2556 28024 2562 28076
rect 2768 28067 2826 28073
rect 2768 28033 2780 28067
rect 2814 28064 2826 28067
rect 4062 28064 4068 28076
rect 2814 28036 4068 28064
rect 2814 28033 2826 28036
rect 2768 28027 2826 28033
rect 4062 28024 4068 28036
rect 4120 28024 4126 28076
rect 9309 28067 9367 28073
rect 9309 28033 9321 28067
rect 9355 28064 9367 28067
rect 9769 28067 9827 28073
rect 9769 28064 9781 28067
rect 9355 28036 9781 28064
rect 9355 28033 9367 28036
rect 9309 28027 9367 28033
rect 9769 28033 9781 28036
rect 9815 28064 9827 28067
rect 9950 28064 9956 28076
rect 9815 28036 9956 28064
rect 9815 28033 9827 28036
rect 9769 28027 9827 28033
rect 9950 28024 9956 28036
rect 10008 28024 10014 28076
rect 10686 28064 10692 28076
rect 10647 28036 10692 28064
rect 10686 28024 10692 28036
rect 10744 28064 10750 28076
rect 11793 28067 11851 28073
rect 11793 28064 11805 28067
rect 10744 28036 11805 28064
rect 10744 28024 10750 28036
rect 11793 28033 11805 28036
rect 11839 28064 11851 28067
rect 11882 28064 11888 28076
rect 11839 28036 11888 28064
rect 11839 28033 11851 28036
rect 11793 28027 11851 28033
rect 11882 28024 11888 28036
rect 11940 28024 11946 28076
rect 12342 28024 12348 28076
rect 12400 28064 12406 28076
rect 12636 28064 12664 28092
rect 14274 28064 14280 28076
rect 12400 28036 12664 28064
rect 14235 28036 14280 28064
rect 12400 28024 12406 28036
rect 14274 28024 14280 28036
rect 14332 28024 14338 28076
rect 14476 28064 14504 28172
rect 17862 28160 17868 28172
rect 17920 28160 17926 28212
rect 18046 28160 18052 28212
rect 18104 28200 18110 28212
rect 18141 28203 18199 28209
rect 18141 28200 18153 28203
rect 18104 28172 18153 28200
rect 18104 28160 18110 28172
rect 18141 28169 18153 28172
rect 18187 28169 18199 28203
rect 18141 28163 18199 28169
rect 18230 28160 18236 28212
rect 18288 28200 18294 28212
rect 18288 28172 18381 28200
rect 18288 28160 18294 28172
rect 14553 28135 14611 28141
rect 14553 28101 14565 28135
rect 14599 28132 14611 28135
rect 18340 28132 18368 28172
rect 18506 28160 18512 28212
rect 18564 28200 18570 28212
rect 21085 28203 21143 28209
rect 21085 28200 21097 28203
rect 18564 28172 21097 28200
rect 18564 28160 18570 28172
rect 14599 28104 18368 28132
rect 14599 28101 14611 28104
rect 14553 28095 14611 28101
rect 18598 28092 18604 28144
rect 18656 28132 18662 28144
rect 18656 28104 19932 28132
rect 18656 28092 18662 28104
rect 14645 28067 14703 28073
rect 14645 28064 14657 28067
rect 14476 28036 14657 28064
rect 14645 28033 14657 28036
rect 14691 28033 14703 28067
rect 14645 28027 14703 28033
rect 15289 28067 15347 28073
rect 15289 28033 15301 28067
rect 15335 28064 15347 28067
rect 17954 28064 17960 28076
rect 15335 28036 17960 28064
rect 15335 28033 15347 28036
rect 15289 28027 15347 28033
rect 17954 28024 17960 28036
rect 18012 28024 18018 28076
rect 18049 28067 18107 28073
rect 18049 28033 18061 28067
rect 18095 28064 18107 28067
rect 18138 28064 18144 28076
rect 18095 28036 18144 28064
rect 18095 28033 18107 28036
rect 18049 28027 18107 28033
rect 18138 28024 18144 28036
rect 18196 28024 18202 28076
rect 18874 28064 18880 28076
rect 18835 28036 18880 28064
rect 18874 28024 18880 28036
rect 18932 28024 18938 28076
rect 19904 28073 19932 28104
rect 19996 28073 20024 28172
rect 21085 28169 21097 28172
rect 21131 28169 21143 28203
rect 21085 28163 21143 28169
rect 20530 28132 20536 28144
rect 20491 28104 20536 28132
rect 20530 28092 20536 28104
rect 20588 28092 20594 28144
rect 19889 28067 19947 28073
rect 19889 28033 19901 28067
rect 19935 28033 19947 28067
rect 19889 28027 19947 28033
rect 19981 28067 20039 28073
rect 19981 28033 19993 28067
rect 20027 28033 20039 28067
rect 19981 28027 20039 28033
rect 9861 27999 9919 28005
rect 9861 27965 9873 27999
rect 9907 27996 9919 27999
rect 10318 27996 10324 28008
rect 9907 27968 10324 27996
rect 9907 27965 9919 27968
rect 9861 27959 9919 27965
rect 10318 27956 10324 27968
rect 10376 27996 10382 28008
rect 10597 27999 10655 28005
rect 10597 27996 10609 27999
rect 10376 27968 10609 27996
rect 10376 27956 10382 27968
rect 10597 27965 10609 27968
rect 10643 27965 10655 27999
rect 10597 27959 10655 27965
rect 10781 27999 10839 28005
rect 10781 27965 10793 27999
rect 10827 27965 10839 27999
rect 10781 27959 10839 27965
rect 8386 27888 8392 27940
rect 8444 27928 8450 27940
rect 10413 27931 10471 27937
rect 10413 27928 10425 27931
rect 8444 27900 10425 27928
rect 8444 27888 8450 27900
rect 10413 27897 10425 27900
rect 10459 27897 10471 27931
rect 10413 27891 10471 27897
rect 10134 27820 10140 27872
rect 10192 27860 10198 27872
rect 10796 27860 10824 27959
rect 10870 27956 10876 28008
rect 10928 27996 10934 28008
rect 12250 27996 12256 28008
rect 10928 27968 10973 27996
rect 12211 27968 12256 27996
rect 10928 27956 10934 27968
rect 12250 27956 12256 27968
rect 12308 27956 12314 28008
rect 14461 27999 14519 28005
rect 14461 27965 14473 27999
rect 14507 27996 14519 27999
rect 17770 27996 17776 28008
rect 14507 27968 17776 27996
rect 14507 27965 14519 27968
rect 14461 27959 14519 27965
rect 17770 27956 17776 27968
rect 17828 27996 17834 28008
rect 18417 27999 18475 28005
rect 18417 27996 18429 27999
rect 17828 27968 18429 27996
rect 17828 27956 17834 27968
rect 18417 27965 18429 27968
rect 18463 27965 18475 27999
rect 18417 27959 18475 27965
rect 18969 27999 19027 28005
rect 18969 27965 18981 27999
rect 19015 27996 19027 27999
rect 19521 27999 19579 28005
rect 19521 27996 19533 27999
rect 19015 27968 19533 27996
rect 19015 27965 19027 27968
rect 18969 27959 19027 27965
rect 19521 27965 19533 27968
rect 19567 27965 19579 27999
rect 19521 27959 19579 27965
rect 19705 27999 19763 28005
rect 19705 27965 19717 27999
rect 19751 27965 19763 27999
rect 19705 27959 19763 27965
rect 19797 27999 19855 28005
rect 19797 27965 19809 27999
rect 19843 27996 19855 27999
rect 20438 27996 20444 28008
rect 19843 27968 20444 27996
rect 19843 27965 19855 27968
rect 19797 27959 19855 27965
rect 14277 27931 14335 27937
rect 14277 27897 14289 27931
rect 14323 27928 14335 27931
rect 16758 27928 16764 27940
rect 14323 27900 16764 27928
rect 14323 27897 14335 27900
rect 14277 27891 14335 27897
rect 16758 27888 16764 27900
rect 16816 27888 16822 27940
rect 17494 27928 17500 27940
rect 17455 27900 17500 27928
rect 17494 27888 17500 27900
rect 17552 27888 17558 27940
rect 18432 27928 18460 27959
rect 19058 27928 19064 27940
rect 18432 27900 19064 27928
rect 19058 27888 19064 27900
rect 19116 27888 19122 27940
rect 19720 27928 19748 27959
rect 20438 27956 20444 27968
rect 20496 27956 20502 28008
rect 20254 27928 20260 27940
rect 19720 27900 20260 27928
rect 20254 27888 20260 27900
rect 20312 27888 20318 27940
rect 10192 27832 10824 27860
rect 11701 27863 11759 27869
rect 10192 27820 10198 27832
rect 11701 27829 11713 27863
rect 11747 27860 11759 27863
rect 11974 27860 11980 27872
rect 11747 27832 11980 27860
rect 11747 27829 11759 27832
rect 11701 27823 11759 27829
rect 11974 27820 11980 27832
rect 12032 27820 12038 27872
rect 15470 27860 15476 27872
rect 15431 27832 15476 27860
rect 15470 27820 15476 27832
rect 15528 27820 15534 27872
rect 18325 27863 18383 27869
rect 18325 27829 18337 27863
rect 18371 27860 18383 27863
rect 18414 27860 18420 27872
rect 18371 27832 18420 27860
rect 18371 27829 18383 27832
rect 18325 27823 18383 27829
rect 18414 27820 18420 27832
rect 18472 27820 18478 27872
rect 19886 27820 19892 27872
rect 19944 27860 19950 27872
rect 20073 27863 20131 27869
rect 20073 27860 20085 27863
rect 19944 27832 20085 27860
rect 19944 27820 19950 27832
rect 20073 27829 20085 27832
rect 20119 27829 20131 27863
rect 20073 27823 20131 27829
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 2777 27659 2835 27665
rect 2777 27625 2789 27659
rect 2823 27625 2835 27659
rect 18046 27656 18052 27668
rect 2777 27619 2835 27625
rect 17880 27628 18052 27656
rect 2792 27588 2820 27619
rect 9858 27588 9864 27600
rect 2792 27560 9864 27588
rect 9858 27548 9864 27560
rect 9916 27588 9922 27600
rect 10505 27591 10563 27597
rect 10505 27588 10517 27591
rect 9916 27560 10517 27588
rect 9916 27548 9922 27560
rect 10505 27557 10517 27560
rect 10551 27588 10563 27591
rect 10686 27588 10692 27600
rect 10551 27560 10692 27588
rect 10551 27557 10563 27560
rect 10505 27551 10563 27557
rect 10686 27548 10692 27560
rect 10744 27548 10750 27600
rect 11790 27588 11796 27600
rect 11751 27560 11796 27588
rect 11790 27548 11796 27560
rect 11848 27548 11854 27600
rect 17313 27591 17371 27597
rect 17313 27557 17325 27591
rect 17359 27588 17371 27591
rect 17880 27588 17908 27628
rect 18046 27616 18052 27628
rect 18104 27616 18110 27668
rect 18509 27659 18567 27665
rect 18509 27625 18521 27659
rect 18555 27656 18567 27659
rect 19426 27656 19432 27668
rect 18555 27628 19432 27656
rect 18555 27625 18567 27628
rect 18509 27619 18567 27625
rect 19426 27616 19432 27628
rect 19484 27616 19490 27668
rect 17359 27560 17908 27588
rect 17359 27557 17371 27560
rect 17313 27551 17371 27557
rect 17954 27548 17960 27600
rect 18012 27588 18018 27600
rect 18325 27591 18383 27597
rect 18325 27588 18337 27591
rect 18012 27560 18337 27588
rect 18012 27548 18018 27560
rect 18325 27557 18337 27560
rect 18371 27557 18383 27591
rect 18325 27551 18383 27557
rect 20530 27548 20536 27600
rect 20588 27588 20594 27600
rect 20901 27591 20959 27597
rect 20901 27588 20913 27591
rect 20588 27560 20913 27588
rect 20588 27548 20594 27560
rect 20901 27557 20913 27560
rect 20947 27557 20959 27591
rect 21634 27588 21640 27600
rect 21595 27560 21640 27588
rect 20901 27551 20959 27557
rect 21634 27548 21640 27560
rect 21692 27548 21698 27600
rect 1394 27520 1400 27532
rect 1355 27492 1400 27520
rect 1394 27480 1400 27492
rect 1452 27480 1458 27532
rect 2774 27480 2780 27532
rect 2832 27520 2838 27532
rect 9585 27523 9643 27529
rect 2832 27492 9352 27520
rect 2832 27480 2838 27492
rect 9324 27461 9352 27492
rect 9585 27489 9597 27523
rect 9631 27520 9643 27523
rect 10870 27520 10876 27532
rect 9631 27492 10876 27520
rect 9631 27489 9643 27492
rect 9585 27483 9643 27489
rect 10870 27480 10876 27492
rect 10928 27520 10934 27532
rect 11241 27523 11299 27529
rect 11241 27520 11253 27523
rect 10928 27492 11253 27520
rect 10928 27480 10934 27492
rect 11241 27489 11253 27492
rect 11287 27520 11299 27523
rect 14182 27520 14188 27532
rect 11287 27492 14188 27520
rect 11287 27489 11299 27492
rect 11241 27483 11299 27489
rect 14182 27480 14188 27492
rect 14240 27480 14246 27532
rect 19334 27520 19340 27532
rect 17052 27492 19340 27520
rect 7653 27455 7711 27461
rect 7653 27421 7665 27455
rect 7699 27452 7711 27455
rect 9309 27455 9367 27461
rect 7699 27424 8984 27452
rect 7699 27421 7711 27424
rect 7653 27415 7711 27421
rect 1664 27387 1722 27393
rect 1664 27353 1676 27387
rect 1710 27384 1722 27387
rect 8386 27384 8392 27396
rect 1710 27356 8392 27384
rect 1710 27353 1722 27356
rect 1664 27347 1722 27353
rect 8386 27344 8392 27356
rect 8444 27344 8450 27396
rect 3878 27276 3884 27328
rect 3936 27316 3942 27328
rect 8956 27325 8984 27424
rect 9309 27421 9321 27455
rect 9355 27452 9367 27455
rect 9950 27452 9956 27464
rect 9355 27424 9956 27452
rect 9355 27421 9367 27424
rect 9309 27415 9367 27421
rect 9950 27412 9956 27424
rect 10008 27412 10014 27464
rect 11425 27455 11483 27461
rect 11425 27421 11437 27455
rect 11471 27452 11483 27455
rect 12342 27452 12348 27464
rect 11471 27424 12348 27452
rect 11471 27421 11483 27424
rect 11425 27415 11483 27421
rect 12342 27412 12348 27424
rect 12400 27412 12406 27464
rect 12986 27452 12992 27464
rect 12947 27424 12992 27452
rect 12986 27412 12992 27424
rect 13044 27412 13050 27464
rect 15933 27455 15991 27461
rect 15933 27421 15945 27455
rect 15979 27452 15991 27455
rect 16666 27452 16672 27464
rect 15979 27424 16672 27452
rect 15979 27421 15991 27424
rect 15933 27415 15991 27421
rect 16666 27412 16672 27424
rect 16724 27412 16730 27464
rect 9858 27344 9864 27396
rect 9916 27384 9922 27396
rect 11974 27384 11980 27396
rect 9916 27356 11980 27384
rect 9916 27344 9922 27356
rect 11974 27344 11980 27356
rect 12032 27344 12038 27396
rect 12897 27387 12955 27393
rect 12897 27353 12909 27387
rect 12943 27384 12955 27387
rect 14458 27384 14464 27396
rect 12943 27356 14464 27384
rect 12943 27353 12955 27356
rect 12897 27347 12955 27353
rect 14458 27344 14464 27356
rect 14516 27344 14522 27396
rect 15470 27344 15476 27396
rect 15528 27384 15534 27396
rect 16178 27387 16236 27393
rect 16178 27384 16190 27387
rect 15528 27356 16190 27384
rect 15528 27344 15534 27356
rect 16178 27353 16190 27356
rect 16224 27353 16236 27387
rect 16178 27347 16236 27353
rect 7469 27319 7527 27325
rect 7469 27316 7481 27319
rect 3936 27288 7481 27316
rect 3936 27276 3942 27288
rect 7469 27285 7481 27288
rect 7515 27285 7527 27319
rect 7469 27279 7527 27285
rect 8941 27319 8999 27325
rect 8941 27285 8953 27319
rect 8987 27285 8999 27319
rect 8941 27279 8999 27285
rect 9398 27276 9404 27328
rect 9456 27316 9462 27328
rect 11330 27316 11336 27328
rect 9456 27288 9501 27316
rect 11291 27288 11336 27316
rect 9456 27276 9462 27288
rect 11330 27276 11336 27288
rect 11388 27316 11394 27328
rect 12253 27319 12311 27325
rect 12253 27316 12265 27319
rect 11388 27288 12265 27316
rect 11388 27276 11394 27288
rect 12253 27285 12265 27288
rect 12299 27285 12311 27319
rect 12253 27279 12311 27285
rect 14185 27319 14243 27325
rect 14185 27285 14197 27319
rect 14231 27316 14243 27319
rect 14734 27316 14740 27328
rect 14231 27288 14740 27316
rect 14231 27285 14243 27288
rect 14185 27279 14243 27285
rect 14734 27276 14740 27288
rect 14792 27276 14798 27328
rect 15194 27316 15200 27328
rect 15155 27288 15200 27316
rect 15194 27276 15200 27288
rect 15252 27276 15258 27328
rect 16022 27276 16028 27328
rect 16080 27316 16086 27328
rect 17052 27316 17080 27492
rect 19334 27480 19340 27492
rect 19392 27520 19398 27532
rect 20073 27523 20131 27529
rect 20073 27520 20085 27523
rect 19392 27492 20085 27520
rect 19392 27480 19398 27492
rect 20073 27489 20085 27492
rect 20119 27489 20131 27523
rect 20073 27483 20131 27489
rect 17126 27412 17132 27464
rect 17184 27452 17190 27464
rect 19886 27452 19892 27464
rect 17184 27424 18736 27452
rect 19847 27424 19892 27452
rect 17184 27412 17190 27424
rect 18414 27344 18420 27396
rect 18472 27393 18478 27396
rect 18708 27393 18736 27424
rect 19886 27412 19892 27424
rect 19944 27412 19950 27464
rect 20165 27455 20223 27461
rect 20165 27421 20177 27455
rect 20211 27452 20223 27455
rect 22094 27452 22100 27464
rect 20211 27424 22100 27452
rect 20211 27421 20223 27424
rect 20165 27415 20223 27421
rect 22094 27412 22100 27424
rect 22152 27412 22158 27464
rect 18472 27387 18535 27393
rect 18472 27353 18489 27387
rect 18523 27353 18535 27387
rect 18472 27347 18535 27353
rect 18693 27387 18751 27393
rect 18693 27353 18705 27387
rect 18739 27353 18751 27387
rect 19702 27384 19708 27396
rect 19663 27356 19708 27384
rect 18693 27347 18751 27353
rect 18472 27344 18478 27347
rect 19702 27344 19708 27356
rect 19760 27344 19766 27396
rect 20622 27384 20628 27396
rect 20583 27356 20628 27384
rect 20622 27344 20628 27356
rect 20680 27344 20686 27396
rect 16080 27288 17080 27316
rect 17865 27319 17923 27325
rect 16080 27276 16086 27288
rect 17865 27285 17877 27319
rect 17911 27316 17923 27319
rect 18874 27316 18880 27328
rect 17911 27288 18880 27316
rect 17911 27285 17923 27288
rect 17865 27279 17923 27285
rect 18874 27276 18880 27288
rect 18932 27276 18938 27328
rect 19242 27276 19248 27328
rect 19300 27316 19306 27328
rect 19518 27316 19524 27328
rect 19300 27288 19524 27316
rect 19300 27276 19306 27288
rect 19518 27276 19524 27288
rect 19576 27276 19582 27328
rect 21082 27316 21088 27328
rect 21043 27288 21088 27316
rect 21082 27276 21088 27288
rect 21140 27276 21146 27328
rect 1104 27226 38824 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 38824 27226
rect 1104 27152 38824 27174
rect 9674 27112 9680 27124
rect 9635 27084 9680 27112
rect 9674 27072 9680 27084
rect 9732 27072 9738 27124
rect 12345 27115 12403 27121
rect 12345 27112 12357 27115
rect 9968 27084 12357 27112
rect 7920 27047 7978 27053
rect 7920 27013 7932 27047
rect 7966 27044 7978 27047
rect 9968 27044 9996 27084
rect 12345 27081 12357 27084
rect 12391 27081 12403 27115
rect 12345 27075 12403 27081
rect 14093 27115 14151 27121
rect 14093 27081 14105 27115
rect 14139 27112 14151 27115
rect 14274 27112 14280 27124
rect 14139 27084 14280 27112
rect 14139 27081 14151 27084
rect 14093 27075 14151 27081
rect 14274 27072 14280 27084
rect 14332 27072 14338 27124
rect 15749 27115 15807 27121
rect 15749 27081 15761 27115
rect 15795 27112 15807 27115
rect 15930 27112 15936 27124
rect 15795 27084 15936 27112
rect 15795 27081 15807 27084
rect 15749 27075 15807 27081
rect 15930 27072 15936 27084
rect 15988 27072 15994 27124
rect 16114 27072 16120 27124
rect 16172 27112 16178 27124
rect 16172 27084 18644 27112
rect 16172 27072 16178 27084
rect 11514 27044 11520 27056
rect 7966 27016 9996 27044
rect 10152 27016 11520 27044
rect 7966 27013 7978 27016
rect 7920 27007 7978 27013
rect 7466 26936 7472 26988
rect 7524 26976 7530 26988
rect 7653 26979 7711 26985
rect 7653 26976 7665 26979
rect 7524 26948 7665 26976
rect 7524 26936 7530 26948
rect 7653 26945 7665 26948
rect 7699 26945 7711 26979
rect 9858 26976 9864 26988
rect 9819 26948 9864 26976
rect 7653 26939 7711 26945
rect 9858 26936 9864 26948
rect 9916 26936 9922 26988
rect 9950 26936 9956 26988
rect 10008 26976 10014 26988
rect 10152 26985 10180 27016
rect 11514 27004 11520 27016
rect 11572 27004 11578 27056
rect 11685 27047 11743 27053
rect 11685 27013 11697 27047
rect 11731 27044 11743 27047
rect 11731 27016 11836 27044
rect 11731 27013 11743 27016
rect 11685 27007 11743 27013
rect 10137 26979 10195 26985
rect 10008 26948 10053 26976
rect 10008 26936 10014 26948
rect 10137 26945 10149 26979
rect 10183 26945 10195 26979
rect 10318 26976 10324 26988
rect 10279 26948 10324 26976
rect 10137 26939 10195 26945
rect 10318 26936 10324 26948
rect 10376 26936 10382 26988
rect 11808 26976 11836 27016
rect 11882 27004 11888 27056
rect 11940 27044 11946 27056
rect 18509 27047 18567 27053
rect 18509 27044 18521 27047
rect 11940 27016 14044 27044
rect 11940 27004 11946 27016
rect 12434 26976 12440 26988
rect 11808 26948 12440 26976
rect 12434 26936 12440 26948
rect 12492 26936 12498 26988
rect 12526 26936 12532 26988
rect 12584 26976 12590 26988
rect 14016 26985 14044 27016
rect 14200 27016 18521 27044
rect 14200 26985 14228 27016
rect 18509 27013 18521 27016
rect 18555 27013 18567 27047
rect 18616 27044 18644 27084
rect 18874 27072 18880 27124
rect 18932 27112 18938 27124
rect 18932 27084 18977 27112
rect 18932 27072 18938 27084
rect 19058 27072 19064 27124
rect 19116 27112 19122 27124
rect 19116 27084 19161 27112
rect 19116 27072 19122 27084
rect 19426 27072 19432 27124
rect 19484 27112 19490 27124
rect 19613 27115 19671 27121
rect 19613 27112 19625 27115
rect 19484 27084 19625 27112
rect 19484 27072 19490 27084
rect 19613 27081 19625 27084
rect 19659 27081 19671 27115
rect 19613 27075 19671 27081
rect 19702 27072 19708 27124
rect 19760 27112 19766 27124
rect 20622 27112 20628 27124
rect 19760 27084 20628 27112
rect 19760 27072 19766 27084
rect 20622 27072 20628 27084
rect 20680 27072 20686 27124
rect 19518 27044 19524 27056
rect 18616 27016 19524 27044
rect 18509 27007 18567 27013
rect 19518 27004 19524 27016
rect 19576 27004 19582 27056
rect 20806 27044 20812 27056
rect 20767 27016 20812 27044
rect 20806 27004 20812 27016
rect 20864 27004 20870 27056
rect 20990 27004 20996 27056
rect 21048 27044 21054 27056
rect 22557 27047 22615 27053
rect 22557 27044 22569 27047
rect 21048 27016 22569 27044
rect 21048 27004 21054 27016
rect 22557 27013 22569 27016
rect 22603 27044 22615 27047
rect 22646 27044 22652 27056
rect 22603 27016 22652 27044
rect 22603 27013 22615 27016
rect 22557 27007 22615 27013
rect 22646 27004 22652 27016
rect 22704 27004 22710 27056
rect 14001 26979 14059 26985
rect 12584 26948 12629 26976
rect 12584 26936 12590 26948
rect 14001 26945 14013 26979
rect 14047 26945 14059 26979
rect 14001 26939 14059 26945
rect 14185 26979 14243 26985
rect 14185 26945 14197 26979
rect 14231 26945 14243 26979
rect 14185 26939 14243 26945
rect 14016 26908 14044 26939
rect 14826 26936 14832 26988
rect 14884 26976 14890 26988
rect 14921 26979 14979 26985
rect 14921 26976 14933 26979
rect 14884 26948 14933 26976
rect 14884 26936 14890 26948
rect 14921 26945 14933 26948
rect 14967 26945 14979 26979
rect 14921 26939 14979 26945
rect 15286 26936 15292 26988
rect 15344 26976 15350 26988
rect 15565 26979 15623 26985
rect 15565 26976 15577 26979
rect 15344 26948 15577 26976
rect 15344 26936 15350 26948
rect 15565 26945 15577 26948
rect 15611 26945 15623 26979
rect 16666 26976 16672 26988
rect 16627 26948 16672 26976
rect 15565 26939 15623 26945
rect 16666 26936 16672 26948
rect 16724 26936 16730 26988
rect 16758 26936 16764 26988
rect 16816 26976 16822 26988
rect 16925 26979 16983 26985
rect 16925 26976 16937 26979
rect 16816 26948 16937 26976
rect 16816 26936 16822 26948
rect 16925 26945 16937 26948
rect 16971 26945 16983 26979
rect 16925 26939 16983 26945
rect 17494 26936 17500 26988
rect 17552 26976 17558 26988
rect 17954 26976 17960 26988
rect 17552 26948 17960 26976
rect 17552 26936 17558 26948
rect 17954 26936 17960 26948
rect 18012 26936 18018 26988
rect 18046 26936 18052 26988
rect 18104 26976 18110 26988
rect 19426 26976 19432 26988
rect 18104 26948 19432 26976
rect 18104 26936 18110 26948
rect 19426 26936 19432 26948
rect 19484 26936 19490 26988
rect 19797 26979 19855 26985
rect 19797 26976 19809 26979
rect 19720 26948 19809 26976
rect 14550 26908 14556 26920
rect 9048 26880 13952 26908
rect 14016 26880 14556 26908
rect 9048 26849 9076 26880
rect 9033 26843 9091 26849
rect 9033 26809 9045 26843
rect 9079 26809 9091 26843
rect 9033 26803 9091 26809
rect 10045 26843 10103 26849
rect 10045 26809 10057 26843
rect 10091 26840 10103 26843
rect 10134 26840 10140 26852
rect 10091 26812 10140 26840
rect 10091 26809 10103 26812
rect 10045 26803 10103 26809
rect 10134 26800 10140 26812
rect 10192 26840 10198 26852
rect 11790 26840 11796 26852
rect 10192 26812 11796 26840
rect 10192 26800 10198 26812
rect 11790 26800 11796 26812
rect 11848 26800 11854 26852
rect 13924 26840 13952 26880
rect 14550 26868 14556 26880
rect 14608 26868 14614 26920
rect 16114 26908 16120 26920
rect 14936 26880 16120 26908
rect 14936 26840 14964 26880
rect 16114 26868 16120 26880
rect 16172 26868 16178 26920
rect 18693 26911 18751 26917
rect 18693 26877 18705 26911
rect 18739 26877 18751 26911
rect 18693 26871 18751 26877
rect 13924 26812 14964 26840
rect 15105 26843 15163 26849
rect 15105 26809 15117 26843
rect 15151 26840 15163 26843
rect 16574 26840 16580 26852
rect 15151 26812 16580 26840
rect 15151 26809 15163 26812
rect 15105 26803 15163 26809
rect 16574 26800 16580 26812
rect 16632 26800 16638 26852
rect 18049 26843 18107 26849
rect 18049 26809 18061 26843
rect 18095 26840 18107 26843
rect 18230 26840 18236 26852
rect 18095 26812 18236 26840
rect 18095 26809 18107 26812
rect 18049 26803 18107 26809
rect 18230 26800 18236 26812
rect 18288 26840 18294 26852
rect 18708 26840 18736 26871
rect 18782 26868 18788 26920
rect 18840 26908 18846 26920
rect 19153 26911 19211 26917
rect 18840 26880 18885 26908
rect 18840 26868 18846 26880
rect 19153 26877 19165 26911
rect 19199 26908 19211 26911
rect 19242 26908 19248 26920
rect 19199 26880 19248 26908
rect 19199 26877 19211 26880
rect 19153 26871 19211 26877
rect 19242 26868 19248 26880
rect 19300 26868 19306 26920
rect 19610 26868 19616 26920
rect 19668 26908 19674 26920
rect 19720 26908 19748 26948
rect 19797 26945 19809 26948
rect 19843 26945 19855 26979
rect 22094 26976 22100 26988
rect 22055 26948 22100 26976
rect 19797 26939 19855 26945
rect 22094 26936 22100 26948
rect 22152 26936 22158 26988
rect 19878 26911 19936 26917
rect 19878 26908 19890 26911
rect 19668 26880 19748 26908
rect 19812 26880 19890 26908
rect 19668 26868 19674 26880
rect 19702 26840 19708 26852
rect 18288 26812 19708 26840
rect 18288 26800 18294 26812
rect 19702 26800 19708 26812
rect 19760 26840 19766 26852
rect 19812 26840 19840 26880
rect 19878 26877 19890 26880
rect 19924 26877 19936 26911
rect 19878 26871 19936 26877
rect 19981 26911 20039 26917
rect 19981 26877 19993 26911
rect 20027 26877 20039 26911
rect 19981 26871 20039 26877
rect 20073 26911 20131 26917
rect 20073 26877 20085 26911
rect 20119 26908 20131 26911
rect 20714 26908 20720 26920
rect 20119 26880 20720 26908
rect 20119 26877 20131 26880
rect 20073 26871 20131 26877
rect 19760 26812 19840 26840
rect 19760 26800 19766 26812
rect 9674 26732 9680 26784
rect 9732 26772 9738 26784
rect 11517 26775 11575 26781
rect 11517 26772 11529 26775
rect 9732 26744 11529 26772
rect 9732 26732 9738 26744
rect 11517 26741 11529 26744
rect 11563 26741 11575 26775
rect 11517 26735 11575 26741
rect 11701 26775 11759 26781
rect 11701 26741 11713 26775
rect 11747 26772 11759 26775
rect 11882 26772 11888 26784
rect 11747 26744 11888 26772
rect 11747 26741 11759 26744
rect 11701 26735 11759 26741
rect 11882 26732 11888 26744
rect 11940 26732 11946 26784
rect 13081 26775 13139 26781
rect 13081 26741 13093 26775
rect 13127 26772 13139 26775
rect 13170 26772 13176 26784
rect 13127 26744 13176 26772
rect 13127 26741 13139 26744
rect 13081 26735 13139 26741
rect 13170 26732 13176 26744
rect 13228 26732 13234 26784
rect 14826 26732 14832 26784
rect 14884 26772 14890 26784
rect 17770 26772 17776 26784
rect 14884 26744 17776 26772
rect 14884 26732 14890 26744
rect 17770 26732 17776 26744
rect 17828 26732 17834 26784
rect 19058 26732 19064 26784
rect 19116 26772 19122 26784
rect 19518 26772 19524 26784
rect 19116 26744 19524 26772
rect 19116 26732 19122 26744
rect 19518 26732 19524 26744
rect 19576 26772 19582 26784
rect 19996 26772 20024 26871
rect 20088 26784 20116 26871
rect 20714 26868 20720 26880
rect 20772 26908 20778 26920
rect 20772 26880 21220 26908
rect 20772 26868 20778 26880
rect 20530 26800 20536 26852
rect 20588 26840 20594 26852
rect 20806 26840 20812 26852
rect 20588 26812 20812 26840
rect 20588 26800 20594 26812
rect 20806 26800 20812 26812
rect 20864 26840 20870 26852
rect 20990 26840 20996 26852
rect 20864 26812 20996 26840
rect 20864 26800 20870 26812
rect 20990 26800 20996 26812
rect 21048 26840 21054 26852
rect 21085 26843 21143 26849
rect 21085 26840 21097 26843
rect 21048 26812 21097 26840
rect 21048 26800 21054 26812
rect 21085 26809 21097 26812
rect 21131 26809 21143 26843
rect 21192 26840 21220 26880
rect 21634 26868 21640 26920
rect 21692 26908 21698 26920
rect 21821 26911 21879 26917
rect 21821 26908 21833 26911
rect 21692 26880 21833 26908
rect 21692 26868 21698 26880
rect 21821 26877 21833 26880
rect 21867 26877 21879 26911
rect 21821 26871 21879 26877
rect 22005 26843 22063 26849
rect 22005 26840 22017 26843
rect 21192 26812 22017 26840
rect 21085 26803 21143 26809
rect 22005 26809 22017 26812
rect 22051 26809 22063 26843
rect 22005 26803 22063 26809
rect 19576 26744 20024 26772
rect 19576 26732 19582 26744
rect 20070 26732 20076 26784
rect 20128 26732 20134 26784
rect 21269 26775 21327 26781
rect 21269 26741 21281 26775
rect 21315 26772 21327 26775
rect 21358 26772 21364 26784
rect 21315 26744 21364 26772
rect 21315 26741 21327 26744
rect 21269 26735 21327 26741
rect 21358 26732 21364 26744
rect 21416 26732 21422 26784
rect 21634 26732 21640 26784
rect 21692 26772 21698 26784
rect 21913 26775 21971 26781
rect 21913 26772 21925 26775
rect 21692 26744 21925 26772
rect 21692 26732 21698 26744
rect 21913 26741 21925 26744
rect 21959 26741 21971 26775
rect 21913 26735 21971 26741
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 2774 26528 2780 26580
rect 2832 26568 2838 26580
rect 2832 26540 2877 26568
rect 2832 26528 2838 26540
rect 8294 26528 8300 26580
rect 8352 26568 8358 26580
rect 8941 26571 8999 26577
rect 8941 26568 8953 26571
rect 8352 26540 8953 26568
rect 8352 26528 8358 26540
rect 8941 26537 8953 26540
rect 8987 26537 8999 26571
rect 8941 26531 8999 26537
rect 9861 26571 9919 26577
rect 9861 26537 9873 26571
rect 9907 26568 9919 26571
rect 10042 26568 10048 26580
rect 9907 26540 10048 26568
rect 9907 26537 9919 26540
rect 9861 26531 9919 26537
rect 10042 26528 10048 26540
rect 10100 26528 10106 26580
rect 11882 26568 11888 26580
rect 11843 26540 11888 26568
rect 11882 26528 11888 26540
rect 11940 26528 11946 26580
rect 12526 26528 12532 26580
rect 12584 26568 12590 26580
rect 17862 26568 17868 26580
rect 12584 26540 17868 26568
rect 12584 26528 12590 26540
rect 17862 26528 17868 26540
rect 17920 26528 17926 26580
rect 18874 26528 18880 26580
rect 18932 26568 18938 26580
rect 19058 26568 19064 26580
rect 18932 26540 19064 26568
rect 18932 26528 18938 26540
rect 19058 26528 19064 26540
rect 19116 26568 19122 26580
rect 19521 26571 19579 26577
rect 19521 26568 19533 26571
rect 19116 26540 19533 26568
rect 19116 26528 19122 26540
rect 19521 26537 19533 26540
rect 19567 26537 19579 26571
rect 19521 26531 19579 26537
rect 19610 26528 19616 26580
rect 19668 26568 19674 26580
rect 19978 26568 19984 26580
rect 19668 26540 19984 26568
rect 19668 26528 19674 26540
rect 19978 26528 19984 26540
rect 20036 26568 20042 26580
rect 20349 26571 20407 26577
rect 20349 26568 20361 26571
rect 20036 26540 20361 26568
rect 20036 26528 20042 26540
rect 20349 26537 20361 26540
rect 20395 26568 20407 26571
rect 20530 26568 20536 26580
rect 20395 26540 20536 26568
rect 20395 26537 20407 26540
rect 20349 26531 20407 26537
rect 20530 26528 20536 26540
rect 20588 26528 20594 26580
rect 5353 26503 5411 26509
rect 5353 26469 5365 26503
rect 5399 26500 5411 26503
rect 15013 26503 15071 26509
rect 5399 26472 14964 26500
rect 5399 26469 5411 26472
rect 5353 26463 5411 26469
rect 1394 26432 1400 26444
rect 1355 26404 1400 26432
rect 1394 26392 1400 26404
rect 1452 26392 1458 26444
rect 4062 26432 4068 26444
rect 4023 26404 4068 26432
rect 4062 26392 4068 26404
rect 4120 26392 4126 26444
rect 11425 26435 11483 26441
rect 11425 26401 11437 26435
rect 11471 26432 11483 26435
rect 12897 26435 12955 26441
rect 12897 26432 12909 26435
rect 11471 26404 12909 26432
rect 11471 26401 11483 26404
rect 11425 26395 11483 26401
rect 1412 26364 1440 26392
rect 3789 26367 3847 26373
rect 3789 26364 3801 26367
rect 1412 26336 3801 26364
rect 3789 26333 3801 26336
rect 3835 26333 3847 26367
rect 3789 26327 3847 26333
rect 9217 26367 9275 26373
rect 9217 26333 9229 26367
rect 9263 26364 9275 26367
rect 9306 26364 9312 26376
rect 9263 26336 9312 26364
rect 9263 26333 9275 26336
rect 9217 26327 9275 26333
rect 9306 26324 9312 26336
rect 9364 26324 9370 26376
rect 9674 26364 9680 26376
rect 9635 26336 9680 26364
rect 9674 26324 9680 26336
rect 9732 26324 9738 26376
rect 12268 26373 12296 26404
rect 12897 26401 12909 26404
rect 12943 26432 12955 26435
rect 13538 26432 13544 26444
rect 12943 26404 13544 26432
rect 12943 26401 12955 26404
rect 12897 26395 12955 26401
rect 13538 26392 13544 26404
rect 13596 26432 13602 26444
rect 14461 26435 14519 26441
rect 14461 26432 14473 26435
rect 13596 26404 14473 26432
rect 13596 26392 13602 26404
rect 14461 26401 14473 26404
rect 14507 26401 14519 26435
rect 14936 26432 14964 26472
rect 15013 26469 15025 26503
rect 15059 26500 15071 26503
rect 15102 26500 15108 26512
rect 15059 26472 15108 26500
rect 15059 26469 15071 26472
rect 15013 26463 15071 26469
rect 15102 26460 15108 26472
rect 15160 26460 15166 26512
rect 16117 26503 16175 26509
rect 16117 26469 16129 26503
rect 16163 26500 16175 26503
rect 17034 26500 17040 26512
rect 16163 26472 17040 26500
rect 16163 26469 16175 26472
rect 16117 26463 16175 26469
rect 17034 26460 17040 26472
rect 17092 26460 17098 26512
rect 17310 26460 17316 26512
rect 17368 26500 17374 26512
rect 18506 26500 18512 26512
rect 17368 26472 18368 26500
rect 18467 26472 18512 26500
rect 17368 26460 17374 26472
rect 14936 26404 16620 26432
rect 14461 26395 14519 26401
rect 12069 26367 12127 26373
rect 12069 26333 12081 26367
rect 12115 26333 12127 26367
rect 12069 26327 12127 26333
rect 12253 26367 12311 26373
rect 12253 26333 12265 26367
rect 12299 26333 12311 26367
rect 12253 26327 12311 26333
rect 12345 26367 12403 26373
rect 12345 26333 12357 26367
rect 12391 26364 12403 26367
rect 13170 26364 13176 26376
rect 12391 26336 13176 26364
rect 12391 26333 12403 26336
rect 12345 26327 12403 26333
rect 1664 26299 1722 26305
rect 1664 26265 1676 26299
rect 1710 26296 1722 26299
rect 3878 26296 3884 26308
rect 1710 26268 3884 26296
rect 1710 26265 1722 26268
rect 1664 26259 1722 26265
rect 3878 26256 3884 26268
rect 3936 26256 3942 26308
rect 8938 26296 8944 26308
rect 8899 26268 8944 26296
rect 8938 26256 8944 26268
rect 8996 26256 9002 26308
rect 9125 26299 9183 26305
rect 9125 26265 9137 26299
rect 9171 26296 9183 26299
rect 9766 26296 9772 26308
rect 9171 26268 9772 26296
rect 9171 26265 9183 26268
rect 9125 26259 9183 26265
rect 9766 26256 9772 26268
rect 9824 26296 9830 26308
rect 10321 26299 10379 26305
rect 10321 26296 10333 26299
rect 9824 26268 10333 26296
rect 9824 26256 9830 26268
rect 10321 26265 10333 26268
rect 10367 26265 10379 26299
rect 12084 26296 12112 26327
rect 13170 26324 13176 26336
rect 13228 26324 13234 26376
rect 14826 26324 14832 26376
rect 14884 26364 14890 26376
rect 14884 26336 14929 26364
rect 14884 26324 14890 26336
rect 13078 26296 13084 26308
rect 12084 26268 13084 26296
rect 10321 26259 10379 26265
rect 13078 26256 13084 26268
rect 13136 26296 13142 26308
rect 13630 26296 13636 26308
rect 13136 26268 13636 26296
rect 13136 26256 13142 26268
rect 13630 26256 13636 26268
rect 13688 26296 13694 26308
rect 14737 26299 14795 26305
rect 14737 26296 14749 26299
rect 13688 26268 14412 26296
rect 13688 26256 13694 26268
rect 13538 26228 13544 26240
rect 13499 26200 13544 26228
rect 13538 26188 13544 26200
rect 13596 26188 13602 26240
rect 14384 26228 14412 26268
rect 14568 26268 14749 26296
rect 14568 26228 14596 26268
rect 14737 26265 14749 26268
rect 14783 26265 14795 26299
rect 15194 26296 15200 26308
rect 14737 26259 14795 26265
rect 14844 26268 15200 26296
rect 14384 26200 14596 26228
rect 14645 26231 14703 26237
rect 14645 26197 14657 26231
rect 14691 26228 14703 26231
rect 14844 26228 14872 26268
rect 15194 26256 15200 26268
rect 15252 26256 15258 26308
rect 16592 26296 16620 26404
rect 16666 26392 16672 26444
rect 16724 26432 16730 26444
rect 18049 26435 18107 26441
rect 18049 26432 18061 26435
rect 16724 26404 18061 26432
rect 16724 26392 16730 26404
rect 18049 26401 18061 26404
rect 18095 26401 18107 26435
rect 18340 26432 18368 26472
rect 18506 26460 18512 26472
rect 18564 26460 18570 26512
rect 19242 26460 19248 26512
rect 19300 26500 19306 26512
rect 19705 26503 19763 26509
rect 19300 26472 19580 26500
rect 19300 26460 19306 26472
rect 19334 26432 19340 26444
rect 18340 26404 19340 26432
rect 18049 26395 18107 26401
rect 19334 26392 19340 26404
rect 19392 26392 19398 26444
rect 19552 26432 19580 26472
rect 19705 26469 19717 26503
rect 19751 26469 19763 26503
rect 19705 26463 19763 26469
rect 19552 26404 19610 26432
rect 17034 26324 17040 26376
rect 17092 26364 17098 26376
rect 17092 26336 18092 26364
rect 17092 26324 17098 26336
rect 17310 26296 17316 26308
rect 16592 26268 17316 26296
rect 17310 26256 17316 26268
rect 17368 26256 17374 26308
rect 17405 26299 17463 26305
rect 17405 26265 17417 26299
rect 17451 26296 17463 26299
rect 17494 26296 17500 26308
rect 17451 26268 17500 26296
rect 17451 26265 17463 26268
rect 17405 26259 17463 26265
rect 17494 26256 17500 26268
rect 17552 26256 17558 26308
rect 17954 26296 17960 26308
rect 17915 26268 17960 26296
rect 17954 26256 17960 26268
rect 18012 26256 18018 26308
rect 18064 26237 18092 26336
rect 18782 26324 18788 26376
rect 18840 26364 18846 26376
rect 18840 26336 19334 26364
rect 19582 26339 19610 26404
rect 19720 26364 19748 26463
rect 21082 26460 21088 26512
rect 21140 26500 21146 26512
rect 21140 26472 21956 26500
rect 21140 26460 21146 26472
rect 21266 26392 21272 26444
rect 21324 26432 21330 26444
rect 21729 26435 21787 26441
rect 21729 26432 21741 26435
rect 21324 26404 21741 26432
rect 21324 26392 21330 26404
rect 21729 26401 21741 26404
rect 21775 26401 21787 26435
rect 21729 26395 21787 26401
rect 20257 26367 20315 26373
rect 20257 26364 20269 26367
rect 18840 26324 18846 26336
rect 19306 26330 19334 26336
rect 19567 26333 19625 26339
rect 19720 26336 20269 26364
rect 19306 26305 19380 26330
rect 19306 26302 19395 26305
rect 19337 26299 19395 26302
rect 19337 26265 19349 26299
rect 19383 26265 19395 26299
rect 19567 26299 19579 26333
rect 19613 26299 19625 26333
rect 20257 26333 20269 26336
rect 20303 26333 20315 26367
rect 21358 26364 21364 26376
rect 21319 26336 21364 26364
rect 20257 26327 20315 26333
rect 21358 26324 21364 26336
rect 21416 26324 21422 26376
rect 21634 26364 21640 26376
rect 21595 26336 21640 26364
rect 21634 26324 21640 26336
rect 21692 26324 21698 26376
rect 21928 26373 21956 26472
rect 21913 26367 21971 26373
rect 21913 26333 21925 26367
rect 21959 26333 21971 26367
rect 22094 26364 22100 26376
rect 22055 26336 22100 26364
rect 21913 26327 21971 26333
rect 22094 26324 22100 26336
rect 22152 26324 22158 26376
rect 22646 26364 22652 26376
rect 22607 26336 22652 26364
rect 22646 26324 22652 26336
rect 22704 26324 22710 26376
rect 19567 26293 19625 26299
rect 19337 26259 19395 26265
rect 14691 26200 14872 26228
rect 18049 26231 18107 26237
rect 14691 26197 14703 26200
rect 14645 26191 14703 26197
rect 18049 26197 18061 26231
rect 18095 26197 18107 26231
rect 18049 26191 18107 26197
rect 22002 26188 22008 26240
rect 22060 26228 22066 26240
rect 22833 26231 22891 26237
rect 22833 26228 22845 26231
rect 22060 26200 22845 26228
rect 22060 26188 22066 26200
rect 22833 26197 22845 26200
rect 22879 26197 22891 26231
rect 22833 26191 22891 26197
rect 1104 26138 38824 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 38824 26138
rect 1104 26064 38824 26086
rect 7837 26027 7895 26033
rect 7837 25993 7849 26027
rect 7883 25993 7895 26027
rect 12986 26024 12992 26036
rect 12947 25996 12992 26024
rect 7837 25987 7895 25993
rect 7852 25956 7880 25987
rect 12986 25984 12992 25996
rect 13044 25984 13050 26036
rect 15562 26024 15568 26036
rect 13924 25996 15568 26024
rect 8542 25959 8600 25965
rect 8542 25956 8554 25959
rect 7852 25928 8554 25956
rect 8542 25925 8554 25928
rect 8588 25925 8600 25959
rect 12250 25956 12256 25968
rect 8542 25919 8600 25925
rect 11624 25928 12256 25956
rect 7653 25891 7711 25897
rect 7653 25857 7665 25891
rect 7699 25888 7711 25891
rect 9490 25888 9496 25900
rect 7699 25860 9496 25888
rect 7699 25857 7711 25860
rect 7653 25851 7711 25857
rect 9490 25848 9496 25860
rect 9548 25848 9554 25900
rect 11624 25897 11652 25928
rect 12250 25916 12256 25928
rect 12308 25956 12314 25968
rect 12308 25928 13676 25956
rect 12308 25916 12314 25928
rect 11609 25891 11667 25897
rect 11609 25857 11621 25891
rect 11655 25857 11667 25891
rect 11609 25851 11667 25857
rect 11876 25891 11934 25897
rect 11876 25857 11888 25891
rect 11922 25888 11934 25891
rect 11922 25860 13308 25888
rect 11922 25857 11934 25860
rect 11876 25851 11934 25857
rect 7466 25780 7472 25832
rect 7524 25820 7530 25832
rect 8297 25823 8355 25829
rect 8297 25820 8309 25823
rect 7524 25792 8309 25820
rect 7524 25780 7530 25792
rect 8297 25789 8309 25792
rect 8343 25789 8355 25823
rect 8297 25783 8355 25789
rect 9674 25644 9680 25696
rect 9732 25684 9738 25696
rect 13280 25684 13308 25860
rect 13648 25752 13676 25928
rect 13814 25897 13820 25900
rect 13812 25888 13820 25897
rect 13775 25860 13820 25888
rect 13812 25851 13820 25860
rect 13814 25848 13820 25851
rect 13872 25848 13878 25900
rect 13924 25897 13952 25996
rect 15562 25984 15568 25996
rect 15620 25984 15626 26036
rect 17494 25984 17500 26036
rect 17552 26024 17558 26036
rect 18322 26024 18328 26036
rect 17552 25996 18328 26024
rect 17552 25984 17558 25996
rect 18322 25984 18328 25996
rect 18380 26024 18386 26036
rect 19061 26027 19119 26033
rect 19061 26024 19073 26027
rect 18380 25996 19073 26024
rect 18380 25984 18386 25996
rect 19061 25993 19073 25996
rect 19107 25993 19119 26027
rect 19061 25987 19119 25993
rect 20717 26027 20775 26033
rect 20717 25993 20729 26027
rect 20763 26024 20775 26027
rect 20806 26024 20812 26036
rect 20763 25996 20812 26024
rect 20763 25993 20775 25996
rect 20717 25987 20775 25993
rect 20806 25984 20812 25996
rect 20864 25984 20870 26036
rect 22094 25984 22100 26036
rect 22152 26024 22158 26036
rect 22189 26027 22247 26033
rect 22189 26024 22201 26027
rect 22152 25996 22201 26024
rect 22152 25984 22158 25996
rect 22189 25993 22201 25996
rect 22235 25993 22247 26027
rect 22189 25987 22247 25993
rect 16666 25956 16672 25968
rect 14752 25928 16672 25956
rect 13909 25891 13967 25897
rect 13909 25857 13921 25891
rect 13955 25857 13967 25891
rect 13909 25851 13967 25857
rect 13998 25848 14004 25900
rect 14056 25888 14062 25900
rect 14185 25891 14243 25897
rect 14056 25860 14101 25888
rect 14056 25848 14062 25860
rect 14185 25857 14197 25891
rect 14231 25888 14243 25891
rect 14458 25888 14464 25900
rect 14231 25860 14464 25888
rect 14231 25857 14243 25860
rect 14185 25851 14243 25857
rect 14458 25848 14464 25860
rect 14516 25848 14522 25900
rect 14752 25897 14780 25928
rect 16666 25916 16672 25928
rect 16724 25916 16730 25968
rect 17126 25956 17132 25968
rect 16868 25928 17132 25956
rect 15010 25897 15016 25900
rect 14737 25891 14795 25897
rect 14737 25857 14749 25891
rect 14783 25857 14795 25891
rect 14737 25851 14795 25857
rect 15004 25851 15016 25897
rect 15068 25888 15074 25900
rect 16868 25897 16896 25928
rect 17126 25916 17132 25928
rect 17184 25916 17190 25968
rect 19150 25916 19156 25968
rect 19208 25956 19214 25968
rect 21177 25959 21235 25965
rect 21177 25956 21189 25959
rect 19208 25928 21189 25956
rect 19208 25916 19214 25928
rect 21177 25925 21189 25928
rect 21223 25925 21235 25959
rect 21177 25919 21235 25925
rect 16853 25891 16911 25897
rect 15068 25860 15104 25888
rect 14752 25752 14780 25851
rect 15010 25848 15016 25851
rect 15068 25848 15074 25860
rect 16853 25857 16865 25891
rect 16899 25857 16911 25891
rect 17034 25888 17040 25900
rect 16995 25860 17040 25888
rect 16853 25851 16911 25857
rect 17034 25848 17040 25860
rect 17092 25848 17098 25900
rect 17773 25891 17831 25897
rect 17773 25857 17785 25891
rect 17819 25888 17831 25891
rect 18046 25888 18052 25900
rect 17819 25860 18052 25888
rect 17819 25857 17831 25860
rect 17773 25851 17831 25857
rect 18046 25848 18052 25860
rect 18104 25848 18110 25900
rect 20990 25848 20996 25900
rect 21048 25888 21054 25900
rect 21913 25891 21971 25897
rect 21913 25888 21925 25891
rect 21048 25860 21925 25888
rect 21048 25848 21054 25860
rect 21913 25857 21925 25860
rect 21959 25888 21971 25891
rect 22002 25888 22008 25900
rect 21959 25860 22008 25888
rect 21959 25857 21971 25860
rect 21913 25851 21971 25857
rect 22002 25848 22008 25860
rect 22060 25848 22066 25900
rect 22094 25848 22100 25900
rect 22152 25888 22158 25900
rect 22152 25860 22197 25888
rect 22152 25848 22158 25860
rect 13648 25724 14780 25752
rect 20073 25755 20131 25761
rect 20073 25721 20085 25755
rect 20119 25752 20131 25755
rect 20346 25752 20352 25764
rect 20119 25724 20352 25752
rect 20119 25721 20131 25724
rect 20073 25715 20131 25721
rect 20346 25712 20352 25724
rect 20404 25712 20410 25764
rect 14185 25687 14243 25693
rect 14185 25684 14197 25687
rect 9732 25656 9777 25684
rect 13280 25656 14197 25684
rect 9732 25644 9738 25656
rect 14185 25653 14197 25656
rect 14231 25653 14243 25687
rect 14185 25647 14243 25653
rect 14918 25644 14924 25696
rect 14976 25684 14982 25696
rect 16117 25687 16175 25693
rect 16117 25684 16129 25687
rect 14976 25656 16129 25684
rect 14976 25644 14982 25656
rect 16117 25653 16129 25656
rect 16163 25653 16175 25687
rect 16117 25647 16175 25653
rect 16850 25644 16856 25696
rect 16908 25684 16914 25696
rect 17037 25687 17095 25693
rect 17037 25684 17049 25687
rect 16908 25656 17049 25684
rect 16908 25644 16914 25656
rect 17037 25653 17049 25656
rect 17083 25653 17095 25687
rect 17037 25647 17095 25653
rect 20162 25644 20168 25696
rect 20220 25684 20226 25696
rect 20806 25684 20812 25696
rect 20220 25656 20812 25684
rect 20220 25644 20226 25656
rect 20806 25644 20812 25656
rect 20864 25644 20870 25696
rect 21726 25644 21732 25696
rect 21784 25684 21790 25696
rect 22373 25687 22431 25693
rect 22373 25684 22385 25687
rect 21784 25656 22385 25684
rect 21784 25644 21790 25656
rect 22373 25653 22385 25656
rect 22419 25653 22431 25687
rect 22373 25647 22431 25653
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 8938 25440 8944 25492
rect 8996 25480 9002 25492
rect 9401 25483 9459 25489
rect 9401 25480 9413 25483
rect 8996 25452 9413 25480
rect 8996 25440 9002 25452
rect 9401 25449 9413 25452
rect 9447 25449 9459 25483
rect 11422 25480 11428 25492
rect 11383 25452 11428 25480
rect 9401 25443 9459 25449
rect 11422 25440 11428 25452
rect 11480 25440 11486 25492
rect 12434 25440 12440 25492
rect 12492 25480 12498 25492
rect 13081 25483 13139 25489
rect 13081 25480 13093 25483
rect 12492 25452 13093 25480
rect 12492 25440 12498 25452
rect 13081 25449 13093 25452
rect 13127 25480 13139 25483
rect 13722 25480 13728 25492
rect 13127 25452 13728 25480
rect 13127 25449 13139 25452
rect 13081 25443 13139 25449
rect 13722 25440 13728 25452
rect 13780 25440 13786 25492
rect 13814 25440 13820 25492
rect 13872 25480 13878 25492
rect 14277 25483 14335 25489
rect 14277 25480 14289 25483
rect 13872 25452 14289 25480
rect 13872 25440 13878 25452
rect 14277 25449 14289 25452
rect 14323 25449 14335 25483
rect 14277 25443 14335 25449
rect 14550 25440 14556 25492
rect 14608 25480 14614 25492
rect 17126 25480 17132 25492
rect 14608 25452 17132 25480
rect 14608 25440 14614 25452
rect 17126 25440 17132 25452
rect 17184 25440 17190 25492
rect 17218 25440 17224 25492
rect 17276 25480 17282 25492
rect 17865 25483 17923 25489
rect 17865 25480 17877 25483
rect 17276 25452 17877 25480
rect 17276 25440 17282 25452
rect 17865 25449 17877 25452
rect 17911 25449 17923 25483
rect 17865 25443 17923 25449
rect 17954 25440 17960 25492
rect 18012 25480 18018 25492
rect 18012 25452 19334 25480
rect 18012 25440 18018 25452
rect 9306 25412 9312 25424
rect 9267 25384 9312 25412
rect 9306 25372 9312 25384
rect 9364 25372 9370 25424
rect 9674 25372 9680 25424
rect 9732 25412 9738 25424
rect 14642 25412 14648 25424
rect 9732 25384 14648 25412
rect 9732 25372 9738 25384
rect 14642 25372 14648 25384
rect 14700 25372 14706 25424
rect 19306 25412 19334 25452
rect 19426 25440 19432 25492
rect 19484 25480 19490 25492
rect 21726 25480 21732 25492
rect 19484 25452 21036 25480
rect 21687 25452 21732 25480
rect 19484 25440 19490 25452
rect 20441 25415 20499 25421
rect 20441 25412 20453 25415
rect 16316 25384 18368 25412
rect 19306 25384 20453 25412
rect 9493 25347 9551 25353
rect 9493 25313 9505 25347
rect 9539 25344 9551 25347
rect 10134 25344 10140 25356
rect 9539 25316 10140 25344
rect 9539 25313 9551 25316
rect 9493 25307 9551 25313
rect 10134 25304 10140 25316
rect 10192 25344 10198 25356
rect 10413 25347 10471 25353
rect 10413 25344 10425 25347
rect 10192 25316 10425 25344
rect 10192 25304 10198 25316
rect 10413 25313 10425 25316
rect 10459 25313 10471 25347
rect 10413 25307 10471 25313
rect 10597 25347 10655 25353
rect 10597 25313 10609 25347
rect 10643 25344 10655 25347
rect 10643 25316 11744 25344
rect 10643 25313 10655 25316
rect 10597 25307 10655 25313
rect 11716 25288 11744 25316
rect 11974 25304 11980 25356
rect 12032 25344 12038 25356
rect 16316 25353 16344 25384
rect 16301 25347 16359 25353
rect 12032 25316 15516 25344
rect 12032 25304 12038 25316
rect 9217 25279 9275 25285
rect 9217 25245 9229 25279
rect 9263 25276 9275 25279
rect 9766 25276 9772 25288
rect 9263 25248 9772 25276
rect 9263 25245 9275 25248
rect 9217 25239 9275 25245
rect 9766 25236 9772 25248
rect 9824 25236 9830 25288
rect 10689 25279 10747 25285
rect 10689 25245 10701 25279
rect 10735 25276 10747 25279
rect 11609 25279 11667 25285
rect 11609 25276 11621 25279
rect 10735 25248 11621 25276
rect 10735 25245 10747 25248
rect 10689 25239 10747 25245
rect 11609 25245 11621 25248
rect 11655 25245 11667 25279
rect 11609 25239 11667 25245
rect 10413 25211 10471 25217
rect 10413 25177 10425 25211
rect 10459 25208 10471 25211
rect 11425 25211 11483 25217
rect 11425 25208 11437 25211
rect 10459 25180 11437 25208
rect 10459 25177 10471 25180
rect 10413 25171 10471 25177
rect 11425 25177 11437 25180
rect 11471 25177 11483 25211
rect 11425 25171 11483 25177
rect 11624 25140 11652 25239
rect 11698 25236 11704 25288
rect 11756 25276 11762 25288
rect 12989 25279 13047 25285
rect 11756 25248 11801 25276
rect 11756 25236 11762 25248
rect 12989 25245 13001 25279
rect 13035 25276 13047 25279
rect 13078 25276 13084 25288
rect 13035 25248 13084 25276
rect 13035 25245 13047 25248
rect 12989 25239 13047 25245
rect 13078 25236 13084 25248
rect 13136 25236 13142 25288
rect 13265 25279 13323 25285
rect 13265 25245 13277 25279
rect 13311 25276 13323 25279
rect 13538 25276 13544 25288
rect 13311 25248 13544 25276
rect 13311 25245 13323 25248
rect 13265 25239 13323 25245
rect 13538 25236 13544 25248
rect 13596 25236 13602 25288
rect 13906 25236 13912 25288
rect 13964 25276 13970 25288
rect 14550 25276 14556 25288
rect 13964 25248 14556 25276
rect 13964 25236 13970 25248
rect 14550 25236 14556 25248
rect 14608 25236 14614 25288
rect 15488 25285 15516 25316
rect 16301 25313 16313 25347
rect 16347 25313 16359 25347
rect 18340 25344 18368 25384
rect 20441 25381 20453 25384
rect 20487 25381 20499 25415
rect 20714 25412 20720 25424
rect 20441 25375 20499 25381
rect 20548 25384 20720 25412
rect 19521 25347 19579 25353
rect 16301 25307 16359 25313
rect 16408 25316 18276 25344
rect 18340 25316 18404 25344
rect 15473 25279 15531 25285
rect 15473 25245 15485 25279
rect 15519 25245 15531 25279
rect 16022 25276 16028 25288
rect 15983 25248 16028 25276
rect 15473 25239 15531 25245
rect 16022 25236 16028 25248
rect 16080 25236 16086 25288
rect 16408 25285 16436 25316
rect 18248 25288 18276 25316
rect 16393 25279 16451 25285
rect 16393 25245 16405 25279
rect 16439 25245 16451 25279
rect 16393 25239 16451 25245
rect 16945 25279 17003 25285
rect 16945 25245 16957 25279
rect 16991 25245 17003 25279
rect 17310 25276 17316 25288
rect 17223 25248 17316 25276
rect 16945 25239 17003 25245
rect 12529 25211 12587 25217
rect 12529 25177 12541 25211
rect 12575 25208 12587 25211
rect 13170 25208 13176 25220
rect 12575 25180 13176 25208
rect 12575 25177 12587 25180
rect 12529 25171 12587 25177
rect 13170 25168 13176 25180
rect 13228 25208 13234 25220
rect 15194 25208 15200 25220
rect 13228 25180 15200 25208
rect 13228 25168 13234 25180
rect 15194 25168 15200 25180
rect 15252 25168 15258 25220
rect 16960 25208 16988 25239
rect 17310 25236 17316 25248
rect 17368 25276 17374 25288
rect 17880 25279 18087 25286
rect 17880 25276 18017 25279
rect 17368 25258 18017 25276
rect 17368 25248 17908 25258
rect 17368 25236 17374 25248
rect 18005 25245 18017 25258
rect 18051 25248 18087 25279
rect 18230 25276 18236 25288
rect 18191 25248 18236 25276
rect 18051 25245 18063 25248
rect 18005 25239 18063 25245
rect 18230 25236 18236 25248
rect 18288 25236 18294 25288
rect 18376 25285 18404 25316
rect 19521 25313 19533 25347
rect 19567 25344 19579 25347
rect 19794 25344 19800 25356
rect 19567 25316 19800 25344
rect 19567 25313 19579 25316
rect 19521 25307 19579 25313
rect 19794 25304 19800 25316
rect 19852 25304 19858 25356
rect 19889 25347 19947 25353
rect 19889 25313 19901 25347
rect 19935 25344 19947 25347
rect 20548 25344 20576 25384
rect 20714 25372 20720 25384
rect 20772 25372 20778 25424
rect 21008 25421 21036 25452
rect 21726 25440 21732 25452
rect 21784 25440 21790 25492
rect 20993 25415 21051 25421
rect 20993 25381 21005 25415
rect 21039 25412 21051 25415
rect 22094 25412 22100 25424
rect 21039 25384 22100 25412
rect 21039 25381 21051 25384
rect 20993 25375 21051 25381
rect 22094 25372 22100 25384
rect 22152 25372 22158 25424
rect 19935 25316 20576 25344
rect 19935 25313 19947 25316
rect 19889 25307 19947 25313
rect 18371 25279 18429 25285
rect 18371 25245 18383 25279
rect 18417 25245 18429 25279
rect 18371 25239 18429 25245
rect 18509 25279 18567 25285
rect 18509 25245 18521 25279
rect 18555 25276 18567 25279
rect 18598 25276 18604 25288
rect 18555 25248 18604 25276
rect 18555 25245 18567 25248
rect 18509 25239 18567 25245
rect 18141 25211 18199 25217
rect 16960 25180 17908 25208
rect 15378 25140 15384 25152
rect 11624 25112 15384 25140
rect 15378 25100 15384 25112
rect 15436 25100 15442 25152
rect 17880 25140 17908 25180
rect 18141 25177 18153 25211
rect 18187 25177 18199 25211
rect 18376 25208 18404 25239
rect 18598 25236 18604 25248
rect 18656 25236 18662 25288
rect 19426 25236 19432 25288
rect 19484 25276 19490 25288
rect 19613 25279 19671 25285
rect 19613 25276 19625 25279
rect 19484 25248 19625 25276
rect 19484 25236 19490 25248
rect 19613 25245 19625 25248
rect 19659 25245 19671 25279
rect 19613 25239 19671 25245
rect 19981 25279 20039 25285
rect 19981 25245 19993 25279
rect 20027 25276 20039 25279
rect 20530 25276 20536 25288
rect 20027 25248 20536 25276
rect 20027 25245 20039 25248
rect 19981 25239 20039 25245
rect 20530 25236 20536 25248
rect 20588 25236 20594 25288
rect 20622 25236 20628 25288
rect 20680 25236 20686 25288
rect 20714 25236 20720 25288
rect 20772 25276 20778 25288
rect 20772 25248 20817 25276
rect 20772 25236 20778 25248
rect 20162 25208 20168 25220
rect 18376 25180 20168 25208
rect 18141 25171 18199 25177
rect 18156 25140 18184 25171
rect 20162 25168 20168 25180
rect 20220 25168 20226 25220
rect 20254 25168 20260 25220
rect 20312 25208 20318 25220
rect 20640 25208 20668 25236
rect 20809 25211 20867 25217
rect 20809 25208 20821 25211
rect 20312 25180 20821 25208
rect 20312 25168 20318 25180
rect 20809 25177 20821 25180
rect 20855 25177 20867 25211
rect 20809 25171 20867 25177
rect 18690 25140 18696 25152
rect 17880 25112 18696 25140
rect 18690 25100 18696 25112
rect 18748 25100 18754 25152
rect 19337 25143 19395 25149
rect 19337 25109 19349 25143
rect 19383 25140 19395 25143
rect 19426 25140 19432 25152
rect 19383 25112 19432 25140
rect 19383 25109 19395 25112
rect 19337 25103 19395 25109
rect 19426 25100 19432 25112
rect 19484 25100 19490 25152
rect 19702 25140 19708 25152
rect 19663 25112 19708 25140
rect 19702 25100 19708 25112
rect 19760 25100 19766 25152
rect 19794 25100 19800 25152
rect 19852 25140 19858 25152
rect 20625 25143 20683 25149
rect 20625 25140 20637 25143
rect 19852 25112 20637 25140
rect 19852 25100 19858 25112
rect 20625 25109 20637 25112
rect 20671 25109 20683 25143
rect 20625 25103 20683 25109
rect 1104 25050 38824 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 38824 25050
rect 1104 24976 38824 24998
rect 9585 24939 9643 24945
rect 9585 24905 9597 24939
rect 9631 24936 9643 24939
rect 9766 24936 9772 24948
rect 9631 24908 9772 24936
rect 9631 24905 9643 24908
rect 9585 24899 9643 24905
rect 9766 24896 9772 24908
rect 9824 24896 9830 24948
rect 12342 24936 12348 24948
rect 12303 24908 12348 24936
rect 12342 24896 12348 24908
rect 12400 24896 12406 24948
rect 13538 24896 13544 24948
rect 13596 24936 13602 24948
rect 18046 24936 18052 24948
rect 13596 24908 14136 24936
rect 18007 24908 18052 24936
rect 13596 24896 13602 24908
rect 9784 24800 9812 24896
rect 13679 24837 13737 24843
rect 11701 24803 11759 24809
rect 11701 24800 11713 24803
rect 9784 24772 11713 24800
rect 11701 24769 11713 24772
rect 11747 24800 11759 24803
rect 11790 24800 11796 24812
rect 11747 24772 11796 24800
rect 11747 24769 11759 24772
rect 11701 24763 11759 24769
rect 11790 24760 11796 24772
rect 11848 24760 11854 24812
rect 12253 24803 12311 24809
rect 12253 24769 12265 24803
rect 12299 24769 12311 24803
rect 12253 24763 12311 24769
rect 9306 24692 9312 24744
rect 9364 24732 9370 24744
rect 12268 24732 12296 24763
rect 12526 24760 12532 24812
rect 12584 24800 12590 24812
rect 13679 24803 13691 24837
rect 13725 24834 13737 24837
rect 13725 24806 13860 24834
rect 13906 24828 13912 24880
rect 13964 24868 13970 24880
rect 14108 24868 14136 24908
rect 18046 24896 18052 24908
rect 18104 24896 18110 24948
rect 18138 24896 18144 24948
rect 18196 24936 18202 24948
rect 24213 24939 24271 24945
rect 24213 24936 24225 24939
rect 18196 24908 24225 24936
rect 18196 24896 18202 24908
rect 24213 24905 24225 24908
rect 24259 24905 24271 24939
rect 24213 24899 24271 24905
rect 17402 24868 17408 24880
rect 13964 24840 14009 24868
rect 14108 24840 17408 24868
rect 13964 24828 13970 24840
rect 17402 24828 17408 24840
rect 17460 24868 17466 24880
rect 19521 24871 19579 24877
rect 17460 24840 19334 24868
rect 17460 24828 17466 24840
rect 19306 24812 19334 24840
rect 19521 24837 19533 24871
rect 19567 24837 19579 24871
rect 19521 24834 19579 24837
rect 19521 24831 19656 24834
rect 13725 24803 13737 24806
rect 12584 24772 12629 24800
rect 13679 24797 13737 24803
rect 13832 24800 13860 24806
rect 14826 24800 14832 24812
rect 13832 24772 14832 24800
rect 12584 24760 12590 24772
rect 14826 24760 14832 24772
rect 14884 24760 14890 24812
rect 16666 24800 16672 24812
rect 16627 24772 16672 24800
rect 16666 24760 16672 24772
rect 16724 24760 16730 24812
rect 16942 24809 16948 24812
rect 16936 24763 16948 24809
rect 17000 24800 17006 24812
rect 17000 24772 17036 24800
rect 16942 24760 16948 24763
rect 17000 24760 17006 24772
rect 17310 24760 17316 24812
rect 17368 24800 17374 24812
rect 18138 24800 18144 24812
rect 17368 24772 18144 24800
rect 17368 24760 17374 24772
rect 18138 24760 18144 24772
rect 18196 24760 18202 24812
rect 19306 24778 19340 24812
rect 19334 24760 19340 24778
rect 19392 24760 19398 24812
rect 19429 24803 19487 24809
rect 19536 24806 19656 24831
rect 19886 24828 19892 24880
rect 19944 24868 19950 24880
rect 20162 24868 20168 24880
rect 19944 24840 20168 24868
rect 19944 24828 19950 24840
rect 20162 24828 20168 24840
rect 20220 24828 20226 24880
rect 21174 24828 21180 24880
rect 21232 24868 21238 24880
rect 21232 24840 24256 24868
rect 21232 24828 21238 24840
rect 19429 24769 19441 24803
rect 19475 24769 19487 24803
rect 19429 24763 19487 24769
rect 15102 24732 15108 24744
rect 9364 24704 15108 24732
rect 9364 24692 9370 24704
rect 15102 24692 15108 24704
rect 15160 24692 15166 24744
rect 19444 24732 19472 24763
rect 19518 24732 19524 24744
rect 18156 24704 19334 24732
rect 19444 24704 19524 24732
rect 9490 24624 9496 24676
rect 9548 24664 9554 24676
rect 13541 24667 13599 24673
rect 13541 24664 13553 24667
rect 9548 24636 13553 24664
rect 9548 24624 9554 24636
rect 13541 24633 13553 24636
rect 13587 24633 13599 24667
rect 13541 24627 13599 24633
rect 11790 24556 11796 24608
rect 11848 24596 11854 24608
rect 12434 24596 12440 24608
rect 11848 24568 12440 24596
rect 11848 24556 11854 24568
rect 12434 24556 12440 24568
rect 12492 24596 12498 24608
rect 12618 24596 12624 24608
rect 12492 24568 12624 24596
rect 12492 24556 12498 24568
rect 12618 24556 12624 24568
rect 12676 24556 12682 24608
rect 12713 24599 12771 24605
rect 12713 24565 12725 24599
rect 12759 24596 12771 24599
rect 13078 24596 13084 24608
rect 12759 24568 13084 24596
rect 12759 24565 12771 24568
rect 12713 24559 12771 24565
rect 13078 24556 13084 24568
rect 13136 24556 13142 24608
rect 13725 24599 13783 24605
rect 13725 24565 13737 24599
rect 13771 24596 13783 24599
rect 14090 24596 14096 24608
rect 13771 24568 14096 24596
rect 13771 24565 13783 24568
rect 13725 24559 13783 24565
rect 14090 24556 14096 24568
rect 14148 24556 14154 24608
rect 14274 24556 14280 24608
rect 14332 24596 14338 24608
rect 14369 24599 14427 24605
rect 14369 24596 14381 24599
rect 14332 24568 14381 24596
rect 14332 24556 14338 24568
rect 14369 24565 14381 24568
rect 14415 24565 14427 24599
rect 14369 24559 14427 24565
rect 14458 24556 14464 24608
rect 14516 24596 14522 24608
rect 18156 24596 18184 24704
rect 19306 24664 19334 24704
rect 19518 24692 19524 24704
rect 19576 24692 19582 24744
rect 19628 24664 19656 24806
rect 19705 24803 19763 24809
rect 19705 24769 19717 24803
rect 19751 24800 19763 24803
rect 20070 24800 20076 24812
rect 19751 24772 20076 24800
rect 19751 24769 19763 24772
rect 19705 24763 19763 24769
rect 20070 24760 20076 24772
rect 20128 24760 20134 24812
rect 20346 24800 20352 24812
rect 20307 24772 20352 24800
rect 20346 24760 20352 24772
rect 20404 24760 20410 24812
rect 20901 24803 20959 24809
rect 20901 24769 20913 24803
rect 20947 24800 20959 24803
rect 21910 24800 21916 24812
rect 20947 24772 21916 24800
rect 20947 24769 20959 24772
rect 20901 24763 20959 24769
rect 21910 24760 21916 24772
rect 21968 24760 21974 24812
rect 23658 24800 23664 24812
rect 23619 24772 23664 24800
rect 23658 24760 23664 24772
rect 23716 24760 23722 24812
rect 23752 24803 23810 24809
rect 23752 24769 23764 24803
rect 23798 24800 23810 24803
rect 23934 24800 23940 24812
rect 23798 24772 23940 24800
rect 23798 24769 23810 24772
rect 23752 24763 23810 24769
rect 23934 24760 23940 24772
rect 23992 24760 23998 24812
rect 24228 24809 24256 24840
rect 24213 24803 24271 24809
rect 24213 24769 24225 24803
rect 24259 24769 24271 24803
rect 24394 24800 24400 24812
rect 24355 24772 24400 24800
rect 24213 24763 24271 24769
rect 24394 24760 24400 24772
rect 24452 24760 24458 24812
rect 21085 24735 21143 24741
rect 21085 24732 21097 24735
rect 19720 24704 21097 24732
rect 19720 24673 19748 24704
rect 21085 24701 21097 24704
rect 21131 24701 21143 24735
rect 21085 24695 21143 24701
rect 21726 24692 21732 24744
rect 21784 24732 21790 24744
rect 22925 24735 22983 24741
rect 22925 24732 22937 24735
rect 21784 24704 22937 24732
rect 21784 24692 21790 24704
rect 22925 24701 22937 24704
rect 22971 24732 22983 24735
rect 23477 24735 23535 24741
rect 23477 24732 23489 24735
rect 22971 24704 23489 24732
rect 22971 24701 22983 24704
rect 22925 24695 22983 24701
rect 23477 24701 23489 24704
rect 23523 24701 23535 24735
rect 23477 24695 23535 24701
rect 19306 24636 19656 24664
rect 19705 24667 19763 24673
rect 19705 24633 19717 24667
rect 19751 24633 19763 24667
rect 19705 24627 19763 24633
rect 14516 24568 18184 24596
rect 18969 24599 19027 24605
rect 14516 24556 14522 24568
rect 18969 24565 18981 24599
rect 19015 24596 19027 24599
rect 19058 24596 19064 24608
rect 19015 24568 19064 24596
rect 19015 24565 19027 24568
rect 18969 24559 19027 24565
rect 19058 24556 19064 24568
rect 19116 24556 19122 24608
rect 22002 24596 22008 24608
rect 21963 24568 22008 24596
rect 22002 24556 22008 24568
rect 22060 24556 22066 24608
rect 23382 24556 23388 24608
rect 23440 24596 23446 24608
rect 23569 24599 23627 24605
rect 23569 24596 23581 24599
rect 23440 24568 23581 24596
rect 23440 24556 23446 24568
rect 23569 24565 23581 24568
rect 23615 24565 23627 24599
rect 23569 24559 23627 24565
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 13538 24392 13544 24404
rect 13499 24364 13544 24392
rect 13538 24352 13544 24364
rect 13596 24352 13602 24404
rect 14090 24392 14096 24404
rect 14051 24364 14096 24392
rect 14090 24352 14096 24364
rect 14148 24352 14154 24404
rect 16942 24392 16948 24404
rect 16903 24364 16948 24392
rect 16942 24352 16948 24364
rect 17000 24352 17006 24404
rect 17862 24352 17868 24404
rect 17920 24392 17926 24404
rect 18233 24395 18291 24401
rect 18233 24392 18245 24395
rect 17920 24364 18245 24392
rect 17920 24352 17926 24364
rect 18233 24361 18245 24364
rect 18279 24361 18291 24395
rect 18233 24355 18291 24361
rect 18417 24395 18475 24401
rect 18417 24361 18429 24395
rect 18463 24392 18475 24395
rect 19334 24392 19340 24404
rect 18463 24364 19340 24392
rect 18463 24361 18475 24364
rect 18417 24355 18475 24361
rect 19334 24352 19340 24364
rect 19392 24352 19398 24404
rect 20070 24392 20076 24404
rect 20031 24364 20076 24392
rect 20070 24352 20076 24364
rect 20128 24352 20134 24404
rect 20809 24395 20867 24401
rect 20809 24361 20821 24395
rect 20855 24392 20867 24395
rect 21726 24392 21732 24404
rect 20855 24364 21732 24392
rect 20855 24361 20867 24364
rect 20809 24355 20867 24361
rect 12437 24327 12495 24333
rect 12437 24293 12449 24327
rect 12483 24324 12495 24327
rect 12526 24324 12532 24336
rect 12483 24296 12532 24324
rect 12483 24293 12495 24296
rect 12437 24287 12495 24293
rect 12526 24284 12532 24296
rect 12584 24324 12590 24336
rect 13354 24324 13360 24336
rect 12584 24296 13360 24324
rect 12584 24284 12590 24296
rect 13354 24284 13360 24296
rect 13412 24324 13418 24336
rect 13412 24296 15240 24324
rect 13412 24284 13418 24296
rect 13906 24256 13912 24268
rect 12912 24228 13912 24256
rect 12912 24197 12940 24228
rect 13906 24216 13912 24228
rect 13964 24216 13970 24268
rect 12897 24191 12955 24197
rect 12897 24157 12909 24191
rect 12943 24157 12955 24191
rect 13078 24188 13084 24200
rect 13039 24160 13084 24188
rect 12897 24151 12955 24157
rect 13078 24148 13084 24160
rect 13136 24148 13142 24200
rect 13170 24148 13176 24200
rect 13228 24188 13234 24200
rect 13311 24191 13369 24197
rect 13228 24160 13273 24188
rect 13228 24148 13234 24160
rect 13311 24157 13323 24191
rect 13357 24188 13369 24191
rect 13722 24188 13728 24200
rect 13357 24160 13728 24188
rect 13357 24157 13369 24160
rect 13311 24151 13369 24157
rect 13722 24148 13728 24160
rect 13780 24148 13786 24200
rect 14200 24188 14228 24296
rect 14277 24259 14335 24265
rect 14277 24225 14289 24259
rect 14323 24256 14335 24259
rect 15102 24256 15108 24268
rect 14323 24228 15108 24256
rect 14323 24225 14335 24228
rect 14277 24219 14335 24225
rect 15102 24216 15108 24228
rect 15160 24216 15166 24268
rect 15212 24265 15240 24296
rect 17586 24284 17592 24336
rect 17644 24324 17650 24336
rect 20165 24327 20223 24333
rect 20165 24324 20177 24327
rect 17644 24296 20177 24324
rect 17644 24284 17650 24296
rect 20165 24293 20177 24296
rect 20211 24293 20223 24327
rect 20165 24287 20223 24293
rect 15197 24259 15255 24265
rect 15197 24225 15209 24259
rect 15243 24256 15255 24259
rect 18414 24256 18420 24268
rect 15243 24228 18420 24256
rect 15243 24225 15255 24228
rect 15197 24219 15255 24225
rect 18414 24216 18420 24228
rect 18472 24256 18478 24268
rect 18874 24256 18880 24268
rect 18472 24228 18880 24256
rect 18472 24216 18478 24228
rect 18874 24216 18880 24228
rect 18932 24216 18938 24268
rect 19981 24259 20039 24265
rect 19981 24225 19993 24259
rect 20027 24256 20039 24259
rect 20824 24256 20852 24355
rect 21726 24352 21732 24364
rect 21784 24352 21790 24404
rect 23385 24395 23443 24401
rect 21928 24364 22416 24392
rect 20898 24284 20904 24336
rect 20956 24324 20962 24336
rect 21545 24327 21603 24333
rect 21545 24324 21557 24327
rect 20956 24296 21557 24324
rect 20956 24284 20962 24296
rect 21545 24293 21557 24296
rect 21591 24324 21603 24327
rect 21928 24324 21956 24364
rect 22388 24336 22416 24364
rect 23385 24361 23397 24395
rect 23431 24392 23443 24395
rect 24394 24392 24400 24404
rect 23431 24364 24400 24392
rect 23431 24361 23443 24364
rect 23385 24355 23443 24361
rect 24394 24352 24400 24364
rect 24452 24352 24458 24404
rect 21591 24296 21956 24324
rect 21591 24293 21603 24296
rect 21545 24287 21603 24293
rect 22002 24284 22008 24336
rect 22060 24324 22066 24336
rect 22370 24324 22376 24336
rect 22060 24296 22140 24324
rect 22283 24296 22376 24324
rect 22060 24284 22066 24296
rect 22112 24265 22140 24296
rect 22370 24284 22376 24296
rect 22428 24284 22434 24336
rect 22557 24327 22615 24333
rect 22557 24293 22569 24327
rect 22603 24324 22615 24327
rect 23474 24324 23480 24336
rect 22603 24296 23480 24324
rect 22603 24293 22615 24296
rect 22557 24287 22615 24293
rect 23474 24284 23480 24296
rect 23532 24284 23538 24336
rect 20027 24228 20852 24256
rect 22097 24259 22155 24265
rect 20027 24225 20039 24228
rect 19981 24219 20039 24225
rect 22097 24225 22109 24259
rect 22143 24225 22155 24259
rect 23382 24256 23388 24268
rect 23343 24228 23388 24256
rect 22097 24219 22155 24225
rect 23382 24216 23388 24228
rect 23440 24216 23446 24268
rect 14369 24191 14427 24197
rect 14369 24188 14381 24191
rect 14200 24160 14381 24188
rect 14369 24157 14381 24160
rect 14415 24157 14427 24191
rect 14369 24151 14427 24157
rect 14461 24191 14519 24197
rect 14461 24157 14473 24191
rect 14507 24157 14519 24191
rect 14461 24151 14519 24157
rect 14553 24191 14611 24197
rect 14553 24157 14565 24191
rect 14599 24188 14611 24191
rect 14642 24188 14648 24200
rect 14599 24160 14648 24188
rect 14599 24157 14611 24160
rect 14553 24151 14611 24157
rect 12618 24080 12624 24132
rect 12676 24120 12682 24132
rect 13446 24120 13452 24132
rect 12676 24092 13452 24120
rect 12676 24080 12682 24092
rect 13446 24080 13452 24092
rect 13504 24120 13510 24132
rect 14274 24120 14280 24132
rect 13504 24092 14280 24120
rect 13504 24080 13510 24092
rect 14274 24080 14280 24092
rect 14332 24120 14338 24132
rect 14476 24120 14504 24151
rect 14642 24148 14648 24160
rect 14700 24148 14706 24200
rect 16850 24188 16856 24200
rect 16811 24160 16856 24188
rect 16850 24148 16856 24160
rect 16908 24148 16914 24200
rect 17126 24188 17132 24200
rect 17087 24160 17132 24188
rect 17126 24148 17132 24160
rect 17184 24148 17190 24200
rect 17236 24160 18736 24188
rect 17236 24120 17264 24160
rect 14332 24092 17264 24120
rect 14332 24080 14338 24092
rect 18138 24080 18144 24132
rect 18196 24120 18202 24132
rect 18601 24123 18659 24129
rect 18601 24120 18613 24123
rect 18196 24092 18613 24120
rect 18196 24080 18202 24092
rect 18601 24089 18613 24092
rect 18647 24089 18659 24123
rect 18708 24120 18736 24160
rect 19518 24148 19524 24200
rect 19576 24188 19582 24200
rect 20257 24191 20315 24197
rect 20257 24188 20269 24191
rect 19576 24160 20269 24188
rect 19576 24148 19582 24160
rect 20257 24157 20269 24160
rect 20303 24188 20315 24191
rect 20990 24188 20996 24200
rect 20303 24160 20996 24188
rect 20303 24157 20315 24160
rect 20257 24151 20315 24157
rect 20990 24148 20996 24160
rect 21048 24148 21054 24200
rect 23566 24188 23572 24200
rect 23527 24160 23572 24188
rect 23566 24148 23572 24160
rect 23624 24148 23630 24200
rect 20806 24120 20812 24132
rect 18708 24092 20812 24120
rect 18601 24083 18659 24089
rect 20806 24080 20812 24092
rect 20864 24080 20870 24132
rect 23198 24120 23204 24132
rect 23159 24092 23204 24120
rect 23198 24080 23204 24092
rect 23256 24080 23262 24132
rect 18414 24061 18420 24064
rect 18401 24055 18420 24061
rect 18401 24021 18413 24055
rect 18401 24015 18420 24021
rect 18414 24012 18420 24015
rect 18472 24012 18478 24064
rect 19150 24012 19156 24064
rect 19208 24052 19214 24064
rect 19337 24055 19395 24061
rect 19337 24052 19349 24055
rect 19208 24024 19349 24052
rect 19208 24012 19214 24024
rect 19337 24021 19349 24024
rect 19383 24052 19395 24055
rect 19426 24052 19432 24064
rect 19383 24024 19432 24052
rect 19383 24021 19395 24024
rect 19337 24015 19395 24021
rect 19426 24012 19432 24024
rect 19484 24012 19490 24064
rect 19610 24012 19616 24064
rect 19668 24052 19674 24064
rect 24302 24052 24308 24064
rect 19668 24024 24308 24052
rect 19668 24012 19674 24024
rect 24302 24012 24308 24024
rect 24360 24052 24366 24064
rect 24397 24055 24455 24061
rect 24397 24052 24409 24055
rect 24360 24024 24409 24052
rect 24360 24012 24366 24024
rect 24397 24021 24409 24024
rect 24443 24021 24455 24055
rect 24397 24015 24455 24021
rect 1104 23962 38824 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 38824 23962
rect 1104 23888 38824 23910
rect 13170 23808 13176 23860
rect 13228 23848 13234 23860
rect 13265 23851 13323 23857
rect 13265 23848 13277 23851
rect 13228 23820 13277 23848
rect 13228 23808 13234 23820
rect 13265 23817 13277 23820
rect 13311 23848 13323 23851
rect 13311 23820 13952 23848
rect 13311 23817 13323 23820
rect 13265 23811 13323 23817
rect 13446 23780 13452 23792
rect 13188 23752 13452 23780
rect 12989 23715 13047 23721
rect 12989 23681 13001 23715
rect 13035 23712 13047 23715
rect 13078 23712 13084 23724
rect 13035 23684 13084 23712
rect 13035 23681 13047 23684
rect 12989 23675 13047 23681
rect 13078 23672 13084 23684
rect 13136 23672 13142 23724
rect 13188 23721 13216 23752
rect 13446 23740 13452 23752
rect 13504 23740 13510 23792
rect 13814 23780 13820 23792
rect 13556 23752 13820 23780
rect 13173 23715 13231 23721
rect 13173 23681 13185 23715
rect 13219 23681 13231 23715
rect 13173 23675 13231 23681
rect 13265 23715 13323 23721
rect 13265 23681 13277 23715
rect 13311 23712 13323 23715
rect 13556 23712 13584 23752
rect 13814 23740 13820 23752
rect 13872 23740 13878 23792
rect 13722 23712 13728 23724
rect 13311 23684 13584 23712
rect 13683 23684 13728 23712
rect 13311 23681 13323 23684
rect 13265 23675 13323 23681
rect 13722 23672 13728 23684
rect 13780 23672 13786 23724
rect 13924 23721 13952 23820
rect 14182 23808 14188 23860
rect 14240 23848 14246 23860
rect 15197 23851 15255 23857
rect 15197 23848 15209 23851
rect 14240 23820 15209 23848
rect 14240 23808 14246 23820
rect 15197 23817 15209 23820
rect 15243 23817 15255 23851
rect 15197 23811 15255 23817
rect 16761 23851 16819 23857
rect 16761 23817 16773 23851
rect 16807 23848 16819 23851
rect 17034 23848 17040 23860
rect 16807 23820 17040 23848
rect 16807 23817 16819 23820
rect 16761 23811 16819 23817
rect 17034 23808 17040 23820
rect 17092 23808 17098 23860
rect 17773 23851 17831 23857
rect 17773 23817 17785 23851
rect 17819 23848 17831 23851
rect 18414 23848 18420 23860
rect 17819 23820 18420 23848
rect 17819 23817 17831 23820
rect 17773 23811 17831 23817
rect 18414 23808 18420 23820
rect 18472 23808 18478 23860
rect 18598 23808 18604 23860
rect 18656 23848 18662 23860
rect 19521 23851 19579 23857
rect 19521 23848 19533 23851
rect 18656 23820 19533 23848
rect 18656 23808 18662 23820
rect 19521 23817 19533 23820
rect 19567 23817 19579 23851
rect 19521 23811 19579 23817
rect 20533 23851 20591 23857
rect 20533 23817 20545 23851
rect 20579 23848 20591 23851
rect 20898 23848 20904 23860
rect 20579 23820 20904 23848
rect 20579 23817 20591 23820
rect 20533 23811 20591 23817
rect 17954 23780 17960 23792
rect 17604 23752 17960 23780
rect 13909 23715 13967 23721
rect 13909 23681 13921 23715
rect 13955 23681 13967 23715
rect 13909 23675 13967 23681
rect 15013 23715 15071 23721
rect 15013 23681 15025 23715
rect 15059 23712 15071 23715
rect 15746 23712 15752 23724
rect 15059 23684 15752 23712
rect 15059 23681 15071 23684
rect 15013 23675 15071 23681
rect 15746 23672 15752 23684
rect 15804 23672 15810 23724
rect 16574 23672 16580 23724
rect 16632 23712 16638 23724
rect 17604 23721 17632 23752
rect 17954 23740 17960 23752
rect 18012 23740 18018 23792
rect 18233 23783 18291 23789
rect 18233 23749 18245 23783
rect 18279 23780 18291 23783
rect 18322 23780 18328 23792
rect 18279 23752 18328 23780
rect 18279 23749 18291 23752
rect 18233 23743 18291 23749
rect 18322 23740 18328 23752
rect 18380 23740 18386 23792
rect 19058 23740 19064 23792
rect 19116 23780 19122 23792
rect 20548 23780 20576 23811
rect 20898 23808 20904 23820
rect 20956 23808 20962 23860
rect 21910 23848 21916 23860
rect 21871 23820 21916 23848
rect 21910 23808 21916 23820
rect 21968 23808 21974 23860
rect 19116 23752 20576 23780
rect 19116 23740 19122 23752
rect 20990 23740 20996 23792
rect 21048 23780 21054 23792
rect 22186 23780 22192 23792
rect 21048 23752 22192 23780
rect 21048 23740 21054 23752
rect 22186 23740 22192 23752
rect 22244 23780 22250 23792
rect 23934 23780 23940 23792
rect 22244 23752 23940 23780
rect 22244 23740 22250 23752
rect 16945 23715 17003 23721
rect 16945 23712 16957 23715
rect 16632 23684 16957 23712
rect 16632 23672 16638 23684
rect 16945 23681 16957 23684
rect 16991 23681 17003 23715
rect 16945 23675 17003 23681
rect 17589 23715 17647 23721
rect 17589 23681 17601 23715
rect 17635 23681 17647 23715
rect 17589 23675 17647 23681
rect 17678 23672 17684 23724
rect 17736 23712 17742 23724
rect 17773 23715 17831 23721
rect 17773 23712 17785 23715
rect 17736 23684 17785 23712
rect 17736 23672 17742 23684
rect 17773 23681 17785 23684
rect 17819 23681 17831 23715
rect 17773 23675 17831 23681
rect 21269 23715 21327 23721
rect 21269 23681 21281 23715
rect 21315 23712 21327 23715
rect 21726 23712 21732 23724
rect 21315 23684 21732 23712
rect 21315 23681 21327 23684
rect 21269 23675 21327 23681
rect 21726 23672 21732 23684
rect 21784 23712 21790 23724
rect 22005 23715 22063 23721
rect 22005 23712 22017 23715
rect 21784 23684 22017 23712
rect 21784 23672 21790 23684
rect 22005 23681 22017 23684
rect 22051 23681 22063 23715
rect 22278 23712 22284 23724
rect 22239 23684 22284 23712
rect 22005 23675 22063 23681
rect 22278 23672 22284 23684
rect 22336 23672 22342 23724
rect 22572 23721 22600 23752
rect 23934 23740 23940 23752
rect 23992 23780 23998 23792
rect 23992 23752 24164 23780
rect 23992 23740 23998 23752
rect 22557 23715 22615 23721
rect 22557 23681 22569 23715
rect 22603 23681 22615 23715
rect 22557 23675 22615 23681
rect 23198 23672 23204 23724
rect 23256 23712 23262 23724
rect 23293 23715 23351 23721
rect 23293 23712 23305 23715
rect 23256 23684 23305 23712
rect 23256 23672 23262 23684
rect 23293 23681 23305 23684
rect 23339 23681 23351 23715
rect 23293 23675 23351 23681
rect 23382 23672 23388 23724
rect 23440 23712 23446 23724
rect 23440 23684 23485 23712
rect 23440 23672 23446 23684
rect 23566 23672 23572 23724
rect 23624 23712 23630 23724
rect 24136 23721 24164 23752
rect 23661 23715 23719 23721
rect 23661 23712 23673 23715
rect 23624 23684 23673 23712
rect 23624 23672 23630 23684
rect 23661 23681 23673 23684
rect 23707 23681 23719 23715
rect 23661 23675 23719 23681
rect 24121 23715 24179 23721
rect 24121 23681 24133 23715
rect 24167 23681 24179 23715
rect 24302 23712 24308 23724
rect 24263 23684 24308 23712
rect 24121 23675 24179 23681
rect 10318 23604 10324 23656
rect 10376 23644 10382 23656
rect 14829 23647 14887 23653
rect 14829 23644 14841 23647
rect 10376 23616 14841 23644
rect 10376 23604 10382 23616
rect 14829 23613 14841 23616
rect 14875 23613 14887 23647
rect 14829 23607 14887 23613
rect 17126 23604 17132 23656
rect 17184 23644 17190 23656
rect 17696 23644 17724 23672
rect 17184 23616 17724 23644
rect 17184 23604 17190 23616
rect 20714 23604 20720 23656
rect 20772 23644 20778 23656
rect 21821 23647 21879 23653
rect 21821 23644 21833 23647
rect 20772 23616 21833 23644
rect 20772 23604 20778 23616
rect 21821 23613 21833 23616
rect 21867 23613 21879 23647
rect 23676 23644 23704 23675
rect 24302 23672 24308 23684
rect 24360 23672 24366 23724
rect 23676 23616 24348 23644
rect 21821 23607 21879 23613
rect 12529 23579 12587 23585
rect 12529 23545 12541 23579
rect 12575 23576 12587 23579
rect 13814 23576 13820 23588
rect 12575 23548 13820 23576
rect 12575 23545 12587 23548
rect 12529 23539 12587 23545
rect 13814 23536 13820 23548
rect 13872 23536 13878 23588
rect 14001 23579 14059 23585
rect 14001 23545 14013 23579
rect 14047 23576 14059 23579
rect 15010 23576 15016 23588
rect 14047 23548 15016 23576
rect 14047 23545 14059 23548
rect 14001 23539 14059 23545
rect 15010 23536 15016 23548
rect 15068 23536 15074 23588
rect 15194 23536 15200 23588
rect 15252 23576 15258 23588
rect 22002 23576 22008 23588
rect 15252 23548 22008 23576
rect 15252 23536 15258 23548
rect 22002 23536 22008 23548
rect 22060 23536 22066 23588
rect 23474 23536 23480 23588
rect 23532 23576 23538 23588
rect 24320 23585 24348 23616
rect 23569 23579 23627 23585
rect 23569 23576 23581 23579
rect 23532 23548 23581 23576
rect 23532 23536 23538 23548
rect 23569 23545 23581 23548
rect 23615 23545 23627 23579
rect 23569 23539 23627 23545
rect 24305 23579 24363 23585
rect 24305 23545 24317 23579
rect 24351 23545 24363 23579
rect 24305 23539 24363 23545
rect 15746 23508 15752 23520
rect 15707 23480 15752 23508
rect 15746 23468 15752 23480
rect 15804 23468 15810 23520
rect 16850 23468 16856 23520
rect 16908 23508 16914 23520
rect 19242 23508 19248 23520
rect 16908 23480 19248 23508
rect 16908 23468 16914 23480
rect 19242 23468 19248 23480
rect 19300 23468 19306 23520
rect 23106 23508 23112 23520
rect 23067 23480 23112 23508
rect 23106 23468 23112 23480
rect 23164 23468 23170 23520
rect 24578 23508 24584 23520
rect 24539 23480 24584 23508
rect 24578 23468 24584 23480
rect 24636 23468 24642 23520
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 12713 23307 12771 23313
rect 12713 23273 12725 23307
rect 12759 23304 12771 23307
rect 13446 23304 13452 23316
rect 12759 23276 13452 23304
rect 12759 23273 12771 23276
rect 12713 23267 12771 23273
rect 13446 23264 13452 23276
rect 13504 23264 13510 23316
rect 15105 23307 15163 23313
rect 15105 23273 15117 23307
rect 15151 23304 15163 23307
rect 15749 23307 15807 23313
rect 15749 23304 15761 23307
rect 15151 23276 15761 23304
rect 15151 23273 15163 23276
rect 15105 23267 15163 23273
rect 15749 23273 15761 23276
rect 15795 23273 15807 23307
rect 15749 23267 15807 23273
rect 15838 23264 15844 23316
rect 15896 23304 15902 23316
rect 16761 23307 16819 23313
rect 16761 23304 16773 23307
rect 15896 23276 16773 23304
rect 15896 23264 15902 23276
rect 16761 23273 16773 23276
rect 16807 23273 16819 23307
rect 16761 23267 16819 23273
rect 17402 23264 17408 23316
rect 17460 23304 17466 23316
rect 17957 23307 18015 23313
rect 17957 23304 17969 23307
rect 17460 23276 17969 23304
rect 17460 23264 17466 23276
rect 17957 23273 17969 23276
rect 18003 23273 18015 23307
rect 19337 23307 19395 23313
rect 19337 23304 19349 23307
rect 17957 23267 18015 23273
rect 18984 23276 19349 23304
rect 13354 23236 13360 23248
rect 13315 23208 13360 23236
rect 13354 23196 13360 23208
rect 13412 23196 13418 23248
rect 15286 23236 15292 23248
rect 15247 23208 15292 23236
rect 15286 23196 15292 23208
rect 15344 23196 15350 23248
rect 15378 23196 15384 23248
rect 15436 23236 15442 23248
rect 17310 23236 17316 23248
rect 15436 23208 16160 23236
rect 17271 23208 17316 23236
rect 15436 23196 15442 23208
rect 11698 23128 11704 23180
rect 11756 23168 11762 23180
rect 15838 23168 15844 23180
rect 11756 23140 15844 23168
rect 11756 23128 11762 23140
rect 15838 23128 15844 23140
rect 15896 23168 15902 23180
rect 16132 23177 16160 23208
rect 17310 23196 17316 23208
rect 17368 23196 17374 23248
rect 17770 23236 17776 23248
rect 17731 23208 17776 23236
rect 17770 23196 17776 23208
rect 17828 23196 17834 23248
rect 17862 23196 17868 23248
rect 17920 23236 17926 23248
rect 18984 23236 19012 23276
rect 19337 23273 19349 23276
rect 19383 23304 19395 23307
rect 19426 23304 19432 23316
rect 19383 23276 19432 23304
rect 19383 23273 19395 23276
rect 19337 23267 19395 23273
rect 19426 23264 19432 23276
rect 19484 23264 19490 23316
rect 20533 23307 20591 23313
rect 20533 23273 20545 23307
rect 20579 23304 20591 23307
rect 20714 23304 20720 23316
rect 20579 23276 20720 23304
rect 20579 23273 20591 23276
rect 20533 23267 20591 23273
rect 20714 23264 20720 23276
rect 20772 23264 20778 23316
rect 21637 23307 21695 23313
rect 21637 23273 21649 23307
rect 21683 23304 21695 23307
rect 22278 23304 22284 23316
rect 21683 23276 22284 23304
rect 21683 23273 21695 23276
rect 21637 23267 21695 23273
rect 22278 23264 22284 23276
rect 22336 23264 22342 23316
rect 23198 23304 23204 23316
rect 23159 23276 23204 23304
rect 23198 23264 23204 23276
rect 23256 23264 23262 23316
rect 20254 23236 20260 23248
rect 17920 23208 19012 23236
rect 19076 23208 20260 23236
rect 17920 23196 17926 23208
rect 15933 23171 15991 23177
rect 15933 23168 15945 23171
rect 15896 23140 15945 23168
rect 15896 23128 15902 23140
rect 15933 23137 15945 23140
rect 15979 23137 15991 23171
rect 15933 23131 15991 23137
rect 16117 23171 16175 23177
rect 16117 23137 16129 23171
rect 16163 23137 16175 23171
rect 17328 23168 17356 23196
rect 18782 23168 18788 23180
rect 17328 23140 18788 23168
rect 16117 23131 16175 23137
rect 18782 23128 18788 23140
rect 18840 23168 18846 23180
rect 19076 23168 19104 23208
rect 20254 23196 20260 23208
rect 20312 23196 20318 23248
rect 21726 23196 21732 23248
rect 21784 23236 21790 23248
rect 22189 23239 22247 23245
rect 22189 23236 22201 23239
rect 21784 23208 22201 23236
rect 21784 23196 21790 23208
rect 22189 23205 22201 23208
rect 22235 23205 22247 23239
rect 22189 23199 22247 23205
rect 22370 23196 22376 23248
rect 22428 23236 22434 23248
rect 23017 23239 23075 23245
rect 23017 23236 23029 23239
rect 22428 23208 23029 23236
rect 22428 23196 22434 23208
rect 23017 23205 23029 23208
rect 23063 23236 23075 23239
rect 23661 23239 23719 23245
rect 23661 23236 23673 23239
rect 23063 23208 23673 23236
rect 23063 23205 23075 23208
rect 23017 23199 23075 23205
rect 23661 23205 23673 23208
rect 23707 23205 23719 23239
rect 23661 23199 23719 23205
rect 22738 23168 22744 23180
rect 18840 23140 19104 23168
rect 19444 23140 21588 23168
rect 22699 23140 22744 23168
rect 18840 23128 18846 23140
rect 16022 23100 16028 23112
rect 15983 23072 16028 23100
rect 16022 23060 16028 23072
rect 16080 23060 16086 23112
rect 16206 23060 16212 23112
rect 16264 23100 16270 23112
rect 16942 23100 16948 23112
rect 16264 23072 16309 23100
rect 16903 23072 16948 23100
rect 16264 23060 16270 23072
rect 16942 23060 16948 23072
rect 17000 23060 17006 23112
rect 18046 23100 18052 23112
rect 17956 23072 18052 23100
rect 14921 23035 14979 23041
rect 14921 23001 14933 23035
rect 14967 23032 14979 23035
rect 16574 23032 16580 23044
rect 14967 23004 16580 23032
rect 14967 23001 14979 23004
rect 14921 22995 14979 23001
rect 16574 22992 16580 23004
rect 16632 22992 16638 23044
rect 16850 22992 16856 23044
rect 16908 23032 16914 23044
rect 17956 23041 17984 23072
rect 18046 23060 18052 23072
rect 18104 23060 18110 23112
rect 19058 23060 19064 23112
rect 19116 23100 19122 23112
rect 19245 23103 19303 23109
rect 19245 23100 19257 23103
rect 19116 23072 19257 23100
rect 19116 23060 19122 23072
rect 19245 23069 19257 23072
rect 19291 23069 19303 23103
rect 19444 23094 19472 23140
rect 20530 23100 20536 23112
rect 19245 23063 19303 23069
rect 19352 23066 19472 23094
rect 20491 23072 20536 23100
rect 17037 23035 17095 23041
rect 17037 23032 17049 23035
rect 16908 23004 17049 23032
rect 16908 22992 16914 23004
rect 17037 23001 17049 23004
rect 17083 23001 17095 23035
rect 17037 22995 17095 23001
rect 17941 23035 17999 23041
rect 17941 23001 17953 23035
rect 17987 23001 17999 23035
rect 18138 23032 18144 23044
rect 18099 23004 18144 23032
rect 17941 22995 17999 23001
rect 18138 22992 18144 23004
rect 18196 22992 18202 23044
rect 18966 22992 18972 23044
rect 19024 23032 19030 23044
rect 19352 23032 19380 23066
rect 20530 23060 20536 23072
rect 20588 23060 20594 23112
rect 20711 23103 20769 23109
rect 20711 23069 20723 23103
rect 20757 23100 20769 23103
rect 20990 23100 20996 23112
rect 20757 23072 20996 23100
rect 20757 23069 20769 23072
rect 20711 23063 20769 23069
rect 20990 23060 20996 23072
rect 21048 23060 21054 23112
rect 21560 23109 21588 23140
rect 22738 23128 22744 23140
rect 22796 23128 22802 23180
rect 21545 23103 21603 23109
rect 21545 23069 21557 23103
rect 21591 23069 21603 23103
rect 21545 23063 21603 23069
rect 21726 23060 21732 23112
rect 21784 23100 21790 23112
rect 24397 23103 24455 23109
rect 24397 23100 24409 23103
rect 21784 23072 24409 23100
rect 21784 23060 21790 23072
rect 24397 23069 24409 23072
rect 24443 23100 24455 23103
rect 24578 23100 24584 23112
rect 24443 23072 24584 23100
rect 24443 23069 24455 23072
rect 24397 23063 24455 23069
rect 24578 23060 24584 23072
rect 24636 23060 24642 23112
rect 19024 23004 19380 23032
rect 19024 22992 19030 23004
rect 13998 22924 14004 22976
rect 14056 22964 14062 22976
rect 15102 22964 15108 22976
rect 15160 22973 15166 22976
rect 15160 22967 15179 22973
rect 14056 22936 15108 22964
rect 14056 22924 14062 22936
rect 15102 22924 15108 22936
rect 15167 22933 15179 22967
rect 15160 22927 15179 22933
rect 15160 22924 15166 22927
rect 16666 22924 16672 22976
rect 16724 22964 16730 22976
rect 17129 22967 17187 22973
rect 17129 22964 17141 22967
rect 16724 22936 17141 22964
rect 16724 22924 16730 22936
rect 17129 22933 17141 22936
rect 17175 22964 17187 22967
rect 17770 22964 17776 22976
rect 17175 22936 17776 22964
rect 17175 22933 17187 22936
rect 17129 22927 17187 22933
rect 17770 22924 17776 22936
rect 17828 22924 17834 22976
rect 18693 22967 18751 22973
rect 18693 22933 18705 22967
rect 18739 22964 18751 22967
rect 18782 22964 18788 22976
rect 18739 22936 18788 22964
rect 18739 22933 18751 22936
rect 18693 22927 18751 22933
rect 18782 22924 18788 22936
rect 18840 22924 18846 22976
rect 19518 22924 19524 22976
rect 19576 22964 19582 22976
rect 19705 22967 19763 22973
rect 19705 22964 19717 22967
rect 19576 22936 19717 22964
rect 19576 22924 19582 22936
rect 19705 22933 19717 22936
rect 19751 22933 19763 22967
rect 19705 22927 19763 22933
rect 1104 22874 38824 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 38824 22874
rect 1104 22800 38824 22822
rect 14826 22760 14832 22772
rect 14787 22732 14832 22760
rect 14826 22720 14832 22732
rect 14884 22720 14890 22772
rect 15102 22720 15108 22772
rect 15160 22760 15166 22772
rect 15473 22763 15531 22769
rect 15473 22760 15485 22763
rect 15160 22732 15485 22760
rect 15160 22720 15166 22732
rect 15473 22729 15485 22732
rect 15519 22729 15531 22763
rect 15473 22723 15531 22729
rect 15749 22763 15807 22769
rect 15749 22729 15761 22763
rect 15795 22760 15807 22763
rect 16206 22760 16212 22772
rect 15795 22732 16212 22760
rect 15795 22729 15807 22732
rect 15749 22723 15807 22729
rect 16206 22720 16212 22732
rect 16264 22720 16270 22772
rect 17126 22760 17132 22772
rect 17087 22732 17132 22760
rect 17126 22720 17132 22732
rect 17184 22720 17190 22772
rect 17402 22760 17408 22772
rect 17363 22732 17408 22760
rect 17402 22720 17408 22732
rect 17460 22720 17466 22772
rect 17865 22763 17923 22769
rect 17865 22729 17877 22763
rect 17911 22760 17923 22763
rect 18046 22760 18052 22772
rect 17911 22732 18052 22760
rect 17911 22729 17923 22732
rect 17865 22723 17923 22729
rect 18046 22720 18052 22732
rect 18104 22720 18110 22772
rect 20530 22760 20536 22772
rect 18248 22732 20536 22760
rect 16850 22692 16856 22704
rect 15028 22664 16856 22692
rect 15028 22636 15056 22664
rect 16850 22652 16856 22664
rect 16908 22652 16914 22704
rect 16942 22652 16948 22704
rect 17000 22692 17006 22704
rect 17000 22664 18000 22692
rect 17000 22652 17006 22664
rect 14642 22584 14648 22636
rect 14700 22624 14706 22636
rect 14829 22627 14887 22633
rect 14829 22624 14841 22627
rect 14700 22596 14841 22624
rect 14700 22584 14706 22596
rect 14829 22593 14841 22596
rect 14875 22593 14887 22627
rect 15010 22624 15016 22636
rect 14971 22596 15016 22624
rect 14829 22587 14887 22593
rect 15010 22584 15016 22596
rect 15068 22584 15074 22636
rect 15378 22584 15384 22636
rect 15436 22624 15442 22636
rect 15473 22627 15531 22633
rect 15473 22624 15485 22627
rect 15436 22596 15485 22624
rect 15436 22584 15442 22596
rect 15473 22593 15485 22596
rect 15519 22593 15531 22627
rect 15473 22587 15531 22593
rect 15637 22627 15695 22633
rect 15637 22593 15649 22627
rect 15683 22624 15695 22627
rect 15838 22624 15844 22636
rect 15683 22593 15700 22624
rect 15799 22596 15844 22624
rect 15637 22587 15700 22593
rect 15672 22556 15700 22587
rect 15838 22584 15844 22596
rect 15896 22584 15902 22636
rect 17052 22633 17080 22664
rect 17972 22636 18000 22664
rect 18248 22636 18276 22732
rect 20530 22720 20536 22732
rect 20588 22720 20594 22772
rect 20714 22720 20720 22772
rect 20772 22760 20778 22772
rect 22005 22763 22063 22769
rect 22005 22760 22017 22763
rect 20772 22732 22017 22760
rect 20772 22720 20778 22732
rect 22005 22729 22017 22732
rect 22051 22729 22063 22763
rect 22005 22723 22063 22729
rect 22738 22720 22744 22772
rect 22796 22760 22802 22772
rect 23845 22763 23903 22769
rect 23845 22760 23857 22763
rect 22796 22732 23857 22760
rect 22796 22720 22802 22732
rect 23845 22729 23857 22732
rect 23891 22729 23903 22763
rect 23845 22723 23903 22729
rect 18966 22692 18972 22704
rect 18340 22664 18972 22692
rect 17037 22627 17095 22633
rect 17037 22593 17049 22627
rect 17083 22593 17095 22627
rect 17251 22627 17309 22633
rect 17251 22624 17263 22627
rect 17037 22587 17095 22593
rect 17144 22596 17263 22624
rect 16022 22556 16028 22568
rect 15672 22528 16028 22556
rect 16022 22516 16028 22528
rect 16080 22556 16086 22568
rect 17144 22556 17172 22596
rect 17251 22593 17263 22596
rect 17297 22624 17309 22627
rect 17297 22596 17816 22624
rect 17297 22593 17309 22596
rect 17251 22587 17309 22593
rect 16080 22528 17172 22556
rect 17405 22559 17463 22565
rect 16080 22516 16086 22528
rect 17405 22525 17417 22559
rect 17451 22525 17463 22559
rect 17405 22519 17463 22525
rect 15378 22380 15384 22432
rect 15436 22420 15442 22432
rect 17420 22420 17448 22519
rect 17788 22488 17816 22596
rect 17954 22584 17960 22636
rect 18012 22624 18018 22636
rect 18049 22627 18107 22633
rect 18049 22624 18061 22627
rect 18012 22596 18061 22624
rect 18012 22584 18018 22596
rect 18049 22593 18061 22596
rect 18095 22593 18107 22627
rect 18230 22624 18236 22636
rect 18191 22596 18236 22624
rect 18049 22587 18107 22593
rect 18230 22584 18236 22596
rect 18288 22584 18294 22636
rect 18340 22633 18368 22664
rect 18966 22652 18972 22664
rect 19024 22652 19030 22704
rect 19058 22652 19064 22704
rect 19116 22692 19122 22704
rect 21174 22692 21180 22704
rect 19116 22664 20300 22692
rect 19116 22652 19122 22664
rect 18325 22627 18383 22633
rect 18325 22593 18337 22627
rect 18371 22593 18383 22627
rect 18325 22587 18383 22593
rect 17862 22516 17868 22568
rect 17920 22556 17926 22568
rect 18141 22559 18199 22565
rect 18141 22556 18153 22559
rect 17920 22528 18153 22556
rect 17920 22516 17926 22528
rect 18141 22525 18153 22528
rect 18187 22525 18199 22559
rect 18141 22519 18199 22525
rect 18340 22488 18368 22587
rect 18782 22584 18788 22636
rect 18840 22624 18846 22636
rect 20272 22633 20300 22664
rect 21100 22664 21180 22692
rect 21100 22633 21128 22664
rect 21174 22652 21180 22664
rect 21232 22692 21238 22704
rect 21232 22664 22048 22692
rect 21232 22652 21238 22664
rect 22020 22636 22048 22664
rect 19981 22627 20039 22633
rect 19981 22624 19993 22627
rect 18840 22596 19993 22624
rect 18840 22584 18846 22596
rect 19981 22593 19993 22596
rect 20027 22624 20039 22627
rect 20257 22627 20315 22633
rect 20027 22596 20208 22624
rect 20027 22593 20039 22596
rect 19981 22587 20039 22593
rect 18874 22556 18880 22568
rect 18835 22528 18880 22556
rect 18874 22516 18880 22528
rect 18932 22516 18938 22568
rect 17788 22460 18368 22488
rect 19058 22448 19064 22500
rect 19116 22488 19122 22500
rect 19245 22491 19303 22497
rect 19245 22488 19257 22491
rect 19116 22460 19257 22488
rect 19116 22448 19122 22460
rect 19245 22457 19257 22460
rect 19291 22457 19303 22491
rect 19245 22451 19303 22457
rect 19337 22491 19395 22497
rect 19337 22457 19349 22491
rect 19383 22488 19395 22491
rect 20070 22488 20076 22500
rect 19383 22460 20076 22488
rect 19383 22457 19395 22460
rect 19337 22451 19395 22457
rect 20070 22448 20076 22460
rect 20128 22448 20134 22500
rect 20180 22488 20208 22596
rect 20257 22593 20269 22627
rect 20303 22593 20315 22627
rect 20257 22587 20315 22593
rect 21085 22627 21143 22633
rect 21085 22593 21097 22627
rect 21131 22593 21143 22627
rect 21266 22624 21272 22636
rect 21227 22596 21272 22624
rect 21085 22587 21143 22593
rect 21266 22584 21272 22596
rect 21324 22584 21330 22636
rect 21726 22584 21732 22636
rect 21784 22624 21790 22636
rect 21821 22627 21879 22633
rect 21821 22624 21833 22627
rect 21784 22596 21833 22624
rect 21784 22584 21790 22596
rect 21821 22593 21833 22596
rect 21867 22593 21879 22627
rect 21821 22587 21879 22593
rect 22002 22584 22008 22636
rect 22060 22584 22066 22636
rect 22097 22627 22155 22633
rect 22097 22593 22109 22627
rect 22143 22593 22155 22627
rect 22097 22587 22155 22593
rect 20806 22516 20812 22568
rect 20864 22556 20870 22568
rect 22112 22556 22140 22587
rect 22186 22584 22192 22636
rect 22244 22624 22250 22636
rect 22281 22627 22339 22633
rect 22281 22624 22293 22627
rect 22244 22596 22293 22624
rect 22244 22584 22250 22596
rect 22281 22593 22293 22596
rect 22327 22593 22339 22627
rect 22281 22587 22339 22593
rect 22741 22559 22799 22565
rect 22741 22556 22753 22559
rect 20864 22528 22753 22556
rect 20864 22516 20870 22528
rect 22741 22525 22753 22528
rect 22787 22525 22799 22559
rect 22741 22519 22799 22525
rect 21726 22488 21732 22500
rect 20180 22460 21732 22488
rect 21726 22448 21732 22460
rect 21784 22448 21790 22500
rect 18230 22420 18236 22432
rect 15436 22392 18236 22420
rect 15436 22380 15442 22392
rect 18230 22380 18236 22392
rect 18288 22380 18294 22432
rect 19797 22423 19855 22429
rect 19797 22389 19809 22423
rect 19843 22420 19855 22423
rect 19978 22420 19984 22432
rect 19843 22392 19984 22420
rect 19843 22389 19855 22392
rect 19797 22383 19855 22389
rect 19978 22380 19984 22392
rect 20036 22380 20042 22432
rect 20165 22423 20223 22429
rect 20165 22389 20177 22423
rect 20211 22420 20223 22423
rect 20254 22420 20260 22432
rect 20211 22392 20260 22420
rect 20211 22389 20223 22392
rect 20165 22383 20223 22389
rect 20254 22380 20260 22392
rect 20312 22380 20318 22432
rect 20898 22380 20904 22432
rect 20956 22420 20962 22432
rect 21177 22423 21235 22429
rect 21177 22420 21189 22423
rect 20956 22392 21189 22420
rect 20956 22380 20962 22392
rect 21177 22389 21189 22392
rect 21223 22389 21235 22423
rect 23290 22420 23296 22432
rect 23251 22392 23296 22420
rect 21177 22383 21235 22389
rect 23290 22380 23296 22392
rect 23348 22380 23354 22432
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 16666 22216 16672 22228
rect 16627 22188 16672 22216
rect 16666 22176 16672 22188
rect 16724 22176 16730 22228
rect 17865 22219 17923 22225
rect 17865 22185 17877 22219
rect 17911 22216 17923 22219
rect 18138 22216 18144 22228
rect 17911 22188 18144 22216
rect 17911 22185 17923 22188
rect 17865 22179 17923 22185
rect 18138 22176 18144 22188
rect 18196 22176 18202 22228
rect 18230 22176 18236 22228
rect 18288 22216 18294 22228
rect 18966 22216 18972 22228
rect 18288 22188 18972 22216
rect 18288 22176 18294 22188
rect 18966 22176 18972 22188
rect 19024 22176 19030 22228
rect 19058 22176 19064 22228
rect 19116 22216 19122 22228
rect 20346 22216 20352 22228
rect 19116 22188 20352 22216
rect 19116 22176 19122 22188
rect 20346 22176 20352 22188
rect 20404 22176 20410 22228
rect 17957 22151 18015 22157
rect 17957 22117 17969 22151
rect 18003 22148 18015 22151
rect 20806 22148 20812 22160
rect 18003 22120 20812 22148
rect 18003 22117 18015 22120
rect 17957 22111 18015 22117
rect 20806 22108 20812 22120
rect 20864 22108 20870 22160
rect 22646 22108 22652 22160
rect 22704 22148 22710 22160
rect 23290 22148 23296 22160
rect 22704 22120 23296 22148
rect 22704 22108 22710 22120
rect 23290 22108 23296 22120
rect 23348 22108 23354 22160
rect 22741 22083 22799 22089
rect 22741 22080 22753 22083
rect 18064 22052 22753 22080
rect 18064 22021 18092 22052
rect 22741 22049 22753 22052
rect 22787 22049 22799 22083
rect 22741 22043 22799 22049
rect 17497 22015 17555 22021
rect 17497 21981 17509 22015
rect 17543 21981 17555 22015
rect 17497 21975 17555 21981
rect 18049 22015 18107 22021
rect 18049 21981 18061 22015
rect 18095 21981 18107 22015
rect 18049 21975 18107 21981
rect 18693 22015 18751 22021
rect 18693 21981 18705 22015
rect 18739 22012 18751 22015
rect 19242 22012 19248 22024
rect 18739 21984 19248 22012
rect 18739 21981 18751 21984
rect 18693 21975 18751 21981
rect 17512 21944 17540 21975
rect 19242 21972 19248 21984
rect 19300 21972 19306 22024
rect 19886 22012 19892 22024
rect 19720 21984 19892 22012
rect 19720 21944 19748 21984
rect 19886 21972 19892 21984
rect 19944 21972 19950 22024
rect 20530 22012 20536 22024
rect 20491 21984 20536 22012
rect 20530 21972 20536 21984
rect 20588 21972 20594 22024
rect 20898 22012 20904 22024
rect 20859 21984 20904 22012
rect 20898 21972 20904 21984
rect 20956 21972 20962 22024
rect 21542 21972 21548 22024
rect 21600 22012 21606 22024
rect 21637 22015 21695 22021
rect 21637 22012 21649 22015
rect 21600 21984 21649 22012
rect 21600 21972 21606 21984
rect 21637 21981 21649 21984
rect 21683 21981 21695 22015
rect 21867 22015 21925 22021
rect 21867 22012 21879 22015
rect 21637 21975 21695 21981
rect 21744 21984 21879 22012
rect 17512 21916 19748 21944
rect 19797 21947 19855 21953
rect 19797 21913 19809 21947
rect 19843 21944 19855 21947
rect 20162 21944 20168 21956
rect 19843 21916 20168 21944
rect 19843 21913 19855 21916
rect 19797 21907 19855 21913
rect 20162 21904 20168 21916
rect 20220 21904 20226 21956
rect 21266 21904 21272 21956
rect 21324 21944 21330 21956
rect 21744 21944 21772 21984
rect 21867 21981 21879 21984
rect 21913 21981 21925 22015
rect 21867 21975 21925 21981
rect 22002 21972 22008 22024
rect 22060 22012 22066 22024
rect 22646 22012 22652 22024
rect 22060 21984 22105 22012
rect 22607 21984 22652 22012
rect 22060 21972 22066 21984
rect 22646 21972 22652 21984
rect 22704 21972 22710 22024
rect 22833 22015 22891 22021
rect 22833 21981 22845 22015
rect 22879 22012 22891 22015
rect 23106 22012 23112 22024
rect 22879 21984 23112 22012
rect 22879 21981 22891 21984
rect 22833 21975 22891 21981
rect 23106 21972 23112 21984
rect 23164 21972 23170 22024
rect 23308 22021 23336 22108
rect 23293 22015 23351 22021
rect 23293 21981 23305 22015
rect 23339 21981 23351 22015
rect 23293 21975 23351 21981
rect 21324 21916 21772 21944
rect 22020 21944 22048 21972
rect 23385 21947 23443 21953
rect 23385 21944 23397 21947
rect 22020 21916 23397 21944
rect 21324 21904 21330 21916
rect 23385 21913 23397 21916
rect 23431 21913 23443 21947
rect 23385 21907 23443 21913
rect 17589 21879 17647 21885
rect 17589 21845 17601 21879
rect 17635 21876 17647 21879
rect 18322 21876 18328 21888
rect 17635 21848 18328 21876
rect 17635 21845 17647 21848
rect 17589 21839 17647 21845
rect 18322 21836 18328 21848
rect 18380 21876 18386 21888
rect 21729 21879 21787 21885
rect 21729 21876 21741 21879
rect 18380 21848 21741 21876
rect 18380 21836 18386 21848
rect 21729 21845 21741 21848
rect 21775 21845 21787 21879
rect 21729 21839 21787 21845
rect 1104 21786 38824 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 38824 21786
rect 1104 21712 38824 21734
rect 18230 21672 18236 21684
rect 18191 21644 18236 21672
rect 18230 21632 18236 21644
rect 18288 21632 18294 21684
rect 18785 21675 18843 21681
rect 18785 21641 18797 21675
rect 18831 21672 18843 21675
rect 18874 21672 18880 21684
rect 18831 21644 18880 21672
rect 18831 21641 18843 21644
rect 18785 21635 18843 21641
rect 18874 21632 18880 21644
rect 18932 21632 18938 21684
rect 19797 21675 19855 21681
rect 19797 21641 19809 21675
rect 19843 21672 19855 21675
rect 19978 21672 19984 21684
rect 19843 21644 19984 21672
rect 19843 21641 19855 21644
rect 19797 21635 19855 21641
rect 19978 21632 19984 21644
rect 20036 21632 20042 21684
rect 20717 21675 20775 21681
rect 20717 21641 20729 21675
rect 20763 21672 20775 21675
rect 20806 21672 20812 21684
rect 20763 21644 20812 21672
rect 20763 21641 20775 21644
rect 20717 21635 20775 21641
rect 20806 21632 20812 21644
rect 20864 21632 20870 21684
rect 23290 21632 23296 21684
rect 23348 21672 23354 21684
rect 23753 21675 23811 21681
rect 23753 21672 23765 21675
rect 23348 21644 23765 21672
rect 23348 21632 23354 21644
rect 23753 21641 23765 21644
rect 23799 21641 23811 21675
rect 23753 21635 23811 21641
rect 20530 21564 20536 21616
rect 20588 21604 20594 21616
rect 20588 21576 20944 21604
rect 20588 21564 20594 21576
rect 19426 21496 19432 21548
rect 19484 21536 19490 21548
rect 19705 21539 19763 21545
rect 19705 21536 19717 21539
rect 19484 21508 19717 21536
rect 19484 21496 19490 21508
rect 19705 21505 19717 21508
rect 19751 21505 19763 21539
rect 20070 21536 20076 21548
rect 20031 21508 20076 21536
rect 19705 21499 19763 21505
rect 20070 21496 20076 21508
rect 20128 21496 20134 21548
rect 20257 21539 20315 21545
rect 20257 21505 20269 21539
rect 20303 21536 20315 21539
rect 20714 21536 20720 21548
rect 20303 21508 20720 21536
rect 20303 21505 20315 21508
rect 20257 21499 20315 21505
rect 20714 21496 20720 21508
rect 20772 21496 20778 21548
rect 20916 21545 20944 21576
rect 20901 21539 20959 21545
rect 20901 21505 20913 21539
rect 20947 21505 20959 21539
rect 21082 21536 21088 21548
rect 21043 21508 21088 21536
rect 20901 21499 20959 21505
rect 21082 21496 21088 21508
rect 21140 21496 21146 21548
rect 21174 21496 21180 21548
rect 21232 21536 21238 21548
rect 21232 21508 21277 21536
rect 21232 21496 21238 21508
rect 21542 21496 21548 21548
rect 21600 21536 21606 21548
rect 22097 21539 22155 21545
rect 22097 21536 22109 21539
rect 21600 21508 22109 21536
rect 21600 21496 21606 21508
rect 22097 21505 22109 21508
rect 22143 21505 22155 21539
rect 22097 21499 22155 21505
rect 22278 21496 22284 21548
rect 22336 21536 22342 21548
rect 22646 21536 22652 21548
rect 22336 21508 22652 21536
rect 22336 21496 22342 21508
rect 22646 21496 22652 21508
rect 22704 21496 22710 21548
rect 22925 21539 22983 21545
rect 22925 21505 22937 21539
rect 22971 21536 22983 21539
rect 23106 21536 23112 21548
rect 22971 21508 23112 21536
rect 22971 21505 22983 21508
rect 22925 21499 22983 21505
rect 23106 21496 23112 21508
rect 23164 21496 23170 21548
rect 20438 21428 20444 21480
rect 20496 21468 20502 21480
rect 21821 21471 21879 21477
rect 21821 21468 21833 21471
rect 20496 21440 21833 21468
rect 20496 21428 20502 21440
rect 21821 21437 21833 21440
rect 21867 21437 21879 21471
rect 21821 21431 21879 21437
rect 22186 21428 22192 21480
rect 22244 21468 22250 21480
rect 22373 21471 22431 21477
rect 22373 21468 22385 21471
rect 22244 21440 22385 21468
rect 22244 21428 22250 21440
rect 22373 21437 22385 21440
rect 22419 21437 22431 21471
rect 22373 21431 22431 21437
rect 20073 21403 20131 21409
rect 20073 21369 20085 21403
rect 20119 21400 20131 21403
rect 21082 21400 21088 21412
rect 20119 21372 21088 21400
rect 20119 21369 20131 21372
rect 20073 21363 20131 21369
rect 21082 21360 21088 21372
rect 21140 21360 21146 21412
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 21542 21128 21548 21140
rect 21503 21100 21548 21128
rect 21542 21088 21548 21100
rect 21600 21088 21606 21140
rect 22186 21128 22192 21140
rect 22147 21100 22192 21128
rect 22186 21088 22192 21100
rect 22244 21088 22250 21140
rect 18690 21020 18696 21072
rect 18748 21060 18754 21072
rect 19429 21063 19487 21069
rect 19429 21060 19441 21063
rect 18748 21032 19441 21060
rect 18748 21020 18754 21032
rect 19429 21029 19441 21032
rect 19475 21029 19487 21063
rect 20533 21063 20591 21069
rect 20533 21060 20545 21063
rect 19429 21023 19487 21029
rect 19582 21032 20545 21060
rect 19058 20952 19064 21004
rect 19116 20992 19122 21004
rect 19582 21001 19610 21032
rect 20533 21029 20545 21032
rect 20579 21060 20591 21063
rect 21174 21060 21180 21072
rect 20579 21032 21180 21060
rect 20579 21029 20591 21032
rect 20533 21023 20591 21029
rect 21174 21020 21180 21032
rect 21232 21020 21238 21072
rect 19567 20995 19625 21001
rect 19567 20992 19579 20995
rect 19116 20964 19579 20992
rect 19116 20952 19122 20964
rect 19567 20961 19579 20964
rect 19613 20961 19625 20995
rect 21082 20992 21088 21004
rect 19567 20955 19625 20961
rect 19720 20964 21088 20992
rect 18693 20927 18751 20933
rect 18693 20893 18705 20927
rect 18739 20924 18751 20927
rect 19334 20924 19340 20936
rect 18739 20896 19340 20924
rect 18739 20893 18751 20896
rect 18693 20887 18751 20893
rect 19334 20884 19340 20896
rect 19392 20884 19398 20936
rect 19720 20933 19748 20964
rect 21082 20952 21088 20964
rect 21140 20992 21146 21004
rect 21140 20964 22140 20992
rect 21140 20952 21146 20964
rect 19705 20927 19763 20933
rect 19705 20893 19717 20927
rect 19751 20893 19763 20927
rect 19705 20887 19763 20893
rect 20530 20884 20536 20936
rect 20588 20924 20594 20936
rect 22112 20933 22140 20964
rect 21453 20927 21511 20933
rect 21453 20924 21465 20927
rect 20588 20896 21465 20924
rect 20588 20884 20594 20896
rect 21453 20893 21465 20896
rect 21499 20893 21511 20927
rect 21453 20887 21511 20893
rect 22097 20927 22155 20933
rect 22097 20893 22109 20927
rect 22143 20893 22155 20927
rect 22278 20924 22284 20936
rect 22239 20896 22284 20924
rect 22097 20887 22155 20893
rect 19352 20856 19380 20884
rect 20548 20856 20576 20884
rect 19352 20828 20576 20856
rect 21468 20856 21496 20887
rect 22278 20884 22284 20896
rect 22336 20884 22342 20936
rect 22741 20859 22799 20865
rect 22741 20856 22753 20859
rect 21468 20828 22753 20856
rect 22741 20825 22753 20828
rect 22787 20825 22799 20859
rect 22741 20819 22799 20825
rect 1104 20698 38824 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 38824 20698
rect 1104 20624 38824 20646
rect 19058 20544 19064 20596
rect 19116 20584 19122 20596
rect 19153 20587 19211 20593
rect 19153 20584 19165 20587
rect 19116 20556 19165 20584
rect 19116 20544 19122 20556
rect 19153 20553 19165 20556
rect 19199 20553 19211 20587
rect 19153 20547 19211 20553
rect 20441 20587 20499 20593
rect 20441 20553 20453 20587
rect 20487 20584 20499 20587
rect 20530 20584 20536 20596
rect 20487 20556 20536 20584
rect 20487 20553 20499 20556
rect 20441 20547 20499 20553
rect 20530 20544 20536 20556
rect 20588 20544 20594 20596
rect 21174 20544 21180 20596
rect 21232 20584 21238 20596
rect 21821 20587 21879 20593
rect 21821 20584 21833 20587
rect 21232 20556 21833 20584
rect 21232 20544 21238 20556
rect 21821 20553 21833 20556
rect 21867 20584 21879 20587
rect 22278 20584 22284 20596
rect 21867 20556 22284 20584
rect 21867 20553 21879 20556
rect 21821 20547 21879 20553
rect 22278 20544 22284 20556
rect 22336 20584 22342 20596
rect 22373 20587 22431 20593
rect 22373 20584 22385 20587
rect 22336 20556 22385 20584
rect 22336 20544 22342 20556
rect 22373 20553 22385 20556
rect 22419 20553 22431 20587
rect 22373 20547 22431 20553
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 1104 19610 38824 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 38824 19610
rect 1104 19536 38824 19558
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 1104 18522 38824 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 38824 18522
rect 1104 18448 38824 18470
rect 1581 18411 1639 18417
rect 1581 18377 1593 18411
rect 1627 18408 1639 18411
rect 9398 18408 9404 18420
rect 1627 18380 9404 18408
rect 1627 18377 1639 18380
rect 1581 18371 1639 18377
rect 9398 18368 9404 18380
rect 9456 18368 9462 18420
rect 1394 18272 1400 18284
rect 1355 18244 1400 18272
rect 1394 18232 1400 18244
rect 1452 18272 1458 18284
rect 2041 18275 2099 18281
rect 2041 18272 2053 18275
rect 1452 18244 2053 18272
rect 1452 18232 1458 18244
rect 2041 18241 2053 18244
rect 2087 18241 2099 18275
rect 2041 18235 2099 18241
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 1104 17434 38824 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 38824 17434
rect 1104 17360 38824 17382
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 1104 16346 38824 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 38824 16346
rect 1104 16272 38824 16294
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 1104 15258 38824 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 38824 15258
rect 1104 15184 38824 15206
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 1104 14170 38824 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 38824 14170
rect 1104 14096 38824 14118
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 1104 13082 38824 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 38824 13082
rect 1104 13008 38824 13030
rect 18506 12792 18512 12844
rect 18564 12832 18570 12844
rect 37277 12835 37335 12841
rect 37277 12832 37289 12835
rect 18564 12804 37289 12832
rect 18564 12792 18570 12804
rect 37277 12801 37289 12804
rect 37323 12832 37335 12835
rect 37829 12835 37887 12841
rect 37829 12832 37841 12835
rect 37323 12804 37841 12832
rect 37323 12801 37335 12804
rect 37277 12795 37335 12801
rect 37829 12801 37841 12804
rect 37875 12801 37887 12835
rect 37829 12795 37887 12801
rect 37918 12588 37924 12640
rect 37976 12628 37982 12640
rect 38013 12631 38071 12637
rect 38013 12628 38025 12631
rect 37976 12600 38025 12628
rect 37976 12588 37982 12600
rect 38013 12597 38025 12600
rect 38059 12597 38071 12631
rect 38013 12591 38071 12597
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 38102 12356 38108 12368
rect 38063 12328 38108 12356
rect 38102 12316 38108 12328
rect 38160 12316 38166 12368
rect 37918 12220 37924 12232
rect 37879 12192 37924 12220
rect 37918 12180 37924 12192
rect 37976 12180 37982 12232
rect 1104 11994 38824 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 38824 11994
rect 1104 11920 38824 11942
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 1104 10906 38824 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 38824 10906
rect 1104 10832 38824 10854
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 1104 9818 38824 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 38824 9818
rect 1104 9744 38824 9766
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 1104 8730 38824 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 38824 8730
rect 1104 8656 38824 8678
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 1104 7642 38824 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 38824 7642
rect 1104 7568 38824 7590
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 1104 6554 38824 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 38824 6554
rect 1104 6480 38824 6502
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 1104 5466 38824 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 38824 5466
rect 1104 5392 38824 5414
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 1104 4378 38824 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 38824 4378
rect 1104 4304 38824 4326
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 1104 3290 38824 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 38824 3290
rect 1104 3216 38824 3238
rect 14 2796 20 2848
rect 72 2836 78 2848
rect 1394 2836 1400 2848
rect 72 2808 1400 2836
rect 72 2796 78 2808
rect 1394 2796 1400 2808
rect 1452 2796 1458 2848
rect 34514 2796 34520 2848
rect 34572 2836 34578 2848
rect 34885 2839 34943 2845
rect 34885 2836 34897 2839
rect 34572 2808 34897 2836
rect 34572 2796 34578 2808
rect 34885 2805 34897 2808
rect 34931 2805 34943 2839
rect 34885 2799 34943 2805
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 15746 2592 15752 2644
rect 15804 2632 15810 2644
rect 16853 2635 16911 2641
rect 16853 2632 16865 2635
rect 15804 2604 16865 2632
rect 15804 2592 15810 2604
rect 16853 2601 16865 2604
rect 16899 2601 16911 2635
rect 16853 2595 16911 2601
rect 1394 2496 1400 2508
rect 1355 2468 1400 2496
rect 1394 2456 1400 2468
rect 1452 2456 1458 2508
rect 1670 2496 1676 2508
rect 1631 2468 1676 2496
rect 1670 2456 1676 2468
rect 1728 2456 1734 2508
rect 11330 2456 11336 2508
rect 11388 2496 11394 2508
rect 35069 2499 35127 2505
rect 35069 2496 35081 2499
rect 11388 2468 35081 2496
rect 11388 2456 11394 2468
rect 35069 2465 35081 2468
rect 35115 2465 35127 2499
rect 35069 2459 35127 2465
rect 16758 2388 16764 2440
rect 16816 2428 16822 2440
rect 17037 2431 17095 2437
rect 17037 2428 17049 2431
rect 16816 2400 17049 2428
rect 16816 2388 16822 2400
rect 17037 2397 17049 2400
rect 17083 2428 17095 2431
rect 17497 2431 17555 2437
rect 17497 2428 17509 2431
rect 17083 2400 17509 2428
rect 17083 2397 17095 2400
rect 17037 2391 17095 2397
rect 17497 2397 17509 2400
rect 17543 2397 17555 2431
rect 17497 2391 17555 2397
rect 34514 2320 34520 2372
rect 34572 2360 34578 2372
rect 35253 2363 35311 2369
rect 35253 2360 35265 2363
rect 34572 2332 35265 2360
rect 34572 2320 34578 2332
rect 35253 2329 35265 2332
rect 35299 2329 35311 2363
rect 35253 2323 35311 2329
rect 1104 2202 38824 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 30932 37408 30984 37460
rect 17776 37272 17828 37324
rect 13544 37204 13596 37256
rect 14280 37204 14332 37256
rect 30932 37204 30984 37256
rect 31024 37111 31076 37120
rect 31024 37077 31033 37111
rect 31033 37077 31067 37111
rect 31067 37077 31076 37111
rect 31024 37068 31076 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 14280 36907 14332 36916
rect 14280 36873 14289 36907
rect 14289 36873 14323 36907
rect 14323 36873 14332 36907
rect 14280 36864 14332 36873
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 3424 35980 3476 36032
rect 9404 35980 9456 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 8300 35708 8352 35760
rect 6644 35683 6696 35692
rect 6644 35649 6678 35683
rect 6678 35649 6696 35683
rect 6644 35640 6696 35649
rect 17224 35640 17276 35692
rect 18788 35504 18840 35556
rect 17684 35436 17736 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 17132 35028 17184 35080
rect 16764 34960 16816 35012
rect 17132 34892 17184 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 18880 34688 18932 34740
rect 16948 34595 17000 34604
rect 16948 34561 16982 34595
rect 16982 34561 17000 34595
rect 16948 34552 17000 34561
rect 17040 34348 17092 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 17316 34144 17368 34196
rect 17040 33940 17092 33992
rect 16672 33872 16724 33924
rect 15844 33804 15896 33856
rect 31024 33804 31076 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 16672 33643 16724 33652
rect 16672 33609 16681 33643
rect 16681 33609 16715 33643
rect 16715 33609 16724 33643
rect 16672 33600 16724 33609
rect 16488 33464 16540 33516
rect 18144 33464 18196 33516
rect 14188 33396 14240 33448
rect 15844 33396 15896 33448
rect 16028 33396 16080 33448
rect 17960 33396 18012 33448
rect 16672 33328 16724 33380
rect 15108 33260 15160 33312
rect 16028 33303 16080 33312
rect 16028 33269 16037 33303
rect 16037 33269 16071 33303
rect 16071 33269 16080 33303
rect 16028 33260 16080 33269
rect 17316 33260 17368 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 15844 33056 15896 33108
rect 14188 32963 14240 32972
rect 14188 32929 14197 32963
rect 14197 32929 14231 32963
rect 14231 32929 14240 32963
rect 14188 32920 14240 32929
rect 13820 32852 13872 32904
rect 17040 32852 17092 32904
rect 15016 32784 15068 32836
rect 15936 32784 15988 32836
rect 11520 32759 11572 32768
rect 11520 32725 11529 32759
rect 11529 32725 11563 32759
rect 11563 32725 11572 32759
rect 11520 32716 11572 32725
rect 14372 32759 14424 32768
rect 14372 32725 14381 32759
rect 14381 32725 14415 32759
rect 14415 32725 14424 32759
rect 14372 32716 14424 32725
rect 14464 32759 14516 32768
rect 14464 32725 14473 32759
rect 14473 32725 14507 32759
rect 14507 32725 14516 32759
rect 14464 32716 14516 32725
rect 14648 32716 14700 32768
rect 17592 32759 17644 32768
rect 17592 32725 17601 32759
rect 17601 32725 17635 32759
rect 17635 32725 17644 32759
rect 17592 32716 17644 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 14648 32419 14700 32428
rect 14648 32385 14657 32419
rect 14657 32385 14691 32419
rect 14691 32385 14700 32419
rect 14648 32376 14700 32385
rect 16672 32419 16724 32428
rect 16672 32385 16681 32419
rect 16681 32385 16715 32419
rect 16715 32385 16724 32419
rect 16672 32376 16724 32385
rect 15752 32308 15804 32360
rect 18236 32308 18288 32360
rect 14372 32240 14424 32292
rect 14924 32172 14976 32224
rect 16856 32215 16908 32224
rect 16856 32181 16865 32215
rect 16865 32181 16899 32215
rect 16899 32181 16908 32215
rect 16856 32172 16908 32181
rect 17684 32172 17736 32224
rect 21640 32172 21692 32224
rect 37832 32172 37884 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 11520 31968 11572 32020
rect 15016 32011 15068 32020
rect 8300 31696 8352 31748
rect 9680 31764 9732 31816
rect 15016 31977 15025 32011
rect 15025 31977 15059 32011
rect 15059 31977 15068 32011
rect 15016 31968 15068 31977
rect 17224 32011 17276 32020
rect 17224 31977 17233 32011
rect 17233 31977 17267 32011
rect 17267 31977 17276 32011
rect 17224 31968 17276 31977
rect 17316 31968 17368 32020
rect 19432 31968 19484 32020
rect 17960 31900 18012 31952
rect 19524 31900 19576 31952
rect 15108 31764 15160 31816
rect 15568 31832 15620 31884
rect 15752 31807 15804 31816
rect 15752 31773 15761 31807
rect 15761 31773 15795 31807
rect 15795 31773 15804 31807
rect 15752 31764 15804 31773
rect 16304 31696 16356 31748
rect 10968 31671 11020 31680
rect 10968 31637 10977 31671
rect 10977 31637 11011 31671
rect 11011 31637 11020 31671
rect 10968 31628 11020 31637
rect 17224 31832 17276 31884
rect 17684 31832 17736 31884
rect 18144 31832 18196 31884
rect 19432 31764 19484 31816
rect 20260 31807 20312 31816
rect 20260 31773 20269 31807
rect 20269 31773 20303 31807
rect 20303 31773 20312 31807
rect 20260 31764 20312 31773
rect 19340 31696 19392 31748
rect 19524 31739 19576 31748
rect 19524 31705 19533 31739
rect 19533 31705 19567 31739
rect 19567 31705 19576 31739
rect 19524 31696 19576 31705
rect 18512 31628 18564 31680
rect 20628 31628 20680 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 1676 31331 1728 31340
rect 1676 31297 1710 31331
rect 1710 31297 1728 31331
rect 1676 31288 1728 31297
rect 1400 31263 1452 31272
rect 1400 31229 1409 31263
rect 1409 31229 1443 31263
rect 1443 31229 1452 31263
rect 1400 31220 1452 31229
rect 7472 31220 7524 31272
rect 8300 31424 8352 31476
rect 16764 31467 16816 31476
rect 16764 31433 16773 31467
rect 16773 31433 16807 31467
rect 16807 31433 16816 31467
rect 16764 31424 16816 31433
rect 17224 31424 17276 31476
rect 19432 31424 19484 31476
rect 18328 31356 18380 31408
rect 8300 31331 8352 31340
rect 8300 31297 8334 31331
rect 8334 31297 8352 31331
rect 8300 31288 8352 31297
rect 16948 31331 17000 31340
rect 16948 31297 16957 31331
rect 16957 31297 16991 31331
rect 16991 31297 17000 31331
rect 16948 31288 17000 31297
rect 17132 31288 17184 31340
rect 17776 31220 17828 31272
rect 18052 31263 18104 31272
rect 18052 31229 18061 31263
rect 18061 31229 18095 31263
rect 18095 31229 18104 31263
rect 18052 31220 18104 31229
rect 16488 31152 16540 31204
rect 18236 31220 18288 31272
rect 18512 31263 18564 31272
rect 18512 31229 18521 31263
rect 18521 31229 18555 31263
rect 18555 31229 18564 31263
rect 18512 31220 18564 31229
rect 20076 31220 20128 31272
rect 2780 31127 2832 31136
rect 2780 31093 2789 31127
rect 2789 31093 2823 31127
rect 2823 31093 2832 31127
rect 2780 31084 2832 31093
rect 9772 31084 9824 31136
rect 17960 31084 18012 31136
rect 20260 31084 20312 31136
rect 20628 31084 20680 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 16948 30880 17000 30932
rect 13820 30744 13872 30796
rect 37832 30787 37884 30796
rect 9404 30719 9456 30728
rect 9404 30685 9413 30719
rect 9413 30685 9447 30719
rect 9447 30685 9456 30719
rect 9404 30676 9456 30685
rect 37832 30753 37841 30787
rect 37841 30753 37875 30787
rect 37875 30753 37884 30787
rect 37832 30744 37884 30753
rect 16672 30676 16724 30728
rect 17132 30676 17184 30728
rect 17776 30676 17828 30728
rect 20444 30719 20496 30728
rect 20444 30685 20458 30719
rect 20458 30685 20492 30719
rect 20492 30685 20496 30719
rect 38108 30719 38160 30728
rect 20444 30676 20496 30685
rect 38108 30685 38117 30719
rect 38117 30685 38151 30719
rect 38151 30685 38160 30719
rect 38108 30676 38160 30685
rect 11428 30608 11480 30660
rect 18052 30608 18104 30660
rect 18512 30608 18564 30660
rect 20076 30651 20128 30660
rect 20076 30617 20085 30651
rect 20085 30617 20119 30651
rect 20119 30617 20128 30651
rect 20076 30608 20128 30617
rect 20260 30651 20312 30660
rect 20260 30617 20269 30651
rect 20269 30617 20303 30651
rect 20303 30617 20312 30651
rect 20260 30608 20312 30617
rect 10692 30583 10744 30592
rect 10692 30549 10701 30583
rect 10701 30549 10735 30583
rect 10735 30549 10744 30583
rect 10692 30540 10744 30549
rect 15384 30540 15436 30592
rect 18328 30583 18380 30592
rect 18328 30549 18337 30583
rect 18337 30549 18371 30583
rect 18371 30549 18380 30583
rect 18328 30540 18380 30549
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 9404 30336 9456 30388
rect 14464 30336 14516 30388
rect 14924 30336 14976 30388
rect 38108 30379 38160 30388
rect 38108 30345 38117 30379
rect 38117 30345 38151 30379
rect 38151 30345 38160 30379
rect 38108 30336 38160 30345
rect 16580 30268 16632 30320
rect 16672 30243 16724 30252
rect 16672 30209 16681 30243
rect 16681 30209 16715 30243
rect 16715 30209 16724 30243
rect 16672 30200 16724 30209
rect 19340 30268 19392 30320
rect 19432 30268 19484 30320
rect 19616 30268 19668 30320
rect 19984 30268 20036 30320
rect 20444 30268 20496 30320
rect 20076 30200 20128 30252
rect 17960 30132 18012 30184
rect 6644 29996 6696 30048
rect 19616 30064 19668 30116
rect 20260 30132 20312 30184
rect 18972 29996 19024 30048
rect 19800 30039 19852 30048
rect 19800 30005 19809 30039
rect 19809 30005 19843 30039
rect 19843 30005 19852 30039
rect 19800 29996 19852 30005
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 12532 29792 12584 29844
rect 13820 29792 13872 29844
rect 15752 29792 15804 29844
rect 16304 29792 16356 29844
rect 17132 29792 17184 29844
rect 11888 29724 11940 29776
rect 18328 29724 18380 29776
rect 12440 29588 12492 29640
rect 18604 29656 18656 29708
rect 19432 29699 19484 29708
rect 19432 29665 19441 29699
rect 19441 29665 19475 29699
rect 19475 29665 19484 29699
rect 19432 29656 19484 29665
rect 8852 29520 8904 29572
rect 14740 29520 14792 29572
rect 15200 29563 15252 29572
rect 15200 29529 15209 29563
rect 15209 29529 15243 29563
rect 15243 29529 15252 29563
rect 15200 29520 15252 29529
rect 11888 29452 11940 29504
rect 15108 29452 15160 29504
rect 16948 29588 17000 29640
rect 15752 29520 15804 29572
rect 15568 29495 15620 29504
rect 15568 29461 15577 29495
rect 15577 29461 15611 29495
rect 15611 29461 15620 29495
rect 15568 29452 15620 29461
rect 16028 29452 16080 29504
rect 17224 29452 17276 29504
rect 18512 29452 18564 29504
rect 20076 29588 20128 29640
rect 20260 29588 20312 29640
rect 19064 29452 19116 29504
rect 19800 29452 19852 29504
rect 20444 29452 20496 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 8852 29291 8904 29300
rect 8852 29257 8861 29291
rect 8861 29257 8895 29291
rect 8895 29257 8904 29291
rect 8852 29248 8904 29257
rect 15200 29248 15252 29300
rect 16948 29291 17000 29300
rect 16948 29257 16957 29291
rect 16957 29257 16991 29291
rect 16991 29257 17000 29291
rect 16948 29248 17000 29257
rect 12532 29223 12584 29232
rect 12532 29189 12541 29223
rect 12541 29189 12575 29223
rect 12575 29189 12584 29223
rect 12532 29180 12584 29189
rect 12624 29180 12676 29232
rect 16028 29223 16080 29232
rect 10968 29155 11020 29164
rect 10968 29121 10977 29155
rect 10977 29121 11011 29155
rect 11011 29121 11020 29155
rect 11704 29155 11756 29164
rect 10968 29112 11020 29121
rect 11704 29121 11713 29155
rect 11713 29121 11747 29155
rect 11747 29121 11756 29155
rect 11704 29112 11756 29121
rect 12808 29112 12860 29164
rect 7472 29087 7524 29096
rect 7472 29053 7481 29087
rect 7481 29053 7515 29087
rect 7515 29053 7524 29087
rect 7472 29044 7524 29053
rect 11888 29044 11940 29096
rect 12256 29044 12308 29096
rect 11520 29019 11572 29028
rect 11520 28985 11529 29019
rect 11529 28985 11563 29019
rect 11563 28985 11572 29019
rect 11520 28976 11572 28985
rect 16028 29189 16037 29223
rect 16037 29189 16071 29223
rect 16071 29189 16080 29223
rect 16028 29180 16080 29189
rect 17224 29248 17276 29300
rect 17408 29248 17460 29300
rect 20076 29248 20128 29300
rect 15200 29112 15252 29164
rect 19248 29180 19300 29232
rect 14740 29044 14792 29096
rect 17224 29155 17276 29164
rect 17224 29121 17233 29155
rect 17233 29121 17267 29155
rect 17267 29121 17276 29155
rect 17224 29112 17276 29121
rect 18420 29112 18472 29164
rect 18880 29112 18932 29164
rect 21180 29112 21232 29164
rect 17132 29044 17184 29096
rect 17408 29044 17460 29096
rect 19064 29087 19116 29096
rect 19064 29053 19073 29087
rect 19073 29053 19107 29087
rect 19107 29053 19116 29087
rect 19064 29044 19116 29053
rect 18880 28976 18932 29028
rect 19156 29019 19208 29028
rect 19156 28985 19165 29019
rect 19165 28985 19199 29019
rect 19199 28985 19208 29019
rect 19156 28976 19208 28985
rect 19432 28976 19484 29028
rect 13360 28908 13412 28960
rect 20536 28908 20588 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 12808 28747 12860 28756
rect 12808 28713 12817 28747
rect 12817 28713 12851 28747
rect 12851 28713 12860 28747
rect 12808 28704 12860 28713
rect 16488 28704 16540 28756
rect 18604 28747 18656 28756
rect 18604 28713 18613 28747
rect 18613 28713 18647 28747
rect 18647 28713 18656 28747
rect 18604 28704 18656 28713
rect 19340 28704 19392 28756
rect 11888 28636 11940 28688
rect 12440 28636 12492 28688
rect 10692 28500 10744 28552
rect 11796 28500 11848 28552
rect 16672 28500 16724 28552
rect 19432 28500 19484 28552
rect 12256 28432 12308 28484
rect 16856 28432 16908 28484
rect 18788 28432 18840 28484
rect 19248 28475 19300 28484
rect 19248 28441 19257 28475
rect 19257 28441 19291 28475
rect 19291 28441 19300 28475
rect 19248 28432 19300 28441
rect 2504 28364 2556 28416
rect 7472 28364 7524 28416
rect 9864 28407 9916 28416
rect 9864 28373 9873 28407
rect 9873 28373 9907 28407
rect 9907 28373 9916 28407
rect 9864 28364 9916 28373
rect 9956 28364 10008 28416
rect 18512 28364 18564 28416
rect 18696 28364 18748 28416
rect 20444 28364 20496 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 13360 28160 13412 28212
rect 13636 28203 13688 28212
rect 13636 28169 13645 28203
rect 13645 28169 13679 28203
rect 13679 28169 13688 28203
rect 13636 28160 13688 28169
rect 10048 28092 10100 28144
rect 12624 28092 12676 28144
rect 1400 28024 1452 28076
rect 2504 28067 2556 28076
rect 2504 28033 2513 28067
rect 2513 28033 2547 28067
rect 2547 28033 2556 28067
rect 2504 28024 2556 28033
rect 4068 28024 4120 28076
rect 9956 28024 10008 28076
rect 10692 28067 10744 28076
rect 10692 28033 10701 28067
rect 10701 28033 10735 28067
rect 10735 28033 10744 28067
rect 10692 28024 10744 28033
rect 11888 28024 11940 28076
rect 12348 28024 12400 28076
rect 14280 28067 14332 28076
rect 14280 28033 14289 28067
rect 14289 28033 14323 28067
rect 14323 28033 14332 28067
rect 14280 28024 14332 28033
rect 17868 28160 17920 28212
rect 18052 28160 18104 28212
rect 18236 28203 18288 28212
rect 18236 28169 18245 28203
rect 18245 28169 18279 28203
rect 18279 28169 18288 28203
rect 18236 28160 18288 28169
rect 18512 28160 18564 28212
rect 18604 28092 18656 28144
rect 17960 28024 18012 28076
rect 18144 28024 18196 28076
rect 18880 28067 18932 28076
rect 18880 28033 18889 28067
rect 18889 28033 18923 28067
rect 18923 28033 18932 28067
rect 18880 28024 18932 28033
rect 20536 28135 20588 28144
rect 20536 28101 20545 28135
rect 20545 28101 20579 28135
rect 20579 28101 20588 28135
rect 20536 28092 20588 28101
rect 10324 27956 10376 28008
rect 8392 27888 8444 27940
rect 10140 27820 10192 27872
rect 10876 27999 10928 28008
rect 10876 27965 10885 27999
rect 10885 27965 10919 27999
rect 10919 27965 10928 27999
rect 12256 27999 12308 28008
rect 10876 27956 10928 27965
rect 12256 27965 12265 27999
rect 12265 27965 12299 27999
rect 12299 27965 12308 27999
rect 12256 27956 12308 27965
rect 17776 27956 17828 28008
rect 16764 27888 16816 27940
rect 17500 27931 17552 27940
rect 17500 27897 17509 27931
rect 17509 27897 17543 27931
rect 17543 27897 17552 27931
rect 17500 27888 17552 27897
rect 19064 27888 19116 27940
rect 20444 27956 20496 28008
rect 20260 27888 20312 27940
rect 11980 27820 12032 27872
rect 15476 27863 15528 27872
rect 15476 27829 15485 27863
rect 15485 27829 15519 27863
rect 15519 27829 15528 27863
rect 15476 27820 15528 27829
rect 18420 27820 18472 27872
rect 19892 27820 19944 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 9864 27548 9916 27600
rect 10692 27548 10744 27600
rect 11796 27591 11848 27600
rect 11796 27557 11805 27591
rect 11805 27557 11839 27591
rect 11839 27557 11848 27591
rect 11796 27548 11848 27557
rect 18052 27616 18104 27668
rect 19432 27616 19484 27668
rect 17960 27548 18012 27600
rect 20536 27548 20588 27600
rect 21640 27591 21692 27600
rect 21640 27557 21649 27591
rect 21649 27557 21683 27591
rect 21683 27557 21692 27591
rect 21640 27548 21692 27557
rect 1400 27523 1452 27532
rect 1400 27489 1409 27523
rect 1409 27489 1443 27523
rect 1443 27489 1452 27523
rect 1400 27480 1452 27489
rect 2780 27480 2832 27532
rect 10876 27480 10928 27532
rect 14188 27480 14240 27532
rect 8392 27344 8444 27396
rect 3884 27276 3936 27328
rect 9956 27412 10008 27464
rect 12348 27412 12400 27464
rect 12992 27455 13044 27464
rect 12992 27421 13001 27455
rect 13001 27421 13035 27455
rect 13035 27421 13044 27455
rect 12992 27412 13044 27421
rect 16672 27412 16724 27464
rect 9864 27344 9916 27396
rect 11980 27344 12032 27396
rect 14464 27344 14516 27396
rect 15476 27344 15528 27396
rect 9404 27319 9456 27328
rect 9404 27285 9413 27319
rect 9413 27285 9447 27319
rect 9447 27285 9456 27319
rect 11336 27319 11388 27328
rect 9404 27276 9456 27285
rect 11336 27285 11345 27319
rect 11345 27285 11379 27319
rect 11379 27285 11388 27319
rect 11336 27276 11388 27285
rect 14740 27276 14792 27328
rect 15200 27319 15252 27328
rect 15200 27285 15209 27319
rect 15209 27285 15243 27319
rect 15243 27285 15252 27319
rect 15200 27276 15252 27285
rect 16028 27276 16080 27328
rect 19340 27480 19392 27532
rect 17132 27412 17184 27464
rect 19892 27455 19944 27464
rect 18420 27344 18472 27396
rect 19892 27421 19901 27455
rect 19901 27421 19935 27455
rect 19935 27421 19944 27455
rect 19892 27412 19944 27421
rect 22100 27412 22152 27464
rect 19708 27387 19760 27396
rect 19708 27353 19717 27387
rect 19717 27353 19751 27387
rect 19751 27353 19760 27387
rect 19708 27344 19760 27353
rect 20628 27387 20680 27396
rect 20628 27353 20637 27387
rect 20637 27353 20671 27387
rect 20671 27353 20680 27387
rect 20628 27344 20680 27353
rect 18880 27276 18932 27328
rect 19248 27276 19300 27328
rect 19524 27276 19576 27328
rect 21088 27319 21140 27328
rect 21088 27285 21097 27319
rect 21097 27285 21131 27319
rect 21131 27285 21140 27319
rect 21088 27276 21140 27285
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 9680 27115 9732 27124
rect 9680 27081 9689 27115
rect 9689 27081 9723 27115
rect 9723 27081 9732 27115
rect 9680 27072 9732 27081
rect 14280 27072 14332 27124
rect 15936 27072 15988 27124
rect 16120 27072 16172 27124
rect 7472 26936 7524 26988
rect 9864 26979 9916 26988
rect 9864 26945 9873 26979
rect 9873 26945 9907 26979
rect 9907 26945 9916 26979
rect 9864 26936 9916 26945
rect 9956 26979 10008 26988
rect 9956 26945 9965 26979
rect 9965 26945 9999 26979
rect 9999 26945 10008 26979
rect 11520 27004 11572 27056
rect 9956 26936 10008 26945
rect 10324 26979 10376 26988
rect 10324 26945 10333 26979
rect 10333 26945 10367 26979
rect 10367 26945 10376 26979
rect 10324 26936 10376 26945
rect 11888 27047 11940 27056
rect 11888 27013 11897 27047
rect 11897 27013 11931 27047
rect 11931 27013 11940 27047
rect 11888 27004 11940 27013
rect 12440 26936 12492 26988
rect 12532 26979 12584 26988
rect 12532 26945 12541 26979
rect 12541 26945 12575 26979
rect 12575 26945 12584 26979
rect 18880 27115 18932 27124
rect 18880 27081 18889 27115
rect 18889 27081 18923 27115
rect 18923 27081 18932 27115
rect 18880 27072 18932 27081
rect 19064 27115 19116 27124
rect 19064 27081 19073 27115
rect 19073 27081 19107 27115
rect 19107 27081 19116 27115
rect 19064 27072 19116 27081
rect 19432 27072 19484 27124
rect 19708 27072 19760 27124
rect 20628 27072 20680 27124
rect 19524 27004 19576 27056
rect 20812 27047 20864 27056
rect 20812 27013 20821 27047
rect 20821 27013 20855 27047
rect 20855 27013 20864 27047
rect 20812 27004 20864 27013
rect 20996 27004 21048 27056
rect 22652 27004 22704 27056
rect 12532 26936 12584 26945
rect 14832 26936 14884 26988
rect 15292 26936 15344 26988
rect 16672 26979 16724 26988
rect 16672 26945 16681 26979
rect 16681 26945 16715 26979
rect 16715 26945 16724 26979
rect 16672 26936 16724 26945
rect 16764 26936 16816 26988
rect 17500 26936 17552 26988
rect 17960 26936 18012 26988
rect 18052 26936 18104 26988
rect 19432 26936 19484 26988
rect 10140 26800 10192 26852
rect 11796 26800 11848 26852
rect 14556 26868 14608 26920
rect 16120 26868 16172 26920
rect 16580 26800 16632 26852
rect 18236 26800 18288 26852
rect 18788 26911 18840 26920
rect 18788 26877 18797 26911
rect 18797 26877 18831 26911
rect 18831 26877 18840 26911
rect 18788 26868 18840 26877
rect 19248 26868 19300 26920
rect 19616 26868 19668 26920
rect 22100 26979 22152 26988
rect 22100 26945 22109 26979
rect 22109 26945 22143 26979
rect 22143 26945 22152 26979
rect 22100 26936 22152 26945
rect 19708 26800 19760 26852
rect 9680 26732 9732 26784
rect 11888 26732 11940 26784
rect 13176 26732 13228 26784
rect 14832 26732 14884 26784
rect 17776 26732 17828 26784
rect 19064 26732 19116 26784
rect 19524 26732 19576 26784
rect 20720 26868 20772 26920
rect 20536 26800 20588 26852
rect 20812 26800 20864 26852
rect 20996 26800 21048 26852
rect 21640 26868 21692 26920
rect 20076 26732 20128 26784
rect 21364 26732 21416 26784
rect 21640 26732 21692 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 2780 26571 2832 26580
rect 2780 26537 2789 26571
rect 2789 26537 2823 26571
rect 2823 26537 2832 26571
rect 2780 26528 2832 26537
rect 8300 26528 8352 26580
rect 10048 26528 10100 26580
rect 11888 26571 11940 26580
rect 11888 26537 11897 26571
rect 11897 26537 11931 26571
rect 11931 26537 11940 26571
rect 11888 26528 11940 26537
rect 12532 26528 12584 26580
rect 17868 26528 17920 26580
rect 18880 26528 18932 26580
rect 19064 26528 19116 26580
rect 19616 26528 19668 26580
rect 19984 26528 20036 26580
rect 20536 26528 20588 26580
rect 1400 26435 1452 26444
rect 1400 26401 1409 26435
rect 1409 26401 1443 26435
rect 1443 26401 1452 26435
rect 1400 26392 1452 26401
rect 4068 26435 4120 26444
rect 4068 26401 4077 26435
rect 4077 26401 4111 26435
rect 4111 26401 4120 26435
rect 4068 26392 4120 26401
rect 9312 26324 9364 26376
rect 9680 26367 9732 26376
rect 9680 26333 9689 26367
rect 9689 26333 9723 26367
rect 9723 26333 9732 26367
rect 9680 26324 9732 26333
rect 13544 26392 13596 26444
rect 15108 26460 15160 26512
rect 17040 26460 17092 26512
rect 17316 26460 17368 26512
rect 18512 26503 18564 26512
rect 3884 26256 3936 26308
rect 8944 26299 8996 26308
rect 8944 26265 8953 26299
rect 8953 26265 8987 26299
rect 8987 26265 8996 26299
rect 8944 26256 8996 26265
rect 9772 26256 9824 26308
rect 13176 26324 13228 26376
rect 14832 26367 14884 26376
rect 14832 26333 14841 26367
rect 14841 26333 14875 26367
rect 14875 26333 14884 26367
rect 14832 26324 14884 26333
rect 13084 26256 13136 26308
rect 13636 26256 13688 26308
rect 13544 26231 13596 26240
rect 13544 26197 13553 26231
rect 13553 26197 13587 26231
rect 13587 26197 13596 26231
rect 13544 26188 13596 26197
rect 15200 26256 15252 26308
rect 16672 26392 16724 26444
rect 18512 26469 18521 26503
rect 18521 26469 18555 26503
rect 18555 26469 18564 26503
rect 18512 26460 18564 26469
rect 19248 26460 19300 26512
rect 19340 26392 19392 26444
rect 17040 26324 17092 26376
rect 17316 26256 17368 26308
rect 17500 26256 17552 26308
rect 17960 26299 18012 26308
rect 17960 26265 17969 26299
rect 17969 26265 18003 26299
rect 18003 26265 18012 26299
rect 17960 26256 18012 26265
rect 18788 26324 18840 26376
rect 21088 26460 21140 26512
rect 21272 26392 21324 26444
rect 21364 26367 21416 26376
rect 21364 26333 21373 26367
rect 21373 26333 21407 26367
rect 21407 26333 21416 26367
rect 21364 26324 21416 26333
rect 21640 26367 21692 26376
rect 21640 26333 21649 26367
rect 21649 26333 21683 26367
rect 21683 26333 21692 26367
rect 21640 26324 21692 26333
rect 22100 26367 22152 26376
rect 22100 26333 22109 26367
rect 22109 26333 22143 26367
rect 22143 26333 22152 26367
rect 22100 26324 22152 26333
rect 22652 26367 22704 26376
rect 22652 26333 22661 26367
rect 22661 26333 22695 26367
rect 22695 26333 22704 26367
rect 22652 26324 22704 26333
rect 22008 26188 22060 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 12992 26027 13044 26036
rect 12992 25993 13001 26027
rect 13001 25993 13035 26027
rect 13035 25993 13044 26027
rect 12992 25984 13044 25993
rect 9496 25848 9548 25900
rect 12256 25916 12308 25968
rect 7472 25780 7524 25832
rect 9680 25687 9732 25696
rect 9680 25653 9689 25687
rect 9689 25653 9723 25687
rect 9723 25653 9732 25687
rect 13820 25891 13872 25900
rect 13820 25857 13824 25891
rect 13824 25857 13858 25891
rect 13858 25857 13872 25891
rect 13820 25848 13872 25857
rect 15568 25984 15620 26036
rect 17500 25984 17552 26036
rect 18328 25984 18380 26036
rect 20812 25984 20864 26036
rect 22100 25984 22152 26036
rect 14004 25891 14056 25900
rect 14004 25857 14013 25891
rect 14013 25857 14047 25891
rect 14047 25857 14056 25891
rect 14004 25848 14056 25857
rect 14464 25848 14516 25900
rect 16672 25916 16724 25968
rect 15016 25891 15068 25900
rect 15016 25857 15050 25891
rect 15050 25857 15068 25891
rect 17132 25916 17184 25968
rect 19156 25916 19208 25968
rect 15016 25848 15068 25857
rect 17040 25891 17092 25900
rect 17040 25857 17049 25891
rect 17049 25857 17083 25891
rect 17083 25857 17092 25891
rect 17040 25848 17092 25857
rect 18052 25848 18104 25900
rect 20996 25848 21048 25900
rect 22008 25848 22060 25900
rect 22100 25891 22152 25900
rect 22100 25857 22109 25891
rect 22109 25857 22143 25891
rect 22143 25857 22152 25891
rect 22100 25848 22152 25857
rect 20352 25712 20404 25764
rect 9680 25644 9732 25653
rect 14924 25644 14976 25696
rect 16856 25644 16908 25696
rect 20168 25644 20220 25696
rect 20812 25644 20864 25696
rect 21732 25644 21784 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 8944 25440 8996 25492
rect 11428 25483 11480 25492
rect 11428 25449 11437 25483
rect 11437 25449 11471 25483
rect 11471 25449 11480 25483
rect 11428 25440 11480 25449
rect 12440 25440 12492 25492
rect 13728 25440 13780 25492
rect 13820 25440 13872 25492
rect 14556 25440 14608 25492
rect 17132 25440 17184 25492
rect 17224 25440 17276 25492
rect 17960 25440 18012 25492
rect 9312 25415 9364 25424
rect 9312 25381 9321 25415
rect 9321 25381 9355 25415
rect 9355 25381 9364 25415
rect 9312 25372 9364 25381
rect 9680 25372 9732 25424
rect 14648 25372 14700 25424
rect 19432 25440 19484 25492
rect 21732 25483 21784 25492
rect 10140 25304 10192 25356
rect 11980 25304 12032 25356
rect 9772 25236 9824 25288
rect 11704 25279 11756 25288
rect 11704 25245 11713 25279
rect 11713 25245 11747 25279
rect 11747 25245 11756 25279
rect 11704 25236 11756 25245
rect 13084 25236 13136 25288
rect 13544 25236 13596 25288
rect 13912 25236 13964 25288
rect 14556 25236 14608 25288
rect 16028 25279 16080 25288
rect 16028 25245 16037 25279
rect 16037 25245 16071 25279
rect 16071 25245 16080 25279
rect 16028 25236 16080 25245
rect 17316 25279 17368 25288
rect 13176 25211 13228 25220
rect 13176 25177 13185 25211
rect 13185 25177 13219 25211
rect 13219 25177 13228 25211
rect 13176 25168 13228 25177
rect 15200 25168 15252 25220
rect 17316 25245 17325 25279
rect 17325 25245 17359 25279
rect 17359 25245 17368 25279
rect 17316 25236 17368 25245
rect 18236 25279 18288 25288
rect 18236 25245 18245 25279
rect 18245 25245 18279 25279
rect 18279 25245 18288 25279
rect 18236 25236 18288 25245
rect 19800 25304 19852 25356
rect 20720 25372 20772 25424
rect 21732 25449 21741 25483
rect 21741 25449 21775 25483
rect 21775 25449 21784 25483
rect 21732 25440 21784 25449
rect 22100 25372 22152 25424
rect 15384 25100 15436 25152
rect 18604 25236 18656 25288
rect 19432 25236 19484 25288
rect 20536 25236 20588 25288
rect 20628 25236 20680 25288
rect 20720 25279 20772 25288
rect 20720 25245 20729 25279
rect 20729 25245 20763 25279
rect 20763 25245 20772 25279
rect 20720 25236 20772 25245
rect 20168 25168 20220 25220
rect 20260 25168 20312 25220
rect 18696 25100 18748 25152
rect 19432 25100 19484 25152
rect 19708 25143 19760 25152
rect 19708 25109 19717 25143
rect 19717 25109 19751 25143
rect 19751 25109 19760 25143
rect 19708 25100 19760 25109
rect 19800 25100 19852 25152
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 9772 24896 9824 24948
rect 12348 24939 12400 24948
rect 12348 24905 12357 24939
rect 12357 24905 12391 24939
rect 12391 24905 12400 24939
rect 12348 24896 12400 24905
rect 13544 24896 13596 24948
rect 18052 24939 18104 24948
rect 11796 24760 11848 24812
rect 9312 24692 9364 24744
rect 12532 24803 12584 24812
rect 12532 24769 12541 24803
rect 12541 24769 12575 24803
rect 12575 24769 12584 24803
rect 13912 24871 13964 24880
rect 13912 24837 13921 24871
rect 13921 24837 13955 24871
rect 13955 24837 13964 24871
rect 18052 24905 18061 24939
rect 18061 24905 18095 24939
rect 18095 24905 18104 24939
rect 18052 24896 18104 24905
rect 18144 24896 18196 24948
rect 13912 24828 13964 24837
rect 17408 24828 17460 24880
rect 12532 24760 12584 24769
rect 14832 24760 14884 24812
rect 16672 24803 16724 24812
rect 16672 24769 16681 24803
rect 16681 24769 16715 24803
rect 16715 24769 16724 24803
rect 16672 24760 16724 24769
rect 16948 24803 17000 24812
rect 16948 24769 16982 24803
rect 16982 24769 17000 24803
rect 16948 24760 17000 24769
rect 17316 24760 17368 24812
rect 18144 24760 18196 24812
rect 19340 24760 19392 24812
rect 19892 24828 19944 24880
rect 20168 24871 20220 24880
rect 20168 24837 20177 24871
rect 20177 24837 20211 24871
rect 20211 24837 20220 24871
rect 20168 24828 20220 24837
rect 21180 24828 21232 24880
rect 15108 24692 15160 24744
rect 9496 24624 9548 24676
rect 11796 24556 11848 24608
rect 12440 24556 12492 24608
rect 12624 24556 12676 24608
rect 13084 24556 13136 24608
rect 14096 24556 14148 24608
rect 14280 24556 14332 24608
rect 14464 24556 14516 24608
rect 19524 24692 19576 24744
rect 20076 24760 20128 24812
rect 20352 24803 20404 24812
rect 20352 24769 20361 24803
rect 20361 24769 20395 24803
rect 20395 24769 20404 24803
rect 20352 24760 20404 24769
rect 21916 24760 21968 24812
rect 23664 24803 23716 24812
rect 23664 24769 23673 24803
rect 23673 24769 23707 24803
rect 23707 24769 23716 24803
rect 23664 24760 23716 24769
rect 23940 24760 23992 24812
rect 24400 24803 24452 24812
rect 24400 24769 24409 24803
rect 24409 24769 24443 24803
rect 24443 24769 24452 24803
rect 24400 24760 24452 24769
rect 21732 24692 21784 24744
rect 19064 24556 19116 24608
rect 22008 24599 22060 24608
rect 22008 24565 22017 24599
rect 22017 24565 22051 24599
rect 22051 24565 22060 24599
rect 22008 24556 22060 24565
rect 23388 24556 23440 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 13544 24395 13596 24404
rect 13544 24361 13553 24395
rect 13553 24361 13587 24395
rect 13587 24361 13596 24395
rect 13544 24352 13596 24361
rect 14096 24395 14148 24404
rect 14096 24361 14105 24395
rect 14105 24361 14139 24395
rect 14139 24361 14148 24395
rect 14096 24352 14148 24361
rect 16948 24395 17000 24404
rect 16948 24361 16957 24395
rect 16957 24361 16991 24395
rect 16991 24361 17000 24395
rect 16948 24352 17000 24361
rect 17868 24352 17920 24404
rect 19340 24352 19392 24404
rect 20076 24395 20128 24404
rect 20076 24361 20085 24395
rect 20085 24361 20119 24395
rect 20119 24361 20128 24395
rect 20076 24352 20128 24361
rect 12532 24284 12584 24336
rect 13360 24284 13412 24336
rect 13912 24216 13964 24268
rect 13084 24191 13136 24200
rect 13084 24157 13093 24191
rect 13093 24157 13127 24191
rect 13127 24157 13136 24191
rect 13084 24148 13136 24157
rect 13176 24191 13228 24200
rect 13176 24157 13185 24191
rect 13185 24157 13219 24191
rect 13219 24157 13228 24191
rect 13176 24148 13228 24157
rect 13728 24148 13780 24200
rect 15108 24216 15160 24268
rect 17592 24284 17644 24336
rect 18420 24216 18472 24268
rect 18880 24216 18932 24268
rect 21732 24352 21784 24404
rect 20904 24284 20956 24336
rect 24400 24352 24452 24404
rect 22008 24284 22060 24336
rect 22376 24327 22428 24336
rect 22376 24293 22385 24327
rect 22385 24293 22419 24327
rect 22419 24293 22428 24327
rect 22376 24284 22428 24293
rect 23480 24327 23532 24336
rect 23480 24293 23489 24327
rect 23489 24293 23523 24327
rect 23523 24293 23532 24327
rect 23480 24284 23532 24293
rect 23388 24259 23440 24268
rect 23388 24225 23397 24259
rect 23397 24225 23431 24259
rect 23431 24225 23440 24259
rect 23388 24216 23440 24225
rect 12624 24080 12676 24132
rect 13452 24080 13504 24132
rect 14280 24080 14332 24132
rect 14648 24148 14700 24200
rect 16856 24191 16908 24200
rect 16856 24157 16865 24191
rect 16865 24157 16899 24191
rect 16899 24157 16908 24191
rect 16856 24148 16908 24157
rect 17132 24191 17184 24200
rect 17132 24157 17141 24191
rect 17141 24157 17175 24191
rect 17175 24157 17184 24191
rect 17132 24148 17184 24157
rect 18144 24080 18196 24132
rect 19524 24148 19576 24200
rect 20996 24148 21048 24200
rect 23572 24191 23624 24200
rect 23572 24157 23581 24191
rect 23581 24157 23615 24191
rect 23615 24157 23624 24191
rect 23572 24148 23624 24157
rect 20812 24080 20864 24132
rect 23204 24123 23256 24132
rect 23204 24089 23213 24123
rect 23213 24089 23247 24123
rect 23247 24089 23256 24123
rect 23204 24080 23256 24089
rect 18420 24055 18472 24064
rect 18420 24021 18447 24055
rect 18447 24021 18472 24055
rect 18420 24012 18472 24021
rect 19156 24012 19208 24064
rect 19432 24012 19484 24064
rect 19616 24012 19668 24064
rect 24308 24012 24360 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 13176 23808 13228 23860
rect 13084 23672 13136 23724
rect 13452 23740 13504 23792
rect 13820 23740 13872 23792
rect 13728 23715 13780 23724
rect 13728 23681 13737 23715
rect 13737 23681 13771 23715
rect 13771 23681 13780 23715
rect 13728 23672 13780 23681
rect 14188 23808 14240 23860
rect 17040 23808 17092 23860
rect 18420 23808 18472 23860
rect 18604 23808 18656 23860
rect 15752 23672 15804 23724
rect 16580 23672 16632 23724
rect 17960 23740 18012 23792
rect 18328 23740 18380 23792
rect 19064 23740 19116 23792
rect 20904 23808 20956 23860
rect 21916 23851 21968 23860
rect 21916 23817 21925 23851
rect 21925 23817 21959 23851
rect 21959 23817 21968 23851
rect 21916 23808 21968 23817
rect 20996 23740 21048 23792
rect 22192 23740 22244 23792
rect 17684 23672 17736 23724
rect 21732 23672 21784 23724
rect 22284 23715 22336 23724
rect 22284 23681 22293 23715
rect 22293 23681 22327 23715
rect 22327 23681 22336 23715
rect 22284 23672 22336 23681
rect 23940 23740 23992 23792
rect 23204 23672 23256 23724
rect 23388 23715 23440 23724
rect 23388 23681 23397 23715
rect 23397 23681 23431 23715
rect 23431 23681 23440 23715
rect 23388 23672 23440 23681
rect 23572 23672 23624 23724
rect 24308 23715 24360 23724
rect 10324 23604 10376 23656
rect 17132 23604 17184 23656
rect 20720 23604 20772 23656
rect 24308 23681 24317 23715
rect 24317 23681 24351 23715
rect 24351 23681 24360 23715
rect 24308 23672 24360 23681
rect 13820 23536 13872 23588
rect 15016 23536 15068 23588
rect 15200 23536 15252 23588
rect 22008 23536 22060 23588
rect 23480 23536 23532 23588
rect 15752 23511 15804 23520
rect 15752 23477 15761 23511
rect 15761 23477 15795 23511
rect 15795 23477 15804 23511
rect 15752 23468 15804 23477
rect 16856 23468 16908 23520
rect 19248 23468 19300 23520
rect 23112 23511 23164 23520
rect 23112 23477 23121 23511
rect 23121 23477 23155 23511
rect 23155 23477 23164 23511
rect 23112 23468 23164 23477
rect 24584 23511 24636 23520
rect 24584 23477 24593 23511
rect 24593 23477 24627 23511
rect 24627 23477 24636 23511
rect 24584 23468 24636 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 13452 23264 13504 23316
rect 15844 23264 15896 23316
rect 17408 23264 17460 23316
rect 13360 23239 13412 23248
rect 13360 23205 13369 23239
rect 13369 23205 13403 23239
rect 13403 23205 13412 23239
rect 13360 23196 13412 23205
rect 15292 23239 15344 23248
rect 15292 23205 15301 23239
rect 15301 23205 15335 23239
rect 15335 23205 15344 23239
rect 15292 23196 15344 23205
rect 15384 23196 15436 23248
rect 17316 23239 17368 23248
rect 11704 23128 11756 23180
rect 15844 23128 15896 23180
rect 17316 23205 17325 23239
rect 17325 23205 17359 23239
rect 17359 23205 17368 23239
rect 17316 23196 17368 23205
rect 17776 23239 17828 23248
rect 17776 23205 17785 23239
rect 17785 23205 17819 23239
rect 17819 23205 17828 23239
rect 17776 23196 17828 23205
rect 17868 23196 17920 23248
rect 19432 23264 19484 23316
rect 20720 23264 20772 23316
rect 22284 23264 22336 23316
rect 23204 23307 23256 23316
rect 23204 23273 23213 23307
rect 23213 23273 23247 23307
rect 23247 23273 23256 23307
rect 23204 23264 23256 23273
rect 18788 23128 18840 23180
rect 20260 23196 20312 23248
rect 21732 23196 21784 23248
rect 22376 23196 22428 23248
rect 22744 23171 22796 23180
rect 16028 23103 16080 23112
rect 16028 23069 16037 23103
rect 16037 23069 16071 23103
rect 16071 23069 16080 23103
rect 16028 23060 16080 23069
rect 16212 23103 16264 23112
rect 16212 23069 16221 23103
rect 16221 23069 16255 23103
rect 16255 23069 16264 23103
rect 16948 23103 17000 23112
rect 16212 23060 16264 23069
rect 16948 23069 16957 23103
rect 16957 23069 16991 23103
rect 16991 23069 17000 23103
rect 16948 23060 17000 23069
rect 16580 22992 16632 23044
rect 16856 22992 16908 23044
rect 18052 23060 18104 23112
rect 19064 23060 19116 23112
rect 20536 23103 20588 23112
rect 18144 23035 18196 23044
rect 18144 23001 18153 23035
rect 18153 23001 18187 23035
rect 18187 23001 18196 23035
rect 18144 22992 18196 23001
rect 18972 22992 19024 23044
rect 20536 23069 20545 23103
rect 20545 23069 20579 23103
rect 20579 23069 20588 23103
rect 20536 23060 20588 23069
rect 20996 23060 21048 23112
rect 22744 23137 22753 23171
rect 22753 23137 22787 23171
rect 22787 23137 22796 23171
rect 22744 23128 22796 23137
rect 21732 23060 21784 23112
rect 24584 23060 24636 23112
rect 14004 22924 14056 22976
rect 15108 22967 15160 22976
rect 15108 22933 15133 22967
rect 15133 22933 15160 22967
rect 15108 22924 15160 22933
rect 16672 22924 16724 22976
rect 17776 22924 17828 22976
rect 18788 22924 18840 22976
rect 19524 22924 19576 22976
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 14832 22763 14884 22772
rect 14832 22729 14841 22763
rect 14841 22729 14875 22763
rect 14875 22729 14884 22763
rect 14832 22720 14884 22729
rect 15108 22720 15160 22772
rect 16212 22720 16264 22772
rect 17132 22763 17184 22772
rect 17132 22729 17141 22763
rect 17141 22729 17175 22763
rect 17175 22729 17184 22763
rect 17132 22720 17184 22729
rect 17408 22763 17460 22772
rect 17408 22729 17417 22763
rect 17417 22729 17451 22763
rect 17451 22729 17460 22763
rect 17408 22720 17460 22729
rect 18052 22720 18104 22772
rect 16856 22652 16908 22704
rect 16948 22652 17000 22704
rect 14648 22584 14700 22636
rect 15016 22627 15068 22636
rect 15016 22593 15025 22627
rect 15025 22593 15059 22627
rect 15059 22593 15068 22627
rect 15016 22584 15068 22593
rect 15384 22584 15436 22636
rect 15844 22627 15896 22636
rect 15844 22593 15853 22627
rect 15853 22593 15887 22627
rect 15887 22593 15896 22627
rect 15844 22584 15896 22593
rect 20536 22720 20588 22772
rect 20720 22720 20772 22772
rect 22744 22720 22796 22772
rect 16028 22516 16080 22568
rect 15384 22380 15436 22432
rect 17960 22584 18012 22636
rect 18236 22627 18288 22636
rect 18236 22593 18245 22627
rect 18245 22593 18279 22627
rect 18279 22593 18288 22627
rect 18236 22584 18288 22593
rect 18972 22652 19024 22704
rect 19064 22652 19116 22704
rect 17868 22516 17920 22568
rect 18788 22584 18840 22636
rect 21180 22652 21232 22704
rect 18880 22559 18932 22568
rect 18880 22525 18889 22559
rect 18889 22525 18923 22559
rect 18923 22525 18932 22559
rect 18880 22516 18932 22525
rect 19064 22448 19116 22500
rect 20076 22448 20128 22500
rect 21272 22627 21324 22636
rect 21272 22593 21281 22627
rect 21281 22593 21315 22627
rect 21315 22593 21324 22627
rect 21272 22584 21324 22593
rect 21732 22584 21784 22636
rect 22008 22584 22060 22636
rect 20812 22516 20864 22568
rect 22192 22584 22244 22636
rect 21732 22448 21784 22500
rect 18236 22380 18288 22432
rect 19984 22380 20036 22432
rect 20260 22380 20312 22432
rect 20904 22380 20956 22432
rect 23296 22423 23348 22432
rect 23296 22389 23305 22423
rect 23305 22389 23339 22423
rect 23339 22389 23348 22423
rect 23296 22380 23348 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 16672 22219 16724 22228
rect 16672 22185 16681 22219
rect 16681 22185 16715 22219
rect 16715 22185 16724 22219
rect 16672 22176 16724 22185
rect 18144 22176 18196 22228
rect 18236 22176 18288 22228
rect 18972 22176 19024 22228
rect 19064 22176 19116 22228
rect 20352 22176 20404 22228
rect 20812 22108 20864 22160
rect 22652 22108 22704 22160
rect 23296 22108 23348 22160
rect 19248 21972 19300 22024
rect 19892 22015 19944 22024
rect 19892 21981 19901 22015
rect 19901 21981 19935 22015
rect 19935 21981 19944 22015
rect 19892 21972 19944 21981
rect 20536 22015 20588 22024
rect 20536 21981 20545 22015
rect 20545 21981 20579 22015
rect 20579 21981 20588 22015
rect 20536 21972 20588 21981
rect 20904 22015 20956 22024
rect 20904 21981 20913 22015
rect 20913 21981 20947 22015
rect 20947 21981 20956 22015
rect 20904 21972 20956 21981
rect 21548 21972 21600 22024
rect 20168 21904 20220 21956
rect 21272 21904 21324 21956
rect 22008 22015 22060 22024
rect 22008 21981 22017 22015
rect 22017 21981 22051 22015
rect 22051 21981 22060 22015
rect 22652 22015 22704 22024
rect 22008 21972 22060 21981
rect 22652 21981 22661 22015
rect 22661 21981 22695 22015
rect 22695 21981 22704 22015
rect 22652 21972 22704 21981
rect 23112 21972 23164 22024
rect 18328 21836 18380 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 18236 21675 18288 21684
rect 18236 21641 18245 21675
rect 18245 21641 18279 21675
rect 18279 21641 18288 21675
rect 18236 21632 18288 21641
rect 18880 21632 18932 21684
rect 19984 21632 20036 21684
rect 20812 21632 20864 21684
rect 23296 21632 23348 21684
rect 20536 21564 20588 21616
rect 19432 21496 19484 21548
rect 20076 21539 20128 21548
rect 20076 21505 20085 21539
rect 20085 21505 20119 21539
rect 20119 21505 20128 21539
rect 20076 21496 20128 21505
rect 20720 21496 20772 21548
rect 21088 21539 21140 21548
rect 21088 21505 21097 21539
rect 21097 21505 21131 21539
rect 21131 21505 21140 21539
rect 21088 21496 21140 21505
rect 21180 21539 21232 21548
rect 21180 21505 21189 21539
rect 21189 21505 21223 21539
rect 21223 21505 21232 21539
rect 21180 21496 21232 21505
rect 21548 21496 21600 21548
rect 22284 21496 22336 21548
rect 22652 21539 22704 21548
rect 22652 21505 22661 21539
rect 22661 21505 22695 21539
rect 22695 21505 22704 21539
rect 22652 21496 22704 21505
rect 23112 21496 23164 21548
rect 20444 21428 20496 21480
rect 22192 21428 22244 21480
rect 21088 21360 21140 21412
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 21548 21131 21600 21140
rect 21548 21097 21557 21131
rect 21557 21097 21591 21131
rect 21591 21097 21600 21131
rect 21548 21088 21600 21097
rect 22192 21131 22244 21140
rect 22192 21097 22201 21131
rect 22201 21097 22235 21131
rect 22235 21097 22244 21131
rect 22192 21088 22244 21097
rect 18696 21020 18748 21072
rect 19064 20952 19116 21004
rect 21180 21020 21232 21072
rect 19340 20927 19392 20936
rect 19340 20893 19349 20927
rect 19349 20893 19383 20927
rect 19383 20893 19392 20927
rect 19340 20884 19392 20893
rect 21088 20952 21140 21004
rect 20536 20884 20588 20936
rect 22284 20927 22336 20936
rect 22284 20893 22293 20927
rect 22293 20893 22327 20927
rect 22327 20893 22336 20927
rect 22284 20884 22336 20893
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 19064 20544 19116 20596
rect 20536 20544 20588 20596
rect 21180 20544 21232 20596
rect 22284 20544 22336 20596
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 9404 18368 9456 18420
rect 1400 18275 1452 18284
rect 1400 18241 1409 18275
rect 1409 18241 1443 18275
rect 1443 18241 1452 18275
rect 1400 18232 1452 18241
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 18512 12792 18564 12844
rect 37924 12588 37976 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 38108 12359 38160 12368
rect 38108 12325 38117 12359
rect 38117 12325 38151 12359
rect 38151 12325 38160 12359
rect 38108 12316 38160 12325
rect 37924 12223 37976 12232
rect 37924 12189 37933 12223
rect 37933 12189 37967 12223
rect 37967 12189 37976 12223
rect 37924 12180 37976 12189
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 20 2796 72 2848
rect 1400 2839 1452 2848
rect 1400 2805 1409 2839
rect 1409 2805 1443 2839
rect 1443 2805 1452 2839
rect 1400 2796 1452 2805
rect 34520 2796 34572 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 15752 2592 15804 2644
rect 1400 2499 1452 2508
rect 1400 2465 1409 2499
rect 1409 2465 1443 2499
rect 1443 2465 1452 2499
rect 1400 2456 1452 2465
rect 1676 2499 1728 2508
rect 1676 2465 1685 2499
rect 1685 2465 1719 2499
rect 1719 2465 1728 2499
rect 1676 2456 1728 2465
rect 11336 2456 11388 2508
rect 16764 2388 16816 2440
rect 34520 2320 34572 2372
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
<< metal2 >>
rect 13542 39200 13598 40000
rect 30930 39200 30986 40000
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 13556 37262 13584 39200
rect 30944 37466 30972 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 30932 37460 30984 37466
rect 30932 37402 30984 37408
rect 17776 37324 17828 37330
rect 17776 37266 17828 37272
rect 13544 37256 13596 37262
rect 13544 37198 13596 37204
rect 14280 37256 14332 37262
rect 14280 37198 14332 37204
rect 14292 36922 14320 37198
rect 14280 36916 14332 36922
rect 14280 36858 14332 36864
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 3422 36136 3478 36145
rect 3422 36071 3478 36080
rect 3436 36038 3464 36071
rect 3424 36032 3476 36038
rect 3424 35974 3476 35980
rect 9404 36032 9456 36038
rect 9404 35974 9456 35980
rect 8300 35760 8352 35766
rect 8300 35702 8352 35708
rect 6644 35692 6696 35698
rect 6644 35634 6696 35640
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 1676 31340 1728 31346
rect 1676 31282 1728 31288
rect 1400 31272 1452 31278
rect 1400 31214 1452 31220
rect 1412 28082 1440 31214
rect 1400 28076 1452 28082
rect 1400 28018 1452 28024
rect 1412 27538 1440 28018
rect 1400 27532 1452 27538
rect 1400 27474 1452 27480
rect 1412 26450 1440 27474
rect 1400 26444 1452 26450
rect 1400 26386 1452 26392
rect 1400 18284 1452 18290
rect 1400 18226 1452 18232
rect 1412 17785 1440 18226
rect 1398 17776 1454 17785
rect 1398 17711 1454 17720
rect 20 2848 72 2854
rect 20 2790 72 2796
rect 1400 2848 1452 2854
rect 1400 2790 1452 2796
rect 32 800 60 2790
rect 1412 2514 1440 2790
rect 1688 2514 1716 31282
rect 2780 31136 2832 31142
rect 2780 31078 2832 31084
rect 2504 28416 2556 28422
rect 2504 28358 2556 28364
rect 2516 28082 2544 28358
rect 2504 28076 2556 28082
rect 2504 28018 2556 28024
rect 2792 27985 2820 31078
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 6656 30054 6684 35634
rect 8312 31754 8340 35702
rect 8300 31748 8352 31754
rect 8300 31690 8352 31696
rect 8312 31482 8340 31690
rect 8300 31476 8352 31482
rect 8300 31418 8352 31424
rect 8300 31340 8352 31346
rect 8300 31282 8352 31288
rect 7472 31272 7524 31278
rect 7472 31214 7524 31220
rect 6644 30048 6696 30054
rect 6644 29990 6696 29996
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 7484 29102 7512 31214
rect 7472 29096 7524 29102
rect 7472 29038 7524 29044
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 7484 28422 7512 29038
rect 7472 28416 7524 28422
rect 7472 28358 7524 28364
rect 4068 28076 4120 28082
rect 4068 28018 4120 28024
rect 2778 27976 2834 27985
rect 2778 27911 2834 27920
rect 2780 27532 2832 27538
rect 2780 27474 2832 27480
rect 2792 26586 2820 27474
rect 4080 27441 4108 28018
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4066 27432 4122 27441
rect 4066 27367 4122 27376
rect 3884 27328 3936 27334
rect 3884 27270 3936 27276
rect 2780 26580 2832 26586
rect 2780 26522 2832 26528
rect 3896 26314 3924 27270
rect 7484 26994 7512 28358
rect 7472 26988 7524 26994
rect 7472 26930 7524 26936
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4066 26480 4122 26489
rect 4066 26415 4068 26424
rect 4120 26415 4122 26424
rect 4068 26386 4120 26392
rect 3884 26308 3936 26314
rect 3884 26250 3936 26256
rect 7484 25838 7512 26930
rect 8312 26586 8340 31282
rect 9416 30734 9444 35974
rect 17224 35692 17276 35698
rect 17224 35634 17276 35640
rect 17132 35080 17184 35086
rect 17052 35028 17132 35034
rect 17052 35022 17184 35028
rect 16764 35012 16816 35018
rect 16764 34954 16816 34960
rect 17052 35006 17172 35022
rect 16672 33924 16724 33930
rect 16672 33866 16724 33872
rect 15844 33856 15896 33862
rect 15844 33798 15896 33804
rect 15856 33454 15884 33798
rect 16684 33658 16712 33866
rect 16672 33652 16724 33658
rect 16672 33594 16724 33600
rect 16488 33516 16540 33522
rect 16488 33458 16540 33464
rect 14188 33448 14240 33454
rect 14188 33390 14240 33396
rect 15844 33448 15896 33454
rect 15844 33390 15896 33396
rect 16028 33448 16080 33454
rect 16028 33390 16080 33396
rect 14200 32978 14228 33390
rect 15108 33312 15160 33318
rect 15108 33254 15160 33260
rect 14188 32972 14240 32978
rect 14188 32914 14240 32920
rect 13820 32904 13872 32910
rect 13820 32846 13872 32852
rect 11520 32768 11572 32774
rect 11520 32710 11572 32716
rect 11532 32026 11560 32710
rect 11520 32020 11572 32026
rect 11520 31962 11572 31968
rect 9680 31816 9732 31822
rect 9680 31758 9732 31764
rect 9404 30728 9456 30734
rect 9404 30670 9456 30676
rect 9416 30394 9444 30670
rect 9404 30388 9456 30394
rect 9404 30330 9456 30336
rect 8852 29572 8904 29578
rect 8852 29514 8904 29520
rect 8864 29306 8892 29514
rect 8852 29300 8904 29306
rect 8852 29242 8904 29248
rect 8392 27940 8444 27946
rect 8392 27882 8444 27888
rect 8404 27402 8432 27882
rect 8392 27396 8444 27402
rect 8392 27338 8444 27344
rect 9404 27328 9456 27334
rect 9404 27270 9456 27276
rect 8300 26580 8352 26586
rect 8300 26522 8352 26528
rect 9312 26376 9364 26382
rect 9312 26318 9364 26324
rect 8944 26308 8996 26314
rect 8944 26250 8996 26256
rect 7472 25832 7524 25838
rect 7472 25774 7524 25780
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 8956 25498 8984 26250
rect 8944 25492 8996 25498
rect 8944 25434 8996 25440
rect 9324 25430 9352 26318
rect 9312 25424 9364 25430
rect 9312 25366 9364 25372
rect 9324 24750 9352 25366
rect 9312 24744 9364 24750
rect 9312 24686 9364 24692
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 9416 18426 9444 27270
rect 9692 27130 9720 31758
rect 10968 31680 11020 31686
rect 10968 31622 11020 31628
rect 9772 31136 9824 31142
rect 9772 31078 9824 31084
rect 9680 27124 9732 27130
rect 9680 27066 9732 27072
rect 9680 26784 9732 26790
rect 9680 26726 9732 26732
rect 9692 26382 9720 26726
rect 9680 26376 9732 26382
rect 9680 26318 9732 26324
rect 9784 26314 9812 31078
rect 10692 30592 10744 30598
rect 10692 30534 10744 30540
rect 10704 28558 10732 30534
rect 10980 29170 11008 31622
rect 13832 30802 13860 32846
rect 13820 30796 13872 30802
rect 13820 30738 13872 30744
rect 11428 30660 11480 30666
rect 11428 30602 11480 30608
rect 10968 29164 11020 29170
rect 10968 29106 11020 29112
rect 10692 28552 10744 28558
rect 10692 28494 10744 28500
rect 9864 28416 9916 28422
rect 9864 28358 9916 28364
rect 9956 28416 10008 28422
rect 9956 28358 10008 28364
rect 9876 27606 9904 28358
rect 9968 28082 9996 28358
rect 10048 28144 10100 28150
rect 10048 28086 10100 28092
rect 9956 28076 10008 28082
rect 9956 28018 10008 28024
rect 9864 27600 9916 27606
rect 9864 27542 9916 27548
rect 9956 27464 10008 27470
rect 9956 27406 10008 27412
rect 9864 27396 9916 27402
rect 9864 27338 9916 27344
rect 9876 26994 9904 27338
rect 9968 26994 9996 27406
rect 9864 26988 9916 26994
rect 9864 26930 9916 26936
rect 9956 26988 10008 26994
rect 9956 26930 10008 26936
rect 10060 26586 10088 28086
rect 10692 28076 10744 28082
rect 10692 28018 10744 28024
rect 10324 28008 10376 28014
rect 10324 27950 10376 27956
rect 10140 27872 10192 27878
rect 10140 27814 10192 27820
rect 10152 26858 10180 27814
rect 10336 26994 10364 27950
rect 10704 27606 10732 28018
rect 10876 28008 10928 28014
rect 10876 27950 10928 27956
rect 10692 27600 10744 27606
rect 10692 27542 10744 27548
rect 10888 27538 10916 27950
rect 10876 27532 10928 27538
rect 10876 27474 10928 27480
rect 11336 27328 11388 27334
rect 11336 27270 11388 27276
rect 10324 26988 10376 26994
rect 10324 26930 10376 26936
rect 10140 26852 10192 26858
rect 10140 26794 10192 26800
rect 10048 26580 10100 26586
rect 10048 26522 10100 26528
rect 9772 26308 9824 26314
rect 9772 26250 9824 26256
rect 9496 25900 9548 25906
rect 9496 25842 9548 25848
rect 9508 24682 9536 25842
rect 9680 25696 9732 25702
rect 9680 25638 9732 25644
rect 9692 25430 9720 25638
rect 9680 25424 9732 25430
rect 9680 25366 9732 25372
rect 9784 25294 9812 26250
rect 10152 25362 10180 26794
rect 10140 25356 10192 25362
rect 10140 25298 10192 25304
rect 9772 25288 9824 25294
rect 9772 25230 9824 25236
rect 9784 24954 9812 25230
rect 9772 24948 9824 24954
rect 9772 24890 9824 24896
rect 9496 24676 9548 24682
rect 9496 24618 9548 24624
rect 10336 23662 10364 26930
rect 10324 23656 10376 23662
rect 10324 23598 10376 23604
rect 9404 18420 9456 18426
rect 9404 18362 9456 18368
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 11348 2514 11376 27270
rect 11440 25498 11468 30602
rect 12532 29844 12584 29850
rect 12532 29786 12584 29792
rect 13820 29844 13872 29850
rect 13820 29786 13872 29792
rect 11888 29776 11940 29782
rect 11888 29718 11940 29724
rect 11900 29510 11928 29718
rect 12440 29640 12492 29646
rect 12440 29582 12492 29588
rect 11888 29504 11940 29510
rect 11888 29446 11940 29452
rect 11702 29200 11758 29209
rect 11702 29135 11704 29144
rect 11756 29135 11758 29144
rect 11704 29106 11756 29112
rect 11900 29102 11928 29446
rect 11888 29096 11940 29102
rect 11888 29038 11940 29044
rect 12256 29096 12308 29102
rect 12256 29038 12308 29044
rect 11520 29028 11572 29034
rect 11520 28970 11572 28976
rect 11532 27062 11560 28970
rect 11900 28694 11928 29038
rect 11888 28688 11940 28694
rect 11888 28630 11940 28636
rect 11796 28552 11848 28558
rect 11796 28494 11848 28500
rect 11808 27606 11836 28494
rect 11900 28082 11928 28630
rect 12268 28490 12296 29038
rect 12452 28694 12480 29582
rect 12544 29238 12572 29786
rect 12532 29232 12584 29238
rect 12532 29174 12584 29180
rect 12624 29232 12676 29238
rect 12624 29174 12676 29180
rect 12440 28688 12492 28694
rect 12440 28630 12492 28636
rect 12256 28484 12308 28490
rect 12256 28426 12308 28432
rect 11888 28076 11940 28082
rect 11888 28018 11940 28024
rect 12268 28014 12296 28426
rect 12636 28150 12664 29174
rect 12808 29164 12860 29170
rect 12808 29106 12860 29112
rect 12820 28762 12848 29106
rect 13360 28960 13412 28966
rect 13360 28902 13412 28908
rect 13634 28928 13690 28937
rect 12808 28756 12860 28762
rect 12808 28698 12860 28704
rect 13372 28218 13400 28902
rect 13634 28863 13690 28872
rect 13648 28218 13676 28863
rect 13360 28212 13412 28218
rect 13360 28154 13412 28160
rect 13636 28212 13688 28218
rect 13636 28154 13688 28160
rect 12624 28144 12676 28150
rect 12624 28086 12676 28092
rect 12348 28076 12400 28082
rect 12348 28018 12400 28024
rect 12256 28008 12308 28014
rect 12256 27950 12308 27956
rect 11980 27872 12032 27878
rect 11980 27814 12032 27820
rect 11796 27600 11848 27606
rect 11796 27542 11848 27548
rect 11992 27402 12020 27814
rect 11980 27396 12032 27402
rect 11980 27338 12032 27344
rect 11520 27056 11572 27062
rect 11520 26998 11572 27004
rect 11888 27056 11940 27062
rect 11888 26998 11940 27004
rect 11900 26874 11928 26998
rect 11808 26858 11928 26874
rect 11796 26852 11928 26858
rect 11848 26846 11928 26852
rect 11796 26794 11848 26800
rect 11888 26784 11940 26790
rect 11888 26726 11940 26732
rect 11900 26586 11928 26726
rect 11888 26580 11940 26586
rect 11888 26522 11940 26528
rect 11428 25492 11480 25498
rect 11428 25434 11480 25440
rect 11992 25362 12020 27338
rect 12268 25974 12296 27950
rect 12360 27470 12388 28018
rect 12348 27464 12400 27470
rect 12348 27406 12400 27412
rect 12992 27464 13044 27470
rect 12992 27406 13044 27412
rect 12440 26988 12492 26994
rect 12440 26930 12492 26936
rect 12532 26988 12584 26994
rect 12532 26930 12584 26936
rect 12256 25968 12308 25974
rect 12256 25910 12308 25916
rect 12452 25498 12480 26930
rect 12544 26586 12572 26930
rect 12532 26580 12584 26586
rect 12532 26522 12584 26528
rect 13004 26042 13032 27406
rect 13176 26784 13228 26790
rect 13176 26726 13228 26732
rect 13188 26382 13216 26726
rect 13544 26444 13596 26450
rect 13544 26386 13596 26392
rect 13176 26376 13228 26382
rect 13176 26318 13228 26324
rect 13084 26308 13136 26314
rect 13084 26250 13136 26256
rect 12992 26036 13044 26042
rect 12992 25978 13044 25984
rect 12440 25492 12492 25498
rect 12440 25434 12492 25440
rect 11980 25356 12032 25362
rect 11980 25298 12032 25304
rect 13096 25294 13124 26250
rect 11704 25288 11756 25294
rect 11704 25230 11756 25236
rect 13084 25288 13136 25294
rect 13084 25230 13136 25236
rect 11716 23186 11744 25230
rect 13188 25226 13216 26318
rect 13556 26246 13584 26386
rect 13648 26314 13676 28154
rect 13636 26308 13688 26314
rect 13636 26250 13688 26256
rect 13544 26240 13596 26246
rect 13544 26182 13596 26188
rect 13556 25294 13584 26182
rect 13832 25906 13860 29786
rect 14200 27538 14228 32914
rect 15016 32836 15068 32842
rect 15016 32778 15068 32784
rect 14372 32768 14424 32774
rect 14372 32710 14424 32716
rect 14464 32768 14516 32774
rect 14464 32710 14516 32716
rect 14648 32768 14700 32774
rect 14648 32710 14700 32716
rect 14384 32298 14412 32710
rect 14372 32292 14424 32298
rect 14372 32234 14424 32240
rect 14476 30394 14504 32710
rect 14660 32434 14688 32710
rect 14648 32428 14700 32434
rect 14648 32370 14700 32376
rect 14924 32224 14976 32230
rect 14924 32166 14976 32172
rect 14936 31754 14964 32166
rect 15028 32026 15056 32778
rect 15016 32020 15068 32026
rect 15016 31962 15068 31968
rect 15120 31822 15148 33254
rect 15856 33114 15884 33390
rect 16040 33318 16068 33390
rect 16028 33312 16080 33318
rect 16028 33254 16080 33260
rect 15844 33108 15896 33114
rect 15844 33050 15896 33056
rect 15936 32836 15988 32842
rect 15936 32778 15988 32784
rect 15752 32360 15804 32366
rect 15752 32302 15804 32308
rect 15568 31884 15620 31890
rect 15568 31826 15620 31832
rect 15108 31816 15160 31822
rect 15108 31758 15160 31764
rect 14936 31726 15056 31754
rect 14464 30388 14516 30394
rect 14464 30330 14516 30336
rect 14924 30388 14976 30394
rect 14924 30330 14976 30336
rect 14740 29572 14792 29578
rect 14740 29514 14792 29520
rect 14752 29102 14780 29514
rect 14740 29096 14792 29102
rect 14740 29038 14792 29044
rect 14280 28076 14332 28082
rect 14280 28018 14332 28024
rect 14188 27532 14240 27538
rect 14188 27474 14240 27480
rect 13820 25900 13872 25906
rect 13820 25842 13872 25848
rect 14004 25900 14056 25906
rect 14004 25842 14056 25848
rect 13832 25498 13860 25842
rect 13728 25492 13780 25498
rect 13728 25434 13780 25440
rect 13820 25492 13872 25498
rect 13820 25434 13872 25440
rect 13544 25288 13596 25294
rect 13544 25230 13596 25236
rect 13176 25220 13228 25226
rect 13176 25162 13228 25168
rect 13556 24954 13584 25230
rect 12348 24948 12400 24954
rect 12348 24890 12400 24896
rect 13544 24948 13596 24954
rect 13544 24890 13596 24896
rect 11796 24812 11848 24818
rect 12360 24800 12388 24890
rect 12532 24812 12584 24818
rect 12360 24772 12480 24800
rect 11796 24754 11848 24760
rect 11808 24614 11836 24754
rect 12452 24614 12480 24772
rect 12532 24754 12584 24760
rect 11796 24608 11848 24614
rect 11796 24550 11848 24556
rect 12440 24608 12492 24614
rect 12440 24550 12492 24556
rect 12544 24342 12572 24754
rect 12624 24608 12676 24614
rect 12624 24550 12676 24556
rect 13084 24608 13136 24614
rect 13084 24550 13136 24556
rect 12532 24336 12584 24342
rect 12532 24278 12584 24284
rect 12636 24138 12664 24550
rect 13096 24206 13124 24550
rect 13542 24440 13598 24449
rect 13542 24375 13544 24384
rect 13596 24375 13598 24384
rect 13544 24346 13596 24352
rect 13360 24336 13412 24342
rect 13360 24278 13412 24284
rect 13084 24200 13136 24206
rect 13084 24142 13136 24148
rect 13176 24200 13228 24206
rect 13176 24142 13228 24148
rect 12624 24132 12676 24138
rect 12624 24074 12676 24080
rect 13188 23866 13216 24142
rect 13176 23860 13228 23866
rect 13176 23802 13228 23808
rect 13084 23724 13136 23730
rect 13372 23712 13400 24278
rect 13740 24206 13768 25434
rect 13912 25288 13964 25294
rect 13912 25230 13964 25236
rect 13924 24886 13952 25230
rect 13912 24880 13964 24886
rect 13912 24822 13964 24828
rect 13924 24274 13952 24822
rect 13912 24268 13964 24274
rect 13912 24210 13964 24216
rect 13728 24200 13780 24206
rect 13728 24142 13780 24148
rect 13452 24132 13504 24138
rect 13452 24074 13504 24080
rect 13464 23798 13492 24074
rect 13452 23792 13504 23798
rect 13452 23734 13504 23740
rect 13136 23684 13400 23712
rect 13084 23666 13136 23672
rect 13372 23254 13400 23684
rect 13464 23322 13492 23734
rect 13740 23730 13768 24142
rect 13820 23792 13872 23798
rect 13818 23760 13820 23769
rect 13872 23760 13874 23769
rect 13728 23724 13780 23730
rect 13818 23695 13874 23704
rect 13728 23666 13780 23672
rect 13832 23594 13860 23695
rect 13820 23588 13872 23594
rect 13820 23530 13872 23536
rect 13452 23316 13504 23322
rect 13452 23258 13504 23264
rect 13360 23248 13412 23254
rect 13360 23190 13412 23196
rect 11704 23180 11756 23186
rect 11704 23122 11756 23128
rect 14016 22982 14044 25842
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 14108 24410 14136 24550
rect 14096 24404 14148 24410
rect 14096 24346 14148 24352
rect 14200 23866 14228 27474
rect 14292 27130 14320 28018
rect 14464 27396 14516 27402
rect 14464 27338 14516 27344
rect 14280 27124 14332 27130
rect 14280 27066 14332 27072
rect 14476 25906 14504 27338
rect 14752 27334 14780 29038
rect 14740 27328 14792 27334
rect 14740 27270 14792 27276
rect 14556 26920 14608 26926
rect 14556 26862 14608 26868
rect 14464 25900 14516 25906
rect 14464 25842 14516 25848
rect 14476 24614 14504 25842
rect 14568 25498 14596 26862
rect 14752 26364 14780 27270
rect 14832 26988 14884 26994
rect 14832 26930 14884 26936
rect 14844 26790 14872 26930
rect 14832 26784 14884 26790
rect 14832 26726 14884 26732
rect 14832 26376 14884 26382
rect 14752 26336 14832 26364
rect 14556 25492 14608 25498
rect 14556 25434 14608 25440
rect 14568 25294 14596 25434
rect 14648 25424 14700 25430
rect 14648 25366 14700 25372
rect 14556 25288 14608 25294
rect 14556 25230 14608 25236
rect 14280 24608 14332 24614
rect 14280 24550 14332 24556
rect 14464 24608 14516 24614
rect 14464 24550 14516 24556
rect 14292 24138 14320 24550
rect 14660 24206 14688 25366
rect 14648 24200 14700 24206
rect 14648 24142 14700 24148
rect 14280 24132 14332 24138
rect 14280 24074 14332 24080
rect 14188 23860 14240 23866
rect 14188 23802 14240 23808
rect 14660 23225 14688 24142
rect 14752 23769 14780 26336
rect 14832 26318 14884 26324
rect 14936 25702 14964 30330
rect 15028 25906 15056 31726
rect 15384 30592 15436 30598
rect 15384 30534 15436 30540
rect 15200 29572 15252 29578
rect 15200 29514 15252 29520
rect 15108 29504 15160 29510
rect 15108 29446 15160 29452
rect 15120 26518 15148 29446
rect 15212 29306 15240 29514
rect 15200 29300 15252 29306
rect 15200 29242 15252 29248
rect 15200 29164 15252 29170
rect 15200 29106 15252 29112
rect 15212 27334 15240 29106
rect 15200 27328 15252 27334
rect 15200 27270 15252 27276
rect 15108 26512 15160 26518
rect 15108 26454 15160 26460
rect 15016 25900 15068 25906
rect 15016 25842 15068 25848
rect 14924 25696 14976 25702
rect 14924 25638 14976 25644
rect 14832 24812 14884 24818
rect 14832 24754 14884 24760
rect 14738 23760 14794 23769
rect 14738 23695 14794 23704
rect 14646 23216 14702 23225
rect 14646 23151 14702 23160
rect 14004 22976 14056 22982
rect 14004 22918 14056 22924
rect 14660 22642 14688 23151
rect 14844 22778 14872 24754
rect 15120 24750 15148 26454
rect 15212 26314 15240 27270
rect 15292 26988 15344 26994
rect 15292 26930 15344 26936
rect 15200 26308 15252 26314
rect 15200 26250 15252 26256
rect 15212 25226 15240 26250
rect 15200 25220 15252 25226
rect 15200 25162 15252 25168
rect 15108 24744 15160 24750
rect 15108 24686 15160 24692
rect 15120 24274 15148 24686
rect 15108 24268 15160 24274
rect 15108 24210 15160 24216
rect 15212 23594 15240 25162
rect 15016 23588 15068 23594
rect 15016 23530 15068 23536
rect 15200 23588 15252 23594
rect 15200 23530 15252 23536
rect 14832 22772 14884 22778
rect 14832 22714 14884 22720
rect 15028 22642 15056 23530
rect 15304 23254 15332 26930
rect 15396 25158 15424 30534
rect 15580 29510 15608 31826
rect 15764 31822 15792 32302
rect 15752 31816 15804 31822
rect 15752 31758 15804 31764
rect 15764 29850 15792 31758
rect 15752 29844 15804 29850
rect 15752 29786 15804 29792
rect 15764 29578 15792 29786
rect 15752 29572 15804 29578
rect 15752 29514 15804 29520
rect 15568 29504 15620 29510
rect 15568 29446 15620 29452
rect 15476 27872 15528 27878
rect 15476 27814 15528 27820
rect 15488 27402 15516 27814
rect 15476 27396 15528 27402
rect 15476 27338 15528 27344
rect 15580 26042 15608 29446
rect 15948 27130 15976 32778
rect 16304 31748 16356 31754
rect 16304 31690 16356 31696
rect 16316 29850 16344 31690
rect 16500 31210 16528 33458
rect 16672 33380 16724 33386
rect 16672 33322 16724 33328
rect 16684 32434 16712 33322
rect 16672 32428 16724 32434
rect 16672 32370 16724 32376
rect 16776 31482 16804 34954
rect 16948 34604 17000 34610
rect 16948 34546 17000 34552
rect 16856 32224 16908 32230
rect 16856 32166 16908 32172
rect 16764 31476 16816 31482
rect 16764 31418 16816 31424
rect 16488 31204 16540 31210
rect 16488 31146 16540 31152
rect 16304 29844 16356 29850
rect 16304 29786 16356 29792
rect 16028 29504 16080 29510
rect 16028 29446 16080 29452
rect 16040 29238 16068 29446
rect 16028 29232 16080 29238
rect 16028 29174 16080 29180
rect 16500 28762 16528 31146
rect 16672 30728 16724 30734
rect 16672 30670 16724 30676
rect 16580 30320 16632 30326
rect 16580 30262 16632 30268
rect 16488 28756 16540 28762
rect 16488 28698 16540 28704
rect 16028 27328 16080 27334
rect 16028 27270 16080 27276
rect 15936 27124 15988 27130
rect 15936 27066 15988 27072
rect 15568 26036 15620 26042
rect 15568 25978 15620 25984
rect 16040 25294 16068 27270
rect 16120 27124 16172 27130
rect 16120 27066 16172 27072
rect 16132 26926 16160 27066
rect 16120 26920 16172 26926
rect 16120 26862 16172 26868
rect 16592 26858 16620 30262
rect 16684 30258 16712 30670
rect 16672 30252 16724 30258
rect 16672 30194 16724 30200
rect 16684 28558 16712 30194
rect 16672 28552 16724 28558
rect 16672 28494 16724 28500
rect 16684 27470 16712 28494
rect 16868 28490 16896 32166
rect 16960 31754 16988 34546
rect 17052 34406 17080 35006
rect 17132 34944 17184 34950
rect 17132 34886 17184 34892
rect 17040 34400 17092 34406
rect 17040 34342 17092 34348
rect 17052 33998 17080 34342
rect 17040 33992 17092 33998
rect 17040 33934 17092 33940
rect 17052 32910 17080 33934
rect 17040 32904 17092 32910
rect 17040 32846 17092 32852
rect 16960 31726 17080 31754
rect 16948 31340 17000 31346
rect 16948 31282 17000 31288
rect 16960 30938 16988 31282
rect 16948 30932 17000 30938
rect 16948 30874 17000 30880
rect 16948 29640 17000 29646
rect 16948 29582 17000 29588
rect 16960 29306 16988 29582
rect 16948 29300 17000 29306
rect 16948 29242 17000 29248
rect 16856 28484 16908 28490
rect 16856 28426 16908 28432
rect 16764 27940 16816 27946
rect 16764 27882 16816 27888
rect 16672 27464 16724 27470
rect 16672 27406 16724 27412
rect 16684 26994 16712 27406
rect 16776 26994 16804 27882
rect 16672 26988 16724 26994
rect 16672 26930 16724 26936
rect 16764 26988 16816 26994
rect 16764 26930 16816 26936
rect 16580 26852 16632 26858
rect 16580 26794 16632 26800
rect 16684 26450 16712 26930
rect 17052 26602 17080 31726
rect 17144 31346 17172 34886
rect 17236 32026 17264 35634
rect 17684 35488 17736 35494
rect 17684 35430 17736 35436
rect 17316 34196 17368 34202
rect 17316 34138 17368 34144
rect 17328 33318 17356 34138
rect 17316 33312 17368 33318
rect 17316 33254 17368 33260
rect 17328 32026 17356 33254
rect 17592 32768 17644 32774
rect 17592 32710 17644 32716
rect 17224 32020 17276 32026
rect 17224 31962 17276 31968
rect 17316 32020 17368 32026
rect 17316 31962 17368 31968
rect 17224 31884 17276 31890
rect 17224 31826 17276 31832
rect 17236 31482 17264 31826
rect 17224 31476 17276 31482
rect 17224 31418 17276 31424
rect 17132 31340 17184 31346
rect 17132 31282 17184 31288
rect 17144 30734 17172 31282
rect 17132 30728 17184 30734
rect 17132 30670 17184 30676
rect 17132 29844 17184 29850
rect 17132 29786 17184 29792
rect 17144 29102 17172 29786
rect 17224 29504 17276 29510
rect 17328 29492 17356 31962
rect 17276 29464 17356 29492
rect 17224 29446 17276 29452
rect 17236 29306 17264 29446
rect 17224 29300 17276 29306
rect 17224 29242 17276 29248
rect 17408 29300 17460 29306
rect 17408 29242 17460 29248
rect 17420 29209 17448 29242
rect 17406 29200 17462 29209
rect 17224 29164 17276 29170
rect 17406 29135 17462 29144
rect 17224 29106 17276 29112
rect 17132 29096 17184 29102
rect 17132 29038 17184 29044
rect 17236 28937 17264 29106
rect 17408 29096 17460 29102
rect 17408 29038 17460 29044
rect 17222 28928 17278 28937
rect 17222 28863 17278 28872
rect 17132 27464 17184 27470
rect 17132 27406 17184 27412
rect 16776 26574 17080 26602
rect 16672 26444 16724 26450
rect 16672 26386 16724 26392
rect 16684 25974 16712 26386
rect 16672 25968 16724 25974
rect 16672 25910 16724 25916
rect 16028 25288 16080 25294
rect 16028 25230 16080 25236
rect 15384 25152 15436 25158
rect 15384 25094 15436 25100
rect 15396 23254 15424 25094
rect 16684 24818 16712 25910
rect 16672 24812 16724 24818
rect 16672 24754 16724 24760
rect 16776 24449 16804 26574
rect 17040 26512 17092 26518
rect 17040 26454 17092 26460
rect 17052 26382 17080 26454
rect 17040 26376 17092 26382
rect 17040 26318 17092 26324
rect 17052 25906 17080 26318
rect 17144 25974 17172 27406
rect 17316 26512 17368 26518
rect 17316 26454 17368 26460
rect 17328 26314 17356 26454
rect 17316 26308 17368 26314
rect 17316 26250 17368 26256
rect 17132 25968 17184 25974
rect 17132 25910 17184 25916
rect 17040 25900 17092 25906
rect 17040 25842 17092 25848
rect 16856 25696 16908 25702
rect 16856 25638 16908 25644
rect 16762 24440 16818 24449
rect 16762 24375 16818 24384
rect 16868 24206 16896 25638
rect 17144 25498 17172 25910
rect 17132 25492 17184 25498
rect 17132 25434 17184 25440
rect 17224 25492 17276 25498
rect 17224 25434 17276 25440
rect 17144 25242 17172 25434
rect 17052 25214 17172 25242
rect 16948 24812 17000 24818
rect 16948 24754 17000 24760
rect 16960 24410 16988 24754
rect 16948 24404 17000 24410
rect 16948 24346 17000 24352
rect 16856 24200 16908 24206
rect 16856 24142 16908 24148
rect 17052 23866 17080 25214
rect 17132 24200 17184 24206
rect 17236 24188 17264 25434
rect 17316 25288 17368 25294
rect 17316 25230 17368 25236
rect 17328 24818 17356 25230
rect 17420 24886 17448 29038
rect 17498 27976 17554 27985
rect 17498 27911 17500 27920
rect 17552 27911 17554 27920
rect 17500 27882 17552 27888
rect 17512 26994 17540 27882
rect 17500 26988 17552 26994
rect 17500 26930 17552 26936
rect 17500 26308 17552 26314
rect 17500 26250 17552 26256
rect 17512 26042 17540 26250
rect 17500 26036 17552 26042
rect 17500 25978 17552 25984
rect 17408 24880 17460 24886
rect 17408 24822 17460 24828
rect 17316 24812 17368 24818
rect 17316 24754 17368 24760
rect 17604 24342 17632 32710
rect 17696 32230 17724 35430
rect 17684 32224 17736 32230
rect 17684 32166 17736 32172
rect 17696 31890 17724 32166
rect 17684 31884 17736 31890
rect 17684 31826 17736 31832
rect 17788 31278 17816 37266
rect 30944 37262 30972 37402
rect 30932 37256 30984 37262
rect 30932 37198 30984 37204
rect 31024 37120 31076 37126
rect 31024 37062 31076 37068
rect 19574 37020 19882 37029
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36955 19882 36964
rect 19574 35932 19882 35941
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35867 19882 35876
rect 18788 35556 18840 35562
rect 18788 35498 18840 35504
rect 18144 33516 18196 33522
rect 18144 33458 18196 33464
rect 17960 33448 18012 33454
rect 17960 33390 18012 33396
rect 17972 31958 18000 33390
rect 17960 31952 18012 31958
rect 17960 31894 18012 31900
rect 18156 31890 18184 33458
rect 18236 32360 18288 32366
rect 18236 32302 18288 32308
rect 18144 31884 18196 31890
rect 18144 31826 18196 31832
rect 18248 31278 18276 32302
rect 18512 31680 18564 31686
rect 18512 31622 18564 31628
rect 18328 31408 18380 31414
rect 18328 31350 18380 31356
rect 17776 31272 17828 31278
rect 17776 31214 17828 31220
rect 18052 31272 18104 31278
rect 18052 31214 18104 31220
rect 18236 31272 18288 31278
rect 18236 31214 18288 31220
rect 17960 31136 18012 31142
rect 17960 31078 18012 31084
rect 17776 30728 17828 30734
rect 17776 30670 17828 30676
rect 17788 28014 17816 30670
rect 17972 30190 18000 31078
rect 18064 30666 18092 31214
rect 18052 30660 18104 30666
rect 18052 30602 18104 30608
rect 18340 30598 18368 31350
rect 18524 31278 18552 31622
rect 18512 31272 18564 31278
rect 18512 31214 18564 31220
rect 18512 30660 18564 30666
rect 18512 30602 18564 30608
rect 18328 30592 18380 30598
rect 18328 30534 18380 30540
rect 17960 30184 18012 30190
rect 17960 30126 18012 30132
rect 17972 28370 18000 30126
rect 18340 29782 18368 30534
rect 18328 29776 18380 29782
rect 18328 29718 18380 29724
rect 18524 29510 18552 30602
rect 18604 29708 18656 29714
rect 18604 29650 18656 29656
rect 18512 29504 18564 29510
rect 18512 29446 18564 29452
rect 18420 29164 18472 29170
rect 18420 29106 18472 29112
rect 17880 28342 18184 28370
rect 17880 28218 17908 28342
rect 17868 28212 17920 28218
rect 17868 28154 17920 28160
rect 18052 28212 18104 28218
rect 18052 28154 18104 28160
rect 17776 28008 17828 28014
rect 17776 27950 17828 27956
rect 17880 26874 17908 28154
rect 17960 28076 18012 28082
rect 17960 28018 18012 28024
rect 17972 27606 18000 28018
rect 18064 27674 18092 28154
rect 18156 28082 18184 28342
rect 18236 28212 18288 28218
rect 18236 28154 18288 28160
rect 18144 28076 18196 28082
rect 18144 28018 18196 28024
rect 18052 27668 18104 27674
rect 18052 27610 18104 27616
rect 17960 27600 18012 27606
rect 17960 27542 18012 27548
rect 18064 26994 18092 27610
rect 17960 26988 18012 26994
rect 17960 26930 18012 26936
rect 18052 26988 18104 26994
rect 18052 26930 18104 26936
rect 17696 26846 17908 26874
rect 17592 24336 17644 24342
rect 17592 24278 17644 24284
rect 17184 24160 17264 24188
rect 17132 24142 17184 24148
rect 17040 23860 17092 23866
rect 17040 23802 17092 23808
rect 15752 23724 15804 23730
rect 15752 23666 15804 23672
rect 16580 23724 16632 23730
rect 16580 23666 16632 23672
rect 15764 23526 15792 23666
rect 15752 23520 15804 23526
rect 15752 23462 15804 23468
rect 16210 23488 16266 23497
rect 15292 23248 15344 23254
rect 15292 23190 15344 23196
rect 15384 23248 15436 23254
rect 15384 23190 15436 23196
rect 15108 22976 15160 22982
rect 15108 22918 15160 22924
rect 15120 22778 15148 22918
rect 15108 22772 15160 22778
rect 15108 22714 15160 22720
rect 15396 22642 15424 23190
rect 14648 22636 14700 22642
rect 14648 22578 14700 22584
rect 15016 22636 15068 22642
rect 15016 22578 15068 22584
rect 15384 22636 15436 22642
rect 15384 22578 15436 22584
rect 15396 22438 15424 22578
rect 15384 22432 15436 22438
rect 15384 22374 15436 22380
rect 15764 2650 15792 23462
rect 16210 23423 16266 23432
rect 15844 23316 15896 23322
rect 15844 23258 15896 23264
rect 15856 23186 15884 23258
rect 15844 23180 15896 23186
rect 15844 23122 15896 23128
rect 15856 22642 15884 23122
rect 16224 23118 16252 23423
rect 16028 23112 16080 23118
rect 16028 23054 16080 23060
rect 16212 23112 16264 23118
rect 16592 23089 16620 23666
rect 17132 23656 17184 23662
rect 17132 23598 17184 23604
rect 16856 23520 16908 23526
rect 16856 23462 16908 23468
rect 16212 23054 16264 23060
rect 16578 23080 16634 23089
rect 15844 22636 15896 22642
rect 15844 22578 15896 22584
rect 16040 22574 16068 23054
rect 16224 22778 16252 23054
rect 16868 23050 16896 23462
rect 16948 23112 17000 23118
rect 16948 23054 17000 23060
rect 16578 23015 16580 23024
rect 16632 23015 16634 23024
rect 16856 23044 16908 23050
rect 16580 22986 16632 22992
rect 16856 22986 16908 22992
rect 16592 22955 16620 22986
rect 16672 22976 16724 22982
rect 16672 22918 16724 22924
rect 16212 22772 16264 22778
rect 16212 22714 16264 22720
rect 16028 22568 16080 22574
rect 16028 22510 16080 22516
rect 16684 22234 16712 22918
rect 16868 22710 16896 22986
rect 16960 22710 16988 23054
rect 17144 22778 17172 23598
rect 17604 23497 17632 24278
rect 17696 23730 17724 26846
rect 17776 26784 17828 26790
rect 17776 26726 17828 26732
rect 17684 23724 17736 23730
rect 17684 23666 17736 23672
rect 17590 23488 17646 23497
rect 17590 23423 17646 23432
rect 17408 23316 17460 23322
rect 17408 23258 17460 23264
rect 17316 23248 17368 23254
rect 17314 23216 17316 23225
rect 17368 23216 17370 23225
rect 17314 23151 17370 23160
rect 17420 22778 17448 23258
rect 17132 22772 17184 22778
rect 17132 22714 17184 22720
rect 17408 22772 17460 22778
rect 17408 22714 17460 22720
rect 16856 22704 16908 22710
rect 16856 22646 16908 22652
rect 16948 22704 17000 22710
rect 16948 22646 17000 22652
rect 17696 22658 17724 23666
rect 17788 23254 17816 26726
rect 17868 26580 17920 26586
rect 17868 26522 17920 26528
rect 17880 24410 17908 26522
rect 17972 26314 18000 26930
rect 18248 26858 18276 28154
rect 18432 27962 18460 29106
rect 18524 28422 18552 29446
rect 18616 28762 18644 29650
rect 18604 28756 18656 28762
rect 18604 28698 18656 28704
rect 18512 28416 18564 28422
rect 18512 28358 18564 28364
rect 18524 28218 18552 28358
rect 18512 28212 18564 28218
rect 18512 28154 18564 28160
rect 18616 28150 18644 28698
rect 18800 28490 18828 35498
rect 19574 34844 19882 34853
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34779 19882 34788
rect 18880 34740 18932 34746
rect 18880 34682 18932 34688
rect 18892 29170 18920 34682
rect 31036 33862 31064 37062
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 31024 33856 31076 33862
rect 31024 33798 31076 33804
rect 19574 33756 19882 33765
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33691 19882 33700
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 19574 32668 19882 32677
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32603 19882 32612
rect 21640 32224 21692 32230
rect 21640 32166 21692 32172
rect 37832 32224 37884 32230
rect 37832 32166 37884 32172
rect 19432 32020 19484 32026
rect 19432 31962 19484 31968
rect 19444 31822 19472 31962
rect 19524 31952 19576 31958
rect 19524 31894 19576 31900
rect 19432 31816 19484 31822
rect 19432 31758 19484 31764
rect 19340 31748 19392 31754
rect 19340 31690 19392 31696
rect 19352 30433 19380 31690
rect 19444 31482 19472 31758
rect 19536 31754 19564 31894
rect 20260 31816 20312 31822
rect 20260 31758 20312 31764
rect 19524 31748 19576 31754
rect 19524 31690 19576 31696
rect 19574 31580 19882 31589
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31515 19882 31524
rect 19432 31476 19484 31482
rect 19432 31418 19484 31424
rect 20076 31272 20128 31278
rect 20272 31260 20300 31758
rect 20628 31680 20680 31686
rect 20628 31622 20680 31628
rect 20128 31232 20300 31260
rect 20076 31214 20128 31220
rect 20088 30666 20116 31214
rect 20640 31142 20668 31622
rect 20260 31136 20312 31142
rect 20260 31078 20312 31084
rect 20628 31136 20680 31142
rect 20628 31078 20680 31084
rect 20272 30666 20300 31078
rect 20444 30728 20496 30734
rect 20444 30670 20496 30676
rect 20076 30660 20128 30666
rect 20076 30602 20128 30608
rect 20260 30660 20312 30666
rect 20260 30602 20312 30608
rect 19574 30492 19882 30501
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19338 30424 19394 30433
rect 19574 30427 19882 30436
rect 19338 30359 19394 30368
rect 19340 30320 19392 30326
rect 19340 30262 19392 30268
rect 19432 30320 19484 30326
rect 19616 30320 19668 30326
rect 19432 30262 19484 30268
rect 19522 30288 19578 30297
rect 18972 30048 19024 30054
rect 18972 29990 19024 29996
rect 18880 29164 18932 29170
rect 18880 29106 18932 29112
rect 18880 29028 18932 29034
rect 18880 28970 18932 28976
rect 18788 28484 18840 28490
rect 18788 28426 18840 28432
rect 18696 28416 18748 28422
rect 18696 28358 18748 28364
rect 18604 28144 18656 28150
rect 18604 28086 18656 28092
rect 18432 27934 18644 27962
rect 18420 27872 18472 27878
rect 18420 27814 18472 27820
rect 18432 27402 18460 27814
rect 18420 27396 18472 27402
rect 18420 27338 18472 27344
rect 18236 26852 18288 26858
rect 18236 26794 18288 26800
rect 18616 26602 18644 27934
rect 18708 27614 18736 28358
rect 18800 27962 18828 28426
rect 18892 28082 18920 28970
rect 18880 28076 18932 28082
rect 18880 28018 18932 28024
rect 18800 27934 18920 27962
rect 18708 27586 18828 27614
rect 18800 26926 18828 27586
rect 18892 27334 18920 27934
rect 18880 27328 18932 27334
rect 18880 27270 18932 27276
rect 18892 27130 18920 27270
rect 18880 27124 18932 27130
rect 18880 27066 18932 27072
rect 18788 26920 18840 26926
rect 18788 26862 18840 26868
rect 18432 26574 18644 26602
rect 17960 26308 18012 26314
rect 17960 26250 18012 26256
rect 18328 26036 18380 26042
rect 18328 25978 18380 25984
rect 18052 25900 18104 25906
rect 18052 25842 18104 25848
rect 17960 25492 18012 25498
rect 17960 25434 18012 25440
rect 17868 24404 17920 24410
rect 17868 24346 17920 24352
rect 17972 23798 18000 25434
rect 18064 24954 18092 25842
rect 18236 25288 18288 25294
rect 18236 25230 18288 25236
rect 18052 24948 18104 24954
rect 18052 24890 18104 24896
rect 18144 24948 18196 24954
rect 18144 24890 18196 24896
rect 18156 24818 18184 24890
rect 18144 24812 18196 24818
rect 18144 24754 18196 24760
rect 18144 24132 18196 24138
rect 18144 24074 18196 24080
rect 17960 23792 18012 23798
rect 17960 23734 18012 23740
rect 17776 23248 17828 23254
rect 17776 23190 17828 23196
rect 17868 23248 17920 23254
rect 17868 23190 17920 23196
rect 17880 23066 17908 23190
rect 17972 23100 18000 23734
rect 17788 23038 17908 23066
rect 17956 23072 18000 23100
rect 18052 23112 18104 23118
rect 17788 22982 17816 23038
rect 17956 23032 17984 23072
rect 18156 23089 18184 24074
rect 18248 23610 18276 25230
rect 18340 23798 18368 25978
rect 18432 24274 18460 26574
rect 18512 26512 18564 26518
rect 18512 26454 18564 26460
rect 18420 24268 18472 24274
rect 18420 24210 18472 24216
rect 18420 24064 18472 24070
rect 18420 24006 18472 24012
rect 18432 23866 18460 24006
rect 18420 23860 18472 23866
rect 18420 23802 18472 23808
rect 18328 23792 18380 23798
rect 18328 23734 18380 23740
rect 18248 23582 18368 23610
rect 18052 23054 18104 23060
rect 18142 23080 18198 23089
rect 17956 23004 18000 23032
rect 17776 22976 17828 22982
rect 17776 22918 17828 22924
rect 17696 22630 17908 22658
rect 17972 22642 18000 23004
rect 18064 22778 18092 23054
rect 18142 23015 18144 23024
rect 18196 23015 18198 23024
rect 18144 22986 18196 22992
rect 18052 22772 18104 22778
rect 18052 22714 18104 22720
rect 17880 22574 17908 22630
rect 17960 22636 18012 22642
rect 17960 22578 18012 22584
rect 17868 22568 17920 22574
rect 17868 22510 17920 22516
rect 18156 22234 18184 22986
rect 18236 22636 18288 22642
rect 18236 22578 18288 22584
rect 18248 22438 18276 22578
rect 18236 22432 18288 22438
rect 18236 22374 18288 22380
rect 16672 22228 16724 22234
rect 16672 22170 16724 22176
rect 18144 22228 18196 22234
rect 18144 22170 18196 22176
rect 18236 22228 18288 22234
rect 18236 22170 18288 22176
rect 18248 21690 18276 22170
rect 18340 21894 18368 23582
rect 18328 21888 18380 21894
rect 18328 21830 18380 21836
rect 18236 21684 18288 21690
rect 18236 21626 18288 21632
rect 18524 12850 18552 26454
rect 18800 26382 18828 26862
rect 18892 26586 18920 27066
rect 18880 26580 18932 26586
rect 18880 26522 18932 26528
rect 18788 26376 18840 26382
rect 18788 26318 18840 26324
rect 18604 25288 18656 25294
rect 18604 25230 18656 25236
rect 18616 23866 18644 25230
rect 18696 25152 18748 25158
rect 18696 25094 18748 25100
rect 18604 23860 18656 23866
rect 18604 23802 18656 23808
rect 18708 21078 18736 25094
rect 18800 23186 18828 26318
rect 18880 24268 18932 24274
rect 18880 24210 18932 24216
rect 18788 23180 18840 23186
rect 18788 23122 18840 23128
rect 18788 22976 18840 22982
rect 18788 22918 18840 22924
rect 18800 22642 18828 22918
rect 18788 22636 18840 22642
rect 18788 22578 18840 22584
rect 18892 22574 18920 24210
rect 18984 23050 19012 29990
rect 19064 29504 19116 29510
rect 19064 29446 19116 29452
rect 19076 29102 19104 29446
rect 19248 29232 19300 29238
rect 19248 29174 19300 29180
rect 19064 29096 19116 29102
rect 19064 29038 19116 29044
rect 19156 29028 19208 29034
rect 19156 28970 19208 28976
rect 19064 27940 19116 27946
rect 19064 27882 19116 27888
rect 19076 27130 19104 27882
rect 19064 27124 19116 27130
rect 19064 27066 19116 27072
rect 19076 26790 19104 27066
rect 19064 26784 19116 26790
rect 19064 26726 19116 26732
rect 19064 26580 19116 26586
rect 19064 26522 19116 26528
rect 19076 26364 19104 26522
rect 19168 26489 19196 28970
rect 19260 28490 19288 29174
rect 19352 28762 19380 30262
rect 19444 29714 19472 30262
rect 19616 30262 19668 30268
rect 19984 30320 20036 30326
rect 19984 30262 20036 30268
rect 19522 30223 19578 30232
rect 19432 29708 19484 29714
rect 19432 29650 19484 29656
rect 19536 29492 19564 30223
rect 19628 30122 19656 30262
rect 19616 30116 19668 30122
rect 19616 30058 19668 30064
rect 19800 30048 19852 30054
rect 19800 29990 19852 29996
rect 19812 29510 19840 29990
rect 19444 29464 19564 29492
rect 19800 29504 19852 29510
rect 19444 29034 19472 29464
rect 19800 29446 19852 29452
rect 19574 29404 19882 29413
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29339 19882 29348
rect 19432 29028 19484 29034
rect 19432 28970 19484 28976
rect 19340 28756 19392 28762
rect 19340 28698 19392 28704
rect 19444 28642 19472 28970
rect 19352 28614 19472 28642
rect 19248 28484 19300 28490
rect 19248 28426 19300 28432
rect 19352 27538 19380 28614
rect 19432 28552 19484 28558
rect 19432 28494 19484 28500
rect 19444 27826 19472 28494
rect 19574 28316 19882 28325
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28251 19882 28260
rect 19892 27872 19944 27878
rect 19444 27798 19564 27826
rect 19892 27814 19944 27820
rect 19432 27668 19484 27674
rect 19432 27610 19484 27616
rect 19340 27532 19392 27538
rect 19340 27474 19392 27480
rect 19248 27328 19300 27334
rect 19248 27270 19300 27276
rect 19260 26926 19288 27270
rect 19444 27130 19472 27610
rect 19536 27334 19564 27798
rect 19904 27470 19932 27814
rect 19892 27464 19944 27470
rect 19706 27432 19762 27441
rect 19892 27406 19944 27412
rect 19706 27367 19708 27376
rect 19760 27367 19762 27376
rect 19708 27338 19760 27344
rect 19524 27328 19576 27334
rect 19524 27270 19576 27276
rect 19574 27228 19882 27237
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27163 19882 27172
rect 19432 27124 19484 27130
rect 19432 27066 19484 27072
rect 19708 27124 19760 27130
rect 19708 27066 19760 27072
rect 19524 27056 19576 27062
rect 19522 27024 19524 27033
rect 19576 27024 19578 27033
rect 19432 26988 19484 26994
rect 19522 26959 19578 26968
rect 19432 26930 19484 26936
rect 19248 26920 19300 26926
rect 19248 26862 19300 26868
rect 19260 26518 19288 26862
rect 19444 26761 19472 26930
rect 19616 26920 19668 26926
rect 19616 26862 19668 26868
rect 19524 26784 19576 26790
rect 19430 26752 19486 26761
rect 19524 26726 19576 26732
rect 19430 26687 19486 26696
rect 19248 26512 19300 26518
rect 19154 26480 19210 26489
rect 19248 26454 19300 26460
rect 19154 26415 19210 26424
rect 19076 26336 19196 26364
rect 19168 25974 19196 26336
rect 19156 25968 19208 25974
rect 19156 25910 19208 25916
rect 19064 24608 19116 24614
rect 19064 24550 19116 24556
rect 19076 23798 19104 24550
rect 19168 24070 19196 25910
rect 19156 24064 19208 24070
rect 19156 24006 19208 24012
rect 19064 23792 19116 23798
rect 19064 23734 19116 23740
rect 19076 23118 19104 23734
rect 19260 23526 19288 26454
rect 19340 26444 19392 26450
rect 19340 26386 19392 26392
rect 19352 26353 19380 26386
rect 19338 26344 19394 26353
rect 19338 26279 19394 26288
rect 19536 26228 19564 26726
rect 19628 26586 19656 26862
rect 19720 26858 19748 27066
rect 19890 26888 19946 26897
rect 19708 26852 19760 26858
rect 19890 26823 19946 26832
rect 19708 26794 19760 26800
rect 19616 26580 19668 26586
rect 19616 26522 19668 26528
rect 19444 26200 19564 26228
rect 19904 26228 19932 26823
rect 19996 26586 20024 30262
rect 20088 30258 20116 30602
rect 20076 30252 20128 30258
rect 20076 30194 20128 30200
rect 20088 29646 20116 30194
rect 20272 30190 20300 30602
rect 20456 30326 20484 30670
rect 20444 30320 20496 30326
rect 20444 30262 20496 30268
rect 20260 30184 20312 30190
rect 20260 30126 20312 30132
rect 20076 29640 20128 29646
rect 20076 29582 20128 29588
rect 20260 29640 20312 29646
rect 20260 29582 20312 29588
rect 20076 29300 20128 29306
rect 20076 29242 20128 29248
rect 20088 26874 20116 29242
rect 20272 27946 20300 29582
rect 20444 29504 20496 29510
rect 20444 29446 20496 29452
rect 20456 28422 20484 29446
rect 21180 29164 21232 29170
rect 21180 29106 21232 29112
rect 20536 28960 20588 28966
rect 20536 28902 20588 28908
rect 20444 28416 20496 28422
rect 20444 28358 20496 28364
rect 20456 28014 20484 28358
rect 20548 28150 20576 28902
rect 20536 28144 20588 28150
rect 20536 28086 20588 28092
rect 20444 28008 20496 28014
rect 20444 27950 20496 27956
rect 20260 27940 20312 27946
rect 20260 27882 20312 27888
rect 20088 26846 20208 26874
rect 20076 26784 20128 26790
rect 20074 26752 20076 26761
rect 20128 26752 20130 26761
rect 20074 26687 20130 26696
rect 19984 26580 20036 26586
rect 19984 26522 20036 26528
rect 19904 26200 20024 26228
rect 19444 25498 19472 26200
rect 19574 26140 19882 26149
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26075 19882 26084
rect 19432 25492 19484 25498
rect 19996 25480 20024 26200
rect 20180 25702 20208 26846
rect 20168 25696 20220 25702
rect 20168 25638 20220 25644
rect 19432 25434 19484 25440
rect 19812 25452 20024 25480
rect 19444 25294 19472 25434
rect 19812 25362 19840 25452
rect 20272 25378 20300 27882
rect 20350 26344 20406 26353
rect 20350 26279 20406 26288
rect 20364 25770 20392 26279
rect 20352 25764 20404 25770
rect 20352 25706 20404 25712
rect 19800 25356 19852 25362
rect 19800 25298 19852 25304
rect 19996 25350 20300 25378
rect 19432 25288 19484 25294
rect 19432 25230 19484 25236
rect 19706 25256 19762 25265
rect 19706 25191 19762 25200
rect 19720 25158 19748 25191
rect 19812 25158 19840 25298
rect 19432 25152 19484 25158
rect 19432 25094 19484 25100
rect 19708 25152 19760 25158
rect 19708 25094 19760 25100
rect 19800 25152 19852 25158
rect 19800 25094 19852 25100
rect 19444 24993 19472 25094
rect 19574 25052 19882 25061
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19430 24984 19486 24993
rect 19574 24987 19882 24996
rect 19430 24919 19486 24928
rect 19892 24880 19944 24886
rect 19352 24818 19656 24834
rect 19892 24822 19944 24828
rect 19340 24812 19656 24818
rect 19392 24806 19656 24812
rect 19340 24754 19392 24760
rect 19524 24744 19576 24750
rect 19338 24712 19394 24721
rect 19524 24686 19576 24692
rect 19338 24647 19394 24656
rect 19352 24410 19380 24647
rect 19340 24404 19392 24410
rect 19340 24346 19392 24352
rect 19536 24206 19564 24686
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 19628 24070 19656 24806
rect 19432 24064 19484 24070
rect 19432 24006 19484 24012
rect 19616 24064 19668 24070
rect 19904 24052 19932 24822
rect 19996 24290 20024 25350
rect 20258 25256 20314 25265
rect 20168 25220 20220 25226
rect 20258 25191 20260 25200
rect 20168 25162 20220 25168
rect 20312 25191 20314 25200
rect 20260 25162 20312 25168
rect 20180 24886 20208 25162
rect 20168 24880 20220 24886
rect 20168 24822 20220 24828
rect 20364 24818 20392 25706
rect 20076 24812 20128 24818
rect 20076 24754 20128 24760
rect 20352 24812 20404 24818
rect 20352 24754 20404 24760
rect 20088 24410 20116 24754
rect 20076 24404 20128 24410
rect 20076 24346 20128 24352
rect 19996 24262 20208 24290
rect 19904 24024 20024 24052
rect 19616 24006 19668 24012
rect 19248 23520 19300 23526
rect 19248 23462 19300 23468
rect 19444 23322 19472 24006
rect 19574 23964 19882 23973
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23899 19882 23908
rect 19432 23316 19484 23322
rect 19432 23258 19484 23264
rect 19064 23112 19116 23118
rect 19064 23054 19116 23060
rect 18972 23044 19024 23050
rect 18972 22986 19024 22992
rect 18984 22710 19012 22986
rect 19076 22710 19104 23054
rect 19524 22976 19576 22982
rect 19444 22936 19524 22964
rect 18972 22704 19024 22710
rect 18972 22646 19024 22652
rect 19064 22704 19116 22710
rect 19064 22646 19116 22652
rect 18880 22568 18932 22574
rect 18880 22510 18932 22516
rect 18892 21690 18920 22510
rect 19076 22506 19104 22646
rect 19064 22500 19116 22506
rect 19064 22442 19116 22448
rect 19076 22386 19104 22442
rect 18984 22358 19104 22386
rect 18984 22234 19012 22358
rect 18972 22228 19024 22234
rect 18972 22170 19024 22176
rect 19064 22228 19116 22234
rect 19064 22170 19116 22176
rect 18880 21684 18932 21690
rect 18880 21626 18932 21632
rect 18696 21072 18748 21078
rect 18696 21014 18748 21020
rect 19076 21010 19104 22170
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 19260 21842 19288 21966
rect 19260 21814 19380 21842
rect 19064 21004 19116 21010
rect 19064 20946 19116 20952
rect 19076 20602 19104 20946
rect 19352 20942 19380 21814
rect 19444 21554 19472 22936
rect 19524 22918 19576 22924
rect 19574 22876 19882 22885
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22811 19882 22820
rect 19996 22556 20024 24024
rect 19904 22528 20024 22556
rect 19904 22030 19932 22528
rect 20076 22500 20128 22506
rect 20076 22442 20128 22448
rect 19984 22432 20036 22438
rect 19984 22374 20036 22380
rect 19892 22024 19944 22030
rect 19892 21966 19944 21972
rect 19574 21788 19882 21797
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21723 19882 21732
rect 19996 21690 20024 22374
rect 19984 21684 20036 21690
rect 19984 21626 20036 21632
rect 20088 21554 20116 22442
rect 20180 21962 20208 24262
rect 20260 23248 20312 23254
rect 20260 23190 20312 23196
rect 20272 22438 20300 23190
rect 20260 22432 20312 22438
rect 20260 22374 20312 22380
rect 20364 22234 20392 24754
rect 20352 22228 20404 22234
rect 20352 22170 20404 22176
rect 20168 21956 20220 21962
rect 20168 21898 20220 21904
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 20076 21548 20128 21554
rect 20076 21490 20128 21496
rect 20456 21486 20484 27950
rect 20548 27606 20576 28086
rect 20536 27600 20588 27606
rect 20536 27542 20588 27548
rect 20548 26858 20576 27542
rect 20628 27396 20680 27402
rect 20628 27338 20680 27344
rect 20640 27130 20668 27338
rect 21088 27328 21140 27334
rect 21088 27270 21140 27276
rect 20628 27124 20680 27130
rect 20628 27066 20680 27072
rect 20536 26852 20588 26858
rect 20536 26794 20588 26800
rect 20536 26580 20588 26586
rect 20536 26522 20588 26528
rect 20548 25294 20576 26522
rect 20640 25294 20668 27066
rect 20812 27056 20864 27062
rect 20810 27024 20812 27033
rect 20996 27056 21048 27062
rect 20864 27024 20866 27033
rect 20996 26998 21048 27004
rect 20810 26959 20866 26968
rect 20720 26920 20772 26926
rect 20720 26862 20772 26868
rect 20732 25430 20760 26862
rect 21008 26858 21036 26998
rect 20812 26852 20864 26858
rect 20812 26794 20864 26800
rect 20996 26852 21048 26858
rect 20996 26794 21048 26800
rect 20824 26042 20852 26794
rect 21100 26518 21128 27270
rect 21088 26512 21140 26518
rect 21088 26454 21140 26460
rect 20812 26036 20864 26042
rect 20864 25996 20944 26024
rect 20812 25978 20864 25984
rect 20812 25696 20864 25702
rect 20812 25638 20864 25644
rect 20720 25424 20772 25430
rect 20720 25366 20772 25372
rect 20732 25294 20760 25366
rect 20536 25288 20588 25294
rect 20536 25230 20588 25236
rect 20628 25288 20680 25294
rect 20628 25230 20680 25236
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 20824 25106 20852 25638
rect 20640 25078 20852 25106
rect 20536 23112 20588 23118
rect 20536 23054 20588 23060
rect 20548 22778 20576 23054
rect 20536 22772 20588 22778
rect 20536 22714 20588 22720
rect 20640 22094 20668 25078
rect 20916 24342 20944 25996
rect 20996 25900 21048 25906
rect 20996 25842 21048 25848
rect 20904 24336 20956 24342
rect 20904 24278 20956 24284
rect 20812 24132 20864 24138
rect 20812 24074 20864 24080
rect 20720 23656 20772 23662
rect 20720 23598 20772 23604
rect 20732 23322 20760 23598
rect 20720 23316 20772 23322
rect 20720 23258 20772 23264
rect 20720 22772 20772 22778
rect 20720 22714 20772 22720
rect 20548 22066 20668 22094
rect 20548 22030 20576 22066
rect 20536 22024 20588 22030
rect 20536 21966 20588 21972
rect 20548 21622 20576 21966
rect 20536 21616 20588 21622
rect 20536 21558 20588 21564
rect 20444 21480 20496 21486
rect 20444 21422 20496 21428
rect 20548 20942 20576 21558
rect 20732 21554 20760 22714
rect 20824 22574 20852 24074
rect 20916 23866 20944 24278
rect 21008 24206 21036 25842
rect 21192 24886 21220 29106
rect 21652 27606 21680 32166
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 37844 30802 37872 32166
rect 37832 30796 37884 30802
rect 37832 30738 37884 30744
rect 38108 30728 38160 30734
rect 38106 30696 38108 30705
rect 38160 30696 38162 30705
rect 38106 30631 38162 30640
rect 38120 30394 38148 30631
rect 38108 30388 38160 30394
rect 38108 30330 38160 30336
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 23662 28928 23718 28937
rect 23662 28863 23718 28872
rect 21640 27600 21692 27606
rect 21640 27542 21692 27548
rect 21652 26926 21680 27542
rect 22100 27464 22152 27470
rect 22100 27406 22152 27412
rect 22112 26994 22140 27406
rect 22652 27056 22704 27062
rect 22652 26998 22704 27004
rect 22100 26988 22152 26994
rect 22020 26948 22100 26976
rect 21640 26920 21692 26926
rect 21692 26868 21772 26874
rect 21640 26862 21772 26868
rect 21652 26846 21772 26862
rect 21364 26784 21416 26790
rect 21364 26726 21416 26732
rect 21640 26784 21692 26790
rect 21640 26726 21692 26732
rect 21272 26444 21324 26450
rect 21272 26386 21324 26392
rect 21180 24880 21232 24886
rect 21180 24822 21232 24828
rect 20996 24200 21048 24206
rect 20996 24142 21048 24148
rect 20904 23860 20956 23866
rect 20904 23802 20956 23808
rect 21008 23798 21036 24142
rect 20996 23792 21048 23798
rect 20996 23734 21048 23740
rect 21008 23118 21036 23734
rect 20996 23112 21048 23118
rect 20996 23054 21048 23060
rect 21192 22710 21220 24822
rect 21180 22704 21232 22710
rect 21180 22646 21232 22652
rect 21284 22642 21312 26386
rect 21376 26382 21404 26726
rect 21652 26382 21680 26726
rect 21364 26376 21416 26382
rect 21364 26318 21416 26324
rect 21640 26376 21692 26382
rect 21640 26318 21692 26324
rect 21744 25702 21772 26846
rect 22020 26246 22048 26948
rect 22100 26930 22152 26936
rect 22664 26382 22692 26998
rect 22100 26376 22152 26382
rect 22100 26318 22152 26324
rect 22652 26376 22704 26382
rect 22652 26318 22704 26324
rect 22008 26240 22060 26246
rect 22008 26182 22060 26188
rect 22020 25906 22048 26182
rect 22112 26042 22140 26318
rect 22100 26036 22152 26042
rect 22100 25978 22152 25984
rect 22008 25900 22060 25906
rect 22008 25842 22060 25848
rect 22100 25900 22152 25906
rect 22100 25842 22152 25848
rect 21732 25696 21784 25702
rect 21732 25638 21784 25644
rect 21744 25498 21772 25638
rect 21732 25492 21784 25498
rect 21732 25434 21784 25440
rect 21744 24750 21772 25434
rect 22112 25430 22140 25842
rect 22100 25424 22152 25430
rect 22100 25366 22152 25372
rect 23676 24818 23704 28863
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 21916 24812 21968 24818
rect 21916 24754 21968 24760
rect 23664 24812 23716 24818
rect 23664 24754 23716 24760
rect 23940 24812 23992 24818
rect 23940 24754 23992 24760
rect 24400 24812 24452 24818
rect 24400 24754 24452 24760
rect 21732 24744 21784 24750
rect 21732 24686 21784 24692
rect 21744 24410 21772 24686
rect 21732 24404 21784 24410
rect 21732 24346 21784 24352
rect 21744 23730 21772 24346
rect 21928 23866 21956 24754
rect 22008 24608 22060 24614
rect 22008 24550 22060 24556
rect 23388 24608 23440 24614
rect 23388 24550 23440 24556
rect 22020 24342 22048 24550
rect 22008 24336 22060 24342
rect 22008 24278 22060 24284
rect 22376 24336 22428 24342
rect 22376 24278 22428 24284
rect 21916 23860 21968 23866
rect 21916 23802 21968 23808
rect 21732 23724 21784 23730
rect 21732 23666 21784 23672
rect 21744 23254 21772 23666
rect 22020 23594 22048 24278
rect 22192 23792 22244 23798
rect 22192 23734 22244 23740
rect 22008 23588 22060 23594
rect 22008 23530 22060 23536
rect 21732 23248 21784 23254
rect 21732 23190 21784 23196
rect 21744 23118 21772 23190
rect 21732 23112 21784 23118
rect 21732 23054 21784 23060
rect 21744 22642 21772 23054
rect 22204 22642 22232 23734
rect 22284 23724 22336 23730
rect 22284 23666 22336 23672
rect 22296 23322 22324 23666
rect 22284 23316 22336 23322
rect 22284 23258 22336 23264
rect 22388 23254 22416 24278
rect 23400 24274 23428 24550
rect 23480 24336 23532 24342
rect 23480 24278 23532 24284
rect 23388 24268 23440 24274
rect 23388 24210 23440 24216
rect 23204 24132 23256 24138
rect 23204 24074 23256 24080
rect 22742 23760 22798 23769
rect 23216 23730 23244 24074
rect 23400 23730 23428 24210
rect 22742 23695 22798 23704
rect 23204 23724 23256 23730
rect 22376 23248 22428 23254
rect 22376 23190 22428 23196
rect 22756 23186 22784 23695
rect 23204 23666 23256 23672
rect 23388 23724 23440 23730
rect 23388 23666 23440 23672
rect 23112 23520 23164 23526
rect 23112 23462 23164 23468
rect 22744 23180 22796 23186
rect 22744 23122 22796 23128
rect 22756 22778 22784 23122
rect 22744 22772 22796 22778
rect 22744 22714 22796 22720
rect 21272 22636 21324 22642
rect 21272 22578 21324 22584
rect 21732 22636 21784 22642
rect 21732 22578 21784 22584
rect 22008 22636 22060 22642
rect 22008 22578 22060 22584
rect 22192 22636 22244 22642
rect 22192 22578 22244 22584
rect 20812 22568 20864 22574
rect 20812 22510 20864 22516
rect 20904 22432 20956 22438
rect 20904 22374 20956 22380
rect 20812 22160 20864 22166
rect 20812 22102 20864 22108
rect 20824 21690 20852 22102
rect 20916 22030 20944 22374
rect 20904 22024 20956 22030
rect 20904 21966 20956 21972
rect 21284 21962 21312 22578
rect 21744 22506 21772 22578
rect 21732 22500 21784 22506
rect 21732 22442 21784 22448
rect 22020 22030 22048 22578
rect 22652 22160 22704 22166
rect 22652 22102 22704 22108
rect 22664 22030 22692 22102
rect 23124 22030 23152 23462
rect 23216 23322 23244 23666
rect 23492 23594 23520 24278
rect 23572 24200 23624 24206
rect 23572 24142 23624 24148
rect 23584 23730 23612 24142
rect 23952 23798 23980 24754
rect 24412 24410 24440 24754
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 24400 24404 24452 24410
rect 24400 24346 24452 24352
rect 24308 24064 24360 24070
rect 24308 24006 24360 24012
rect 23940 23792 23992 23798
rect 23940 23734 23992 23740
rect 24320 23730 24348 24006
rect 23572 23724 23624 23730
rect 23572 23666 23624 23672
rect 24308 23724 24360 23730
rect 24308 23666 24360 23672
rect 23480 23588 23532 23594
rect 23480 23530 23532 23536
rect 24584 23520 24636 23526
rect 24584 23462 24636 23468
rect 23204 23316 23256 23322
rect 23204 23258 23256 23264
rect 24596 23118 24624 23462
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 24584 23112 24636 23118
rect 24584 23054 24636 23060
rect 23296 22432 23348 22438
rect 23296 22374 23348 22380
rect 23308 22166 23336 22374
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 23296 22160 23348 22166
rect 23296 22102 23348 22108
rect 21548 22024 21600 22030
rect 21548 21966 21600 21972
rect 22008 22024 22060 22030
rect 22008 21966 22060 21972
rect 22652 22024 22704 22030
rect 22652 21966 22704 21972
rect 23112 22024 23164 22030
rect 23112 21966 23164 21972
rect 21272 21956 21324 21962
rect 21272 21898 21324 21904
rect 20812 21684 20864 21690
rect 20812 21626 20864 21632
rect 21560 21554 21588 21966
rect 22664 21554 22692 21966
rect 23124 21554 23152 21966
rect 23308 21690 23336 22102
rect 23296 21684 23348 21690
rect 23296 21626 23348 21632
rect 20720 21548 20772 21554
rect 20720 21490 20772 21496
rect 21088 21548 21140 21554
rect 21088 21490 21140 21496
rect 21180 21548 21232 21554
rect 21180 21490 21232 21496
rect 21548 21548 21600 21554
rect 21548 21490 21600 21496
rect 22284 21548 22336 21554
rect 22284 21490 22336 21496
rect 22652 21548 22704 21554
rect 22652 21490 22704 21496
rect 23112 21548 23164 21554
rect 23112 21490 23164 21496
rect 21100 21418 21128 21490
rect 21088 21412 21140 21418
rect 21088 21354 21140 21360
rect 21100 21010 21128 21354
rect 21192 21078 21220 21490
rect 21560 21146 21588 21490
rect 22192 21480 22244 21486
rect 22192 21422 22244 21428
rect 22204 21146 22232 21422
rect 21548 21140 21600 21146
rect 21548 21082 21600 21088
rect 22192 21140 22244 21146
rect 22192 21082 22244 21088
rect 21180 21072 21232 21078
rect 21180 21014 21232 21020
rect 21088 21004 21140 21010
rect 21088 20946 21140 20952
rect 19340 20936 19392 20942
rect 19340 20878 19392 20884
rect 20536 20936 20588 20942
rect 20536 20878 20588 20884
rect 19574 20700 19882 20709
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20635 19882 20644
rect 20548 20602 20576 20878
rect 21192 20602 21220 21014
rect 22296 20942 22324 21490
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 22284 20936 22336 20942
rect 22284 20878 22336 20884
rect 22296 20602 22324 20878
rect 19064 20596 19116 20602
rect 19064 20538 19116 20544
rect 20536 20596 20588 20602
rect 20536 20538 20588 20544
rect 21180 20596 21232 20602
rect 21180 20538 21232 20544
rect 22284 20596 22336 20602
rect 22284 20538 22336 20544
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 19574 19612 19882 19621
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19547 19882 19556
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 19574 18524 19882 18533
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18459 19882 18468
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 19574 17436 19882 17445
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17371 19882 17380
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 19574 16348 19882 16357
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16283 19882 16292
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 19574 15260 19882 15269
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15195 19882 15204
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 19574 14172 19882 14181
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14107 19882 14116
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 19574 13084 19882 13093
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13019 19882 13028
rect 18512 12844 18564 12850
rect 18512 12786 18564 12792
rect 37924 12640 37976 12646
rect 37924 12582 37976 12588
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 37936 12238 37964 12582
rect 38108 12368 38160 12374
rect 38106 12336 38108 12345
rect 38160 12336 38162 12345
rect 38106 12271 38162 12280
rect 37924 12232 37976 12238
rect 37924 12174 37976 12180
rect 19574 11996 19882 12005
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11931 19882 11940
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 19574 10908 19882 10917
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10843 19882 10852
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 19574 9820 19882 9829
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9755 19882 9764
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 19574 8732 19882 8741
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8667 19882 8676
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 19574 7644 19882 7653
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7579 19882 7588
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 19574 6556 19882 6565
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6491 19882 6500
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 19574 5468 19882 5477
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5403 19882 5412
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 19574 4380 19882 4389
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4315 19882 4324
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 19574 3292 19882 3301
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3227 19882 3236
rect 34520 2848 34572 2854
rect 34520 2790 34572 2796
rect 15752 2644 15804 2650
rect 15752 2586 15804 2592
rect 1400 2508 1452 2514
rect 1400 2450 1452 2456
rect 1676 2508 1728 2514
rect 1676 2450 1728 2456
rect 11336 2508 11388 2514
rect 11336 2450 11388 2456
rect 16764 2440 16816 2446
rect 16764 2382 16816 2388
rect 16776 800 16804 2382
rect 34532 2378 34560 2790
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 34520 2372 34572 2378
rect 34520 2314 34572 2320
rect 34532 2258 34560 2314
rect 34440 2230 34560 2258
rect 19574 2204 19882 2213
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2139 19882 2148
rect 34164 870 34284 898
rect 34164 800 34192 870
rect 18 0 74 800
rect 16762 0 16818 800
rect 34150 0 34206 800
rect 34256 762 34284 870
rect 34440 762 34468 2230
rect 34256 734 34468 762
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 3422 36080 3478 36136
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 1398 17720 1454 17776
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 2778 27920 2834 27976
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4066 27376 4122 27432
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4066 26444 4122 26480
rect 4066 26424 4068 26444
rect 4068 26424 4120 26444
rect 4120 26424 4122 26444
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 11702 29164 11758 29200
rect 11702 29144 11704 29164
rect 11704 29144 11756 29164
rect 11756 29144 11758 29164
rect 13634 28872 13690 28928
rect 13542 24404 13598 24440
rect 13542 24384 13544 24404
rect 13544 24384 13596 24404
rect 13596 24384 13598 24404
rect 13818 23740 13820 23760
rect 13820 23740 13872 23760
rect 13872 23740 13874 23760
rect 13818 23704 13874 23740
rect 14738 23704 14794 23760
rect 14646 23160 14702 23216
rect 17406 29144 17462 29200
rect 17222 28872 17278 28928
rect 16762 24384 16818 24440
rect 17498 27940 17554 27976
rect 17498 27920 17500 27940
rect 17500 27920 17552 27940
rect 17552 27920 17554 27940
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 16210 23432 16266 23488
rect 16578 23044 16634 23080
rect 16578 23024 16580 23044
rect 16580 23024 16632 23044
rect 16632 23024 16634 23044
rect 17590 23432 17646 23488
rect 17314 23196 17316 23216
rect 17316 23196 17368 23216
rect 17368 23196 17370 23216
rect 17314 23160 17370 23196
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19338 30368 19394 30424
rect 18142 23044 18198 23080
rect 18142 23024 18144 23044
rect 18144 23024 18196 23044
rect 18196 23024 18198 23044
rect 19522 30232 19578 30288
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19706 27396 19762 27432
rect 19706 27376 19708 27396
rect 19708 27376 19760 27396
rect 19760 27376 19762 27396
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19522 27004 19524 27024
rect 19524 27004 19576 27024
rect 19576 27004 19578 27024
rect 19522 26968 19578 27004
rect 19430 26696 19486 26752
rect 19154 26424 19210 26480
rect 19338 26288 19394 26344
rect 19890 26832 19946 26888
rect 20074 26732 20076 26752
rect 20076 26732 20128 26752
rect 20128 26732 20130 26752
rect 20074 26696 20130 26732
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 20350 26288 20406 26344
rect 19706 25200 19762 25256
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 19430 24928 19486 24984
rect 19338 24656 19394 24712
rect 20258 25220 20314 25256
rect 20258 25200 20260 25220
rect 20260 25200 20312 25220
rect 20312 25200 20314 25220
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 20810 27004 20812 27024
rect 20812 27004 20864 27024
rect 20864 27004 20866 27024
rect 20810 26968 20866 27004
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 38106 30676 38108 30696
rect 38108 30676 38160 30696
rect 38160 30676 38162 30696
rect 38106 30640 38162 30676
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 23662 28872 23718 28928
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 22742 23704 22798 23760
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 38106 12316 38108 12336
rect 38108 12316 38160 12336
rect 38160 12316 38162 12336
rect 38106 12280 38162 12316
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
<< metal3 >>
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 19570 37024 19886 37025
rect 19570 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19886 37024
rect 19570 36959 19886 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 0 36138 800 36168
rect 3417 36138 3483 36141
rect 0 36136 3483 36138
rect 0 36080 3422 36136
rect 3478 36080 3483 36136
rect 0 36078 3483 36080
rect 0 36048 800 36078
rect 3417 36075 3483 36078
rect 19570 35936 19886 35937
rect 19570 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19886 35936
rect 19570 35871 19886 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 19570 34848 19886 34849
rect 19570 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19886 34848
rect 19570 34783 19886 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19570 33760 19886 33761
rect 19570 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19886 33760
rect 19570 33695 19886 33696
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 19570 32672 19886 32673
rect 19570 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19886 32672
rect 19570 32607 19886 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 19570 31584 19886 31585
rect 19570 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19886 31584
rect 19570 31519 19886 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 38101 30698 38167 30701
rect 39200 30698 40000 30728
rect 38101 30696 40000 30698
rect 38101 30640 38106 30696
rect 38162 30640 40000 30696
rect 38101 30638 40000 30640
rect 38101 30635 38167 30638
rect 39200 30608 40000 30638
rect 19570 30496 19886 30497
rect 19570 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19886 30496
rect 19570 30431 19886 30432
rect 19333 30426 19399 30429
rect 19333 30424 19442 30426
rect 19333 30368 19338 30424
rect 19394 30368 19442 30424
rect 19333 30363 19442 30368
rect 19382 30290 19442 30363
rect 19517 30290 19583 30293
rect 19382 30288 19583 30290
rect 19382 30232 19522 30288
rect 19578 30232 19583 30288
rect 19382 30230 19583 30232
rect 19517 30227 19583 30230
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 19570 29408 19886 29409
rect 19570 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19886 29408
rect 19570 29343 19886 29344
rect 11697 29202 11763 29205
rect 17401 29202 17467 29205
rect 11697 29200 17467 29202
rect 11697 29144 11702 29200
rect 11758 29144 17406 29200
rect 17462 29144 17467 29200
rect 11697 29142 17467 29144
rect 11697 29139 11763 29142
rect 17401 29139 17467 29142
rect 13629 28930 13695 28933
rect 17217 28930 17283 28933
rect 23657 28930 23723 28933
rect 13629 28928 23723 28930
rect 13629 28872 13634 28928
rect 13690 28872 17222 28928
rect 17278 28872 23662 28928
rect 23718 28872 23723 28928
rect 13629 28870 23723 28872
rect 13629 28867 13695 28870
rect 17217 28867 17283 28870
rect 23657 28867 23723 28870
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 19570 28320 19886 28321
rect 19570 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19886 28320
rect 19570 28255 19886 28256
rect 2773 27978 2839 27981
rect 17493 27978 17559 27981
rect 2773 27976 17559 27978
rect 2773 27920 2778 27976
rect 2834 27920 17498 27976
rect 17554 27920 17559 27976
rect 2773 27918 17559 27920
rect 2773 27915 2839 27918
rect 17493 27915 17559 27918
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 4061 27434 4127 27437
rect 19701 27434 19767 27437
rect 4061 27432 19767 27434
rect 4061 27376 4066 27432
rect 4122 27376 19706 27432
rect 19762 27376 19767 27432
rect 4061 27374 19767 27376
rect 4061 27371 4127 27374
rect 19701 27371 19767 27374
rect 19570 27232 19886 27233
rect 19570 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19886 27232
rect 19570 27167 19886 27168
rect 19517 27026 19583 27029
rect 20805 27026 20871 27029
rect 19517 27024 20871 27026
rect 19517 26968 19522 27024
rect 19578 26968 20810 27024
rect 20866 26968 20871 27024
rect 19517 26966 20871 26968
rect 19517 26963 19583 26966
rect 19934 26893 19994 26966
rect 20805 26963 20871 26966
rect 19885 26888 19994 26893
rect 19885 26832 19890 26888
rect 19946 26832 19994 26888
rect 19885 26830 19994 26832
rect 19885 26827 19951 26830
rect 19425 26754 19491 26757
rect 20069 26754 20135 26757
rect 19425 26752 20135 26754
rect 19425 26696 19430 26752
rect 19486 26696 20074 26752
rect 20130 26696 20135 26752
rect 19425 26694 20135 26696
rect 19425 26691 19491 26694
rect 20069 26691 20135 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 4061 26482 4127 26485
rect 19149 26482 19215 26485
rect 4061 26480 19215 26482
rect 4061 26424 4066 26480
rect 4122 26424 19154 26480
rect 19210 26424 19215 26480
rect 4061 26422 19215 26424
rect 4061 26419 4127 26422
rect 19149 26419 19215 26422
rect 19333 26346 19399 26349
rect 20345 26346 20411 26349
rect 19333 26344 20411 26346
rect 19333 26288 19338 26344
rect 19394 26288 20350 26344
rect 20406 26288 20411 26344
rect 19333 26286 20411 26288
rect 19333 26283 19399 26286
rect 20345 26283 20411 26286
rect 19570 26144 19886 26145
rect 19570 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19886 26144
rect 19570 26079 19886 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 19701 25258 19767 25261
rect 20253 25258 20319 25261
rect 19701 25256 20319 25258
rect 19701 25200 19706 25256
rect 19762 25200 20258 25256
rect 20314 25200 20319 25256
rect 19701 25198 20319 25200
rect 19701 25195 19767 25198
rect 20253 25195 20319 25198
rect 19570 25056 19886 25057
rect 19570 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19886 25056
rect 19570 24991 19886 24992
rect 19425 24986 19491 24989
rect 19382 24984 19491 24986
rect 19382 24928 19430 24984
rect 19486 24928 19491 24984
rect 19382 24923 19491 24928
rect 19382 24717 19442 24923
rect 19333 24712 19442 24717
rect 19333 24656 19338 24712
rect 19394 24656 19442 24712
rect 19333 24654 19442 24656
rect 19333 24651 19399 24654
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 13537 24442 13603 24445
rect 16757 24442 16823 24445
rect 13537 24440 16823 24442
rect 13537 24384 13542 24440
rect 13598 24384 16762 24440
rect 16818 24384 16823 24440
rect 13537 24382 16823 24384
rect 13537 24379 13603 24382
rect 16757 24379 16823 24382
rect 19570 23968 19886 23969
rect 19570 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19886 23968
rect 19570 23903 19886 23904
rect 13813 23762 13879 23765
rect 14733 23762 14799 23765
rect 22737 23762 22803 23765
rect 13813 23760 22803 23762
rect 13813 23704 13818 23760
rect 13874 23704 14738 23760
rect 14794 23704 22742 23760
rect 22798 23704 22803 23760
rect 13813 23702 22803 23704
rect 13813 23699 13879 23702
rect 14733 23699 14799 23702
rect 22737 23699 22803 23702
rect 16205 23490 16271 23493
rect 17585 23490 17651 23493
rect 16205 23488 17651 23490
rect 16205 23432 16210 23488
rect 16266 23432 17590 23488
rect 17646 23432 17651 23488
rect 16205 23430 17651 23432
rect 16205 23427 16271 23430
rect 17585 23427 17651 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 14641 23218 14707 23221
rect 17309 23218 17375 23221
rect 14641 23216 17375 23218
rect 14641 23160 14646 23216
rect 14702 23160 17314 23216
rect 17370 23160 17375 23216
rect 14641 23158 17375 23160
rect 14641 23155 14707 23158
rect 17309 23155 17375 23158
rect 16573 23082 16639 23085
rect 18137 23082 18203 23085
rect 16573 23080 18203 23082
rect 16573 23024 16578 23080
rect 16634 23024 18142 23080
rect 18198 23024 18203 23080
rect 16573 23022 18203 23024
rect 16573 23019 16639 23022
rect 18137 23019 18203 23022
rect 19570 22880 19886 22881
rect 19570 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19886 22880
rect 19570 22815 19886 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19570 21792 19886 21793
rect 19570 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19886 21792
rect 19570 21727 19886 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 19570 20704 19886 20705
rect 19570 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19886 20704
rect 19570 20639 19886 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 19570 19616 19886 19617
rect 19570 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19886 19616
rect 19570 19551 19886 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 19570 18528 19886 18529
rect 19570 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19886 18528
rect 19570 18463 19886 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 0 17778 800 17808
rect 1393 17778 1459 17781
rect 0 17776 1459 17778
rect 0 17720 1398 17776
rect 1454 17720 1459 17776
rect 0 17718 1459 17720
rect 0 17688 800 17718
rect 1393 17715 1459 17718
rect 19570 17440 19886 17441
rect 19570 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19886 17440
rect 19570 17375 19886 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 19570 16352 19886 16353
rect 19570 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19886 16352
rect 19570 16287 19886 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 19570 15264 19886 15265
rect 19570 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19886 15264
rect 19570 15199 19886 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 19570 14176 19886 14177
rect 19570 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19886 14176
rect 19570 14111 19886 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 19570 13088 19886 13089
rect 19570 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19886 13088
rect 19570 13023 19886 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 38101 12338 38167 12341
rect 39200 12338 40000 12368
rect 38101 12336 40000 12338
rect 38101 12280 38106 12336
rect 38162 12280 40000 12336
rect 38101 12278 40000 12280
rect 38101 12275 38167 12278
rect 39200 12248 40000 12278
rect 19570 12000 19886 12001
rect 19570 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19886 12000
rect 19570 11935 19886 11936
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 19570 10912 19886 10913
rect 19570 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19886 10912
rect 19570 10847 19886 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 19570 9824 19886 9825
rect 19570 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19886 9824
rect 19570 9759 19886 9760
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 19570 8736 19886 8737
rect 19570 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19886 8736
rect 19570 8671 19886 8672
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 19570 7648 19886 7649
rect 19570 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19886 7648
rect 19570 7583 19886 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 19570 6560 19886 6561
rect 19570 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19886 6560
rect 19570 6495 19886 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 19570 5472 19886 5473
rect 19570 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19886 5472
rect 19570 5407 19886 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 19570 4384 19886 4385
rect 19570 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19886 4384
rect 19570 4319 19886 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 19570 3296 19886 3297
rect 19570 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19886 3296
rect 19570 3231 19886 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 19570 2208 19886 2209
rect 19570 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19886 2208
rect 19570 2143 19886 2144
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA__114__S opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17480 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__115__A
timestamp 1649977179
transform -1 0 37444 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__117__A
timestamp 1649977179
transform 1 0 22540 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__118__B1
timestamp 1649977179
transform 1 0 20700 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__122__B1
timestamp 1649977179
transform 1 0 21160 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__123__B1
timestamp 1649977179
transform 1 0 19964 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__124__A
timestamp 1649977179
transform -1 0 23920 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__125__B1_N
timestamp 1649977179
transform 1 0 21712 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__126__B
timestamp 1649977179
transform 1 0 20516 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__127__B
timestamp 1649977179
transform 1 0 20608 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__128__B1
timestamp 1649977179
transform 1 0 21620 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__131__B
timestamp 1649977179
transform 1 0 18584 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__A2
timestamp 1649977179
transform -1 0 24564 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__132__B1_N
timestamp 1649977179
transform -1 0 24564 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__A_N
timestamp 1649977179
transform 1 0 21896 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__133__B
timestamp 1649977179
transform 1 0 21528 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__A_N
timestamp 1649977179
transform -1 0 24012 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__134__B
timestamp 1649977179
transform -1 0 23828 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__135__B1
timestamp 1649977179
transform 1 0 22908 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__A
timestamp 1649977179
transform 1 0 19228 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__137__B_N
timestamp 1649977179
transform 1 0 18860 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__A1
timestamp 1649977179
transform 1 0 20424 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__138__B1
timestamp 1649977179
transform 1 0 18584 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__A2
timestamp 1649977179
transform -1 0 22908 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__139__B1_N
timestamp 1649977179
transform 1 0 22172 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__A_N
timestamp 1649977179
transform -1 0 18860 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__140__B
timestamp 1649977179
transform -1 0 18308 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__142__B
timestamp 1649977179
transform -1 0 22540 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__143__A
timestamp 1649977179
transform -1 0 22908 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__144__A1
timestamp 1649977179
transform -1 0 21988 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__A2
timestamp 1649977179
transform -1 0 15916 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__145__B1
timestamp 1649977179
transform 1 0 14444 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A1
timestamp 1649977179
transform 1 0 19412 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__A2
timestamp 1649977179
transform 1 0 19596 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__146__B2
timestamp 1649977179
transform -1 0 21068 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A1
timestamp 1649977179
transform 1 0 16008 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__147__A2
timestamp 1649977179
transform 1 0 17572 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__149__A
timestamp 1649977179
transform 1 0 23276 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__A2
timestamp 1649977179
transform 1 0 20516 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__150__B1
timestamp 1649977179
transform -1 0 20516 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__A1
timestamp 1649977179
transform -1 0 11500 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__153__A2
timestamp 1649977179
transform 1 0 12972 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__A
timestamp 1649977179
transform 1 0 12788 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__154__B
timestamp 1649977179
transform 1 0 12420 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A1
timestamp 1649977179
transform 1 0 16652 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__A2
timestamp 1649977179
transform 1 0 16008 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__157__B1
timestamp 1649977179
transform 1 0 15456 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__A
timestamp 1649977179
transform 1 0 13432 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__B
timestamp 1649977179
transform 1 0 15180 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__158__D
timestamp 1649977179
transform 1 0 14076 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__159__A2
timestamp 1649977179
transform 1 0 16100 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__160__A1
timestamp 1649977179
transform 1 0 9568 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__161__A1
timestamp 1649977179
transform 1 0 10304 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__A
timestamp 1649977179
transform 1 0 12420 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__B
timestamp 1649977179
transform 1 0 12604 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__162__C
timestamp 1649977179
transform 1 0 13340 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__A1
timestamp 1649977179
transform 1 0 11684 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__163__B1
timestamp 1649977179
transform -1 0 12512 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__165__A1
timestamp 1649977179
transform 1 0 14352 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__165__A2
timestamp 1649977179
transform 1 0 15088 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__170__B1
timestamp 1649977179
transform 1 0 19780 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__171__B
timestamp 1649977179
transform -1 0 21344 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__173__A2
timestamp 1649977179
transform 1 0 19780 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__174__B1
timestamp 1649977179
transform 1 0 20976 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__176__A2
timestamp 1649977179
transform 1 0 17756 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__188__B
timestamp 1649977179
transform -1 0 16744 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__199__A2
timestamp 1649977179
transform 1 0 14260 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__200__A2
timestamp 1649977179
transform -1 0 19320 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__200__B1
timestamp 1649977179
transform 1 0 18584 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__203__A
timestamp 1649977179
transform 1 0 10488 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__A3
timestamp 1649977179
transform 1 0 20148 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__A4
timestamp 1649977179
transform 1 0 18584 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__206__B1
timestamp 1649977179
transform -1 0 21252 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__208__A
timestamp 1649977179
transform 1 0 18492 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__A2
timestamp 1649977179
transform 1 0 18952 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__A3
timestamp 1649977179
transform 1 0 18308 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__209__B1
timestamp 1649977179
transform 1 0 17756 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A2
timestamp 1649977179
transform 1 0 20240 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__A3
timestamp 1649977179
transform 1 0 18032 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__211__B1
timestamp 1649977179
transform 1 0 18584 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A1
timestamp 1649977179
transform 1 0 12420 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__A2
timestamp 1649977179
transform 1 0 11132 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__213__B1
timestamp 1649977179
transform -1 0 11040 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__214__A
timestamp 1649977179
transform -1 0 9384 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__216__B
timestamp 1649977179
transform 1 0 15732 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__217__A2
timestamp 1649977179
transform 1 0 9844 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__218__A1
timestamp 1649977179
transform -1 0 12420 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__220__A1
timestamp 1649977179
transform -1 0 15640 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__222__A1
timestamp 1649977179
transform 1 0 15272 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__245__D
timestamp 1649977179
transform -1 0 3404 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_clkbuf_0_i_clk_A
timestamp 1649977179
transform -1 0 9384 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1649977179
transform -1 0 1564 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1649977179
transform -1 0 35052 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1649977179
transform -1 0 30636 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1649977179
transform -1 0 38180 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1649977179
transform -1 0 2208 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1649977179
transform -1 0 17664 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1649977179
transform -1 0 14444 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 2300 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29
timestamp 1649977179
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41
timestamp 1649977179
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53
timestamp 1649977179
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57
timestamp 1649977179
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69
timestamp 1649977179
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_81
timestamp 1649977179
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_85
timestamp 1649977179
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_97
timestamp 1649977179
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_109
timestamp 1649977179
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_113
timestamp 1649977179
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_125
timestamp 1649977179
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1649977179
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_141
timestamp 1649977179
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_153
timestamp 1649977179
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_165
timestamp 1649977179
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_169 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 16652 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_174 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 17112 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_180
timestamp 1649977179
transform 1 0 17664 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_192
timestamp 1649977179
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_197
timestamp 1649977179
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_209
timestamp 1649977179
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_221
timestamp 1649977179
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_225
timestamp 1649977179
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_237
timestamp 1649977179
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_249
timestamp 1649977179
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_253
timestamp 1649977179
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_265
timestamp 1649977179
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_277
timestamp 1649977179
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_281
timestamp 1649977179
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_293
timestamp 1649977179
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_305
timestamp 1649977179
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_309
timestamp 1649977179
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_321
timestamp 1649977179
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_333
timestamp 1649977179
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_337
timestamp 1649977179
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_349
timestamp 1649977179
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_361
timestamp 1649977179
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_365
timestamp 1649977179
transform 1 0 34684 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_373
timestamp 1649977179
transform 1 0 35420 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_393
timestamp 1649977179
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_405
timestamp 1649977179
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_1_5
timestamp 1649977179
transform 1 0 1564 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_17
timestamp 1649977179
transform 1 0 2668 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_29
timestamp 1649977179
transform 1 0 3772 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_41
timestamp 1649977179
transform 1 0 4876 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_53
timestamp 1649977179
transform 1 0 5980 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_57
timestamp 1649977179
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_69
timestamp 1649977179
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_81
timestamp 1649977179
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_93
timestamp 1649977179
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_105
timestamp 1649977179
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_111
timestamp 1649977179
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_113
timestamp 1649977179
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_125
timestamp 1649977179
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_137
timestamp 1649977179
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_149
timestamp 1649977179
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_161
timestamp 1649977179
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1649977179
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_169
timestamp 1649977179
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_181
timestamp 1649977179
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_193
timestamp 1649977179
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_205
timestamp 1649977179
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_217
timestamp 1649977179
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1649977179
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_225
timestamp 1649977179
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_237
timestamp 1649977179
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_249
timestamp 1649977179
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_261
timestamp 1649977179
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_273
timestamp 1649977179
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_279
timestamp 1649977179
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_281
timestamp 1649977179
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_293
timestamp 1649977179
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_305
timestamp 1649977179
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_317
timestamp 1649977179
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_329
timestamp 1649977179
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1649977179
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_1_337
timestamp 1649977179
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_1_349
timestamp 1649977179
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_361
timestamp 1649977179
transform 1 0 34316 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_1_369
timestamp 1649977179
transform 1 0 35052 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_381 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 36156 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_389
timestamp 1649977179
transform 1 0 36892 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_1_393
timestamp 1649977179
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1649977179
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_2_3
timestamp 1649977179
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_15
timestamp 1649977179
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_27
timestamp 1649977179
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_29
timestamp 1649977179
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_41
timestamp 1649977179
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_53
timestamp 1649977179
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_65
timestamp 1649977179
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1649977179
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1649977179
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_85
timestamp 1649977179
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_97
timestamp 1649977179
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_109
timestamp 1649977179
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_121
timestamp 1649977179
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_133
timestamp 1649977179
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_139
timestamp 1649977179
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_141
timestamp 1649977179
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_153
timestamp 1649977179
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_165
timestamp 1649977179
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_177
timestamp 1649977179
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_189
timestamp 1649977179
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1649977179
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_197
timestamp 1649977179
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_209
timestamp 1649977179
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_221
timestamp 1649977179
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_233
timestamp 1649977179
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_245
timestamp 1649977179
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_251
timestamp 1649977179
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_253
timestamp 1649977179
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_265
timestamp 1649977179
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_277
timestamp 1649977179
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_289
timestamp 1649977179
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_301
timestamp 1649977179
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_307
timestamp 1649977179
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_309
timestamp 1649977179
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_321
timestamp 1649977179
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_333
timestamp 1649977179
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_345
timestamp 1649977179
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1649977179
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1649977179
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_2_365
timestamp 1649977179
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_377
timestamp 1649977179
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_2_389
timestamp 1649977179
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_401
timestamp 1649977179
transform 1 0 37996 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_3_3
timestamp 1649977179
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_15
timestamp 1649977179
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_27
timestamp 1649977179
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_39
timestamp 1649977179
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1649977179
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1649977179
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_57
timestamp 1649977179
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_69
timestamp 1649977179
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_81
timestamp 1649977179
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_93
timestamp 1649977179
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_105
timestamp 1649977179
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1649977179
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_113
timestamp 1649977179
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_125
timestamp 1649977179
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_137
timestamp 1649977179
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_149
timestamp 1649977179
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_161
timestamp 1649977179
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_167
timestamp 1649977179
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_169
timestamp 1649977179
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_181
timestamp 1649977179
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_193
timestamp 1649977179
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_205
timestamp 1649977179
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1649977179
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1649977179
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_225
timestamp 1649977179
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_237
timestamp 1649977179
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_249
timestamp 1649977179
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_261
timestamp 1649977179
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_273
timestamp 1649977179
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1649977179
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_281
timestamp 1649977179
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_293
timestamp 1649977179
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_305
timestamp 1649977179
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_317
timestamp 1649977179
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1649977179
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1649977179
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_337
timestamp 1649977179
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_349
timestamp 1649977179
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_361
timestamp 1649977179
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_3_373
timestamp 1649977179
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_385
timestamp 1649977179
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1649977179
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_3_393
timestamp 1649977179
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_405
timestamp 1649977179
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_4_3
timestamp 1649977179
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_15
timestamp 1649977179
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1649977179
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_29
timestamp 1649977179
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_41
timestamp 1649977179
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_53
timestamp 1649977179
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_65
timestamp 1649977179
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_77
timestamp 1649977179
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1649977179
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_85
timestamp 1649977179
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_97
timestamp 1649977179
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_109
timestamp 1649977179
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_121
timestamp 1649977179
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1649977179
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1649977179
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_141
timestamp 1649977179
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_153
timestamp 1649977179
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_165
timestamp 1649977179
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_177
timestamp 1649977179
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1649977179
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1649977179
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_197
timestamp 1649977179
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_209
timestamp 1649977179
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_221
timestamp 1649977179
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_233
timestamp 1649977179
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_245
timestamp 1649977179
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_251
timestamp 1649977179
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_253
timestamp 1649977179
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_265
timestamp 1649977179
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_277
timestamp 1649977179
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_289
timestamp 1649977179
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1649977179
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1649977179
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_309
timestamp 1649977179
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_321
timestamp 1649977179
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_333
timestamp 1649977179
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_345
timestamp 1649977179
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_357
timestamp 1649977179
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1649977179
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_4_365
timestamp 1649977179
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_377
timestamp 1649977179
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_4_389
timestamp 1649977179
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_401
timestamp 1649977179
transform 1 0 37996 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_5_3
timestamp 1649977179
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_15
timestamp 1649977179
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_27
timestamp 1649977179
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_39
timestamp 1649977179
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_51
timestamp 1649977179
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1649977179
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_57
timestamp 1649977179
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_69
timestamp 1649977179
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_81
timestamp 1649977179
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_93
timestamp 1649977179
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1649977179
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1649977179
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_113
timestamp 1649977179
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_125
timestamp 1649977179
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_137
timestamp 1649977179
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_149
timestamp 1649977179
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1649977179
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1649977179
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_169
timestamp 1649977179
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_181
timestamp 1649977179
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_193
timestamp 1649977179
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_205
timestamp 1649977179
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1649977179
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1649977179
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_225
timestamp 1649977179
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_237
timestamp 1649977179
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_249
timestamp 1649977179
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_261
timestamp 1649977179
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1649977179
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1649977179
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_281
timestamp 1649977179
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_293
timestamp 1649977179
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_305
timestamp 1649977179
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_317
timestamp 1649977179
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1649977179
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1649977179
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_337
timestamp 1649977179
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_349
timestamp 1649977179
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_361
timestamp 1649977179
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_5_373
timestamp 1649977179
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1649977179
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1649977179
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_5_393
timestamp 1649977179
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_405
timestamp 1649977179
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_6_3
timestamp 1649977179
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_15
timestamp 1649977179
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1649977179
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_29
timestamp 1649977179
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_41
timestamp 1649977179
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_53
timestamp 1649977179
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_65
timestamp 1649977179
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1649977179
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1649977179
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_85
timestamp 1649977179
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_97
timestamp 1649977179
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_109
timestamp 1649977179
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_121
timestamp 1649977179
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1649977179
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1649977179
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_141
timestamp 1649977179
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_153
timestamp 1649977179
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_165
timestamp 1649977179
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_177
timestamp 1649977179
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1649977179
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1649977179
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_197
timestamp 1649977179
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_209
timestamp 1649977179
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_221
timestamp 1649977179
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_233
timestamp 1649977179
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1649977179
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1649977179
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_253
timestamp 1649977179
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_265
timestamp 1649977179
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_277
timestamp 1649977179
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_289
timestamp 1649977179
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_301
timestamp 1649977179
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1649977179
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_309
timestamp 1649977179
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_321
timestamp 1649977179
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_333
timestamp 1649977179
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_345
timestamp 1649977179
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1649977179
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1649977179
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_6_365
timestamp 1649977179
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_377
timestamp 1649977179
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_6_389
timestamp 1649977179
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_401
timestamp 1649977179
transform 1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_7_3
timestamp 1649977179
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_15
timestamp 1649977179
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_27
timestamp 1649977179
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_39
timestamp 1649977179
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_51
timestamp 1649977179
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_55
timestamp 1649977179
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_57
timestamp 1649977179
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_69
timestamp 1649977179
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_81
timestamp 1649977179
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_93
timestamp 1649977179
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1649977179
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1649977179
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_113
timestamp 1649977179
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_125
timestamp 1649977179
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_137
timestamp 1649977179
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_149
timestamp 1649977179
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1649977179
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1649977179
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_169
timestamp 1649977179
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_181
timestamp 1649977179
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_193
timestamp 1649977179
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_205
timestamp 1649977179
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1649977179
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1649977179
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_225
timestamp 1649977179
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_237
timestamp 1649977179
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_249
timestamp 1649977179
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_261
timestamp 1649977179
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_273
timestamp 1649977179
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_279
timestamp 1649977179
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_281
timestamp 1649977179
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_293
timestamp 1649977179
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_305
timestamp 1649977179
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_317
timestamp 1649977179
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1649977179
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1649977179
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_337
timestamp 1649977179
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_349
timestamp 1649977179
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_361
timestamp 1649977179
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_7_373
timestamp 1649977179
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1649977179
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1649977179
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_7_393
timestamp 1649977179
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_405
timestamp 1649977179
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_8_3
timestamp 1649977179
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_15
timestamp 1649977179
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1649977179
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_29
timestamp 1649977179
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_41
timestamp 1649977179
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_53
timestamp 1649977179
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_65
timestamp 1649977179
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1649977179
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1649977179
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_85
timestamp 1649977179
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_97
timestamp 1649977179
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_109
timestamp 1649977179
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_121
timestamp 1649977179
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1649977179
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1649977179
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_141
timestamp 1649977179
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_153
timestamp 1649977179
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_165
timestamp 1649977179
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_177
timestamp 1649977179
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1649977179
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1649977179
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_197
timestamp 1649977179
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_209
timestamp 1649977179
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_221
timestamp 1649977179
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_233
timestamp 1649977179
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1649977179
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1649977179
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_253
timestamp 1649977179
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_265
timestamp 1649977179
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_277
timestamp 1649977179
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_289
timestamp 1649977179
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1649977179
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1649977179
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_309
timestamp 1649977179
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_321
timestamp 1649977179
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_333
timestamp 1649977179
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_345
timestamp 1649977179
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_357
timestamp 1649977179
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_363
timestamp 1649977179
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_8_365
timestamp 1649977179
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_377
timestamp 1649977179
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_8_389
timestamp 1649977179
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_401
timestamp 1649977179
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_9_3
timestamp 1649977179
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_15
timestamp 1649977179
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_27
timestamp 1649977179
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_39
timestamp 1649977179
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1649977179
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1649977179
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_57
timestamp 1649977179
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_69
timestamp 1649977179
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_81
timestamp 1649977179
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_93
timestamp 1649977179
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1649977179
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1649977179
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_113
timestamp 1649977179
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_125
timestamp 1649977179
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_137
timestamp 1649977179
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_149
timestamp 1649977179
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1649977179
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1649977179
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_169
timestamp 1649977179
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_181
timestamp 1649977179
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_193
timestamp 1649977179
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_205
timestamp 1649977179
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_217
timestamp 1649977179
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_223
timestamp 1649977179
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_225
timestamp 1649977179
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_237
timestamp 1649977179
transform 1 0 22908 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_249
timestamp 1649977179
transform 1 0 24012 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_261
timestamp 1649977179
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1649977179
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1649977179
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_281
timestamp 1649977179
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_293
timestamp 1649977179
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_305
timestamp 1649977179
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_317
timestamp 1649977179
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_329
timestamp 1649977179
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1649977179
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_337
timestamp 1649977179
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_349
timestamp 1649977179
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_361
timestamp 1649977179
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_9_373
timestamp 1649977179
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1649977179
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1649977179
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_9_393
timestamp 1649977179
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_405
timestamp 1649977179
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_10_3
timestamp 1649977179
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_15
timestamp 1649977179
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1649977179
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_29
timestamp 1649977179
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_41
timestamp 1649977179
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_53
timestamp 1649977179
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_65
timestamp 1649977179
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1649977179
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1649977179
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_85
timestamp 1649977179
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_97
timestamp 1649977179
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_109
timestamp 1649977179
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_121
timestamp 1649977179
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1649977179
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1649977179
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_141
timestamp 1649977179
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_153
timestamp 1649977179
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_165
timestamp 1649977179
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_177
timestamp 1649977179
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_189
timestamp 1649977179
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1649977179
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_197
timestamp 1649977179
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_209
timestamp 1649977179
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_221
timestamp 1649977179
transform 1 0 21436 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_233
timestamp 1649977179
transform 1 0 22540 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_245
timestamp 1649977179
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_251
timestamp 1649977179
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_253
timestamp 1649977179
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_265
timestamp 1649977179
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_277
timestamp 1649977179
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_289
timestamp 1649977179
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_301
timestamp 1649977179
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_307
timestamp 1649977179
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_309
timestamp 1649977179
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_321
timestamp 1649977179
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_333
timestamp 1649977179
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_345
timestamp 1649977179
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_357
timestamp 1649977179
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1649977179
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_10_365
timestamp 1649977179
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_377
timestamp 1649977179
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_10_389
timestamp 1649977179
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_401
timestamp 1649977179
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_11_3
timestamp 1649977179
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_15
timestamp 1649977179
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_27
timestamp 1649977179
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_39
timestamp 1649977179
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1649977179
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1649977179
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_57
timestamp 1649977179
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_69
timestamp 1649977179
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_81
timestamp 1649977179
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_93
timestamp 1649977179
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1649977179
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1649977179
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_113
timestamp 1649977179
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_125
timestamp 1649977179
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_137
timestamp 1649977179
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_149
timestamp 1649977179
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1649977179
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1649977179
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_169
timestamp 1649977179
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_181
timestamp 1649977179
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_193
timestamp 1649977179
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_205
timestamp 1649977179
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_217
timestamp 1649977179
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_223
timestamp 1649977179
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_225
timestamp 1649977179
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_237
timestamp 1649977179
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_249
timestamp 1649977179
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_261
timestamp 1649977179
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1649977179
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1649977179
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_281
timestamp 1649977179
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_293
timestamp 1649977179
transform 1 0 28060 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_305
timestamp 1649977179
transform 1 0 29164 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_317
timestamp 1649977179
transform 1 0 30268 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_329
timestamp 1649977179
transform 1 0 31372 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1649977179
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_337
timestamp 1649977179
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_349
timestamp 1649977179
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_361
timestamp 1649977179
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_11_373
timestamp 1649977179
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1649977179
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1649977179
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_11_393
timestamp 1649977179
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_405
timestamp 1649977179
transform 1 0 38364 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_12_3
timestamp 1649977179
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_15
timestamp 1649977179
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1649977179
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_29
timestamp 1649977179
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_41
timestamp 1649977179
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_53
timestamp 1649977179
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_65
timestamp 1649977179
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1649977179
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1649977179
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_85
timestamp 1649977179
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_97
timestamp 1649977179
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_109
timestamp 1649977179
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_121
timestamp 1649977179
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1649977179
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1649977179
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_141
timestamp 1649977179
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_153
timestamp 1649977179
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_165
timestamp 1649977179
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_177
timestamp 1649977179
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_189
timestamp 1649977179
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_195
timestamp 1649977179
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_197
timestamp 1649977179
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_209
timestamp 1649977179
transform 1 0 20332 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_221
timestamp 1649977179
transform 1 0 21436 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_233
timestamp 1649977179
transform 1 0 22540 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_245
timestamp 1649977179
transform 1 0 23644 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1649977179
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_253
timestamp 1649977179
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_265
timestamp 1649977179
transform 1 0 25484 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_277
timestamp 1649977179
transform 1 0 26588 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_289
timestamp 1649977179
transform 1 0 27692 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_301
timestamp 1649977179
transform 1 0 28796 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1649977179
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_309
timestamp 1649977179
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_321
timestamp 1649977179
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_333
timestamp 1649977179
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_345
timestamp 1649977179
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1649977179
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1649977179
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_12_365
timestamp 1649977179
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_377
timestamp 1649977179
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_12_389
timestamp 1649977179
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_401
timestamp 1649977179
transform 1 0 37996 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_13_3
timestamp 1649977179
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_15
timestamp 1649977179
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_27
timestamp 1649977179
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_39
timestamp 1649977179
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1649977179
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1649977179
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_57
timestamp 1649977179
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_69
timestamp 1649977179
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_81
timestamp 1649977179
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_93
timestamp 1649977179
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1649977179
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1649977179
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_113
timestamp 1649977179
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_125
timestamp 1649977179
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_137
timestamp 1649977179
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_149
timestamp 1649977179
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1649977179
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1649977179
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_169
timestamp 1649977179
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_181
timestamp 1649977179
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_193
timestamp 1649977179
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_205
timestamp 1649977179
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_217
timestamp 1649977179
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1649977179
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_225
timestamp 1649977179
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_237
timestamp 1649977179
transform 1 0 22908 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_249
timestamp 1649977179
transform 1 0 24012 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_261
timestamp 1649977179
transform 1 0 25116 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_273
timestamp 1649977179
transform 1 0 26220 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_279
timestamp 1649977179
transform 1 0 26772 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_281
timestamp 1649977179
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_293
timestamp 1649977179
transform 1 0 28060 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_305
timestamp 1649977179
transform 1 0 29164 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_317
timestamp 1649977179
transform 1 0 30268 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_329
timestamp 1649977179
transform 1 0 31372 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1649977179
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_337
timestamp 1649977179
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_349
timestamp 1649977179
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_361
timestamp 1649977179
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_13_373
timestamp 1649977179
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1649977179
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1649977179
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_13_393
timestamp 1649977179
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_405
timestamp 1649977179
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_14_3
timestamp 1649977179
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_15
timestamp 1649977179
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1649977179
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_29
timestamp 1649977179
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_41
timestamp 1649977179
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_53
timestamp 1649977179
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_65
timestamp 1649977179
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1649977179
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1649977179
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_85
timestamp 1649977179
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_97
timestamp 1649977179
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_109
timestamp 1649977179
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_121
timestamp 1649977179
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1649977179
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1649977179
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_141
timestamp 1649977179
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_153
timestamp 1649977179
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_165
timestamp 1649977179
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_177
timestamp 1649977179
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1649977179
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1649977179
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_197
timestamp 1649977179
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_209
timestamp 1649977179
transform 1 0 20332 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_221
timestamp 1649977179
transform 1 0 21436 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_233
timestamp 1649977179
transform 1 0 22540 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_245
timestamp 1649977179
transform 1 0 23644 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_251
timestamp 1649977179
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_253
timestamp 1649977179
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_265
timestamp 1649977179
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_277
timestamp 1649977179
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_289
timestamp 1649977179
transform 1 0 27692 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_301
timestamp 1649977179
transform 1 0 28796 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1649977179
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_309
timestamp 1649977179
transform 1 0 29532 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_321
timestamp 1649977179
transform 1 0 30636 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_333
timestamp 1649977179
transform 1 0 31740 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_345
timestamp 1649977179
transform 1 0 32844 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_357
timestamp 1649977179
transform 1 0 33948 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1649977179
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_14_365
timestamp 1649977179
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_377
timestamp 1649977179
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_14_389
timestamp 1649977179
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_401
timestamp 1649977179
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_15_3
timestamp 1649977179
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_15
timestamp 1649977179
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_27
timestamp 1649977179
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_39
timestamp 1649977179
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1649977179
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1649977179
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_57
timestamp 1649977179
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_69
timestamp 1649977179
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_81
timestamp 1649977179
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_93
timestamp 1649977179
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1649977179
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1649977179
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_113
timestamp 1649977179
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_125
timestamp 1649977179
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_137
timestamp 1649977179
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_149
timestamp 1649977179
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1649977179
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1649977179
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_169
timestamp 1649977179
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_181
timestamp 1649977179
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_193
timestamp 1649977179
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_205
timestamp 1649977179
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_217
timestamp 1649977179
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1649977179
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_225
timestamp 1649977179
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_237
timestamp 1649977179
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_249
timestamp 1649977179
transform 1 0 24012 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_261
timestamp 1649977179
transform 1 0 25116 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_273
timestamp 1649977179
transform 1 0 26220 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_279
timestamp 1649977179
transform 1 0 26772 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_281
timestamp 1649977179
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_293
timestamp 1649977179
transform 1 0 28060 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_305
timestamp 1649977179
transform 1 0 29164 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_317
timestamp 1649977179
transform 1 0 30268 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_329
timestamp 1649977179
transform 1 0 31372 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_335
timestamp 1649977179
transform 1 0 31924 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_337
timestamp 1649977179
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_349
timestamp 1649977179
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_361
timestamp 1649977179
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_15_373
timestamp 1649977179
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1649977179
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1649977179
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_15_393
timestamp 1649977179
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_405
timestamp 1649977179
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_16_3
timestamp 1649977179
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_15
timestamp 1649977179
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1649977179
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_29
timestamp 1649977179
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_41
timestamp 1649977179
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_53
timestamp 1649977179
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_65
timestamp 1649977179
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1649977179
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1649977179
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_85
timestamp 1649977179
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_97
timestamp 1649977179
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_109
timestamp 1649977179
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_121
timestamp 1649977179
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1649977179
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1649977179
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_141
timestamp 1649977179
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_153
timestamp 1649977179
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_165
timestamp 1649977179
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_177
timestamp 1649977179
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_189
timestamp 1649977179
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1649977179
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_197
timestamp 1649977179
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_209
timestamp 1649977179
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_221
timestamp 1649977179
transform 1 0 21436 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_233
timestamp 1649977179
transform 1 0 22540 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_245
timestamp 1649977179
transform 1 0 23644 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1649977179
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_253
timestamp 1649977179
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_265
timestamp 1649977179
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_277
timestamp 1649977179
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_289
timestamp 1649977179
transform 1 0 27692 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_301
timestamp 1649977179
transform 1 0 28796 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1649977179
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_309
timestamp 1649977179
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_321
timestamp 1649977179
transform 1 0 30636 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_333
timestamp 1649977179
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_345
timestamp 1649977179
transform 1 0 32844 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_357
timestamp 1649977179
transform 1 0 33948 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_363
timestamp 1649977179
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_16_365
timestamp 1649977179
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_377
timestamp 1649977179
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_16_389
timestamp 1649977179
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_401
timestamp 1649977179
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_17_3
timestamp 1649977179
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_15
timestamp 1649977179
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_27
timestamp 1649977179
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_39
timestamp 1649977179
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_51
timestamp 1649977179
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_55
timestamp 1649977179
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_57
timestamp 1649977179
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_69
timestamp 1649977179
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_81
timestamp 1649977179
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_93
timestamp 1649977179
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1649977179
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1649977179
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_113
timestamp 1649977179
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_125
timestamp 1649977179
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_137
timestamp 1649977179
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_149
timestamp 1649977179
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1649977179
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1649977179
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_169
timestamp 1649977179
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_181
timestamp 1649977179
transform 1 0 17756 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_193
timestamp 1649977179
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_205
timestamp 1649977179
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_217
timestamp 1649977179
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1649977179
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_225
timestamp 1649977179
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_237
timestamp 1649977179
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_249
timestamp 1649977179
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_261
timestamp 1649977179
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_273
timestamp 1649977179
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1649977179
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_281
timestamp 1649977179
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_293
timestamp 1649977179
transform 1 0 28060 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_305
timestamp 1649977179
transform 1 0 29164 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_317
timestamp 1649977179
transform 1 0 30268 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_329
timestamp 1649977179
transform 1 0 31372 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_335
timestamp 1649977179
transform 1 0 31924 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_337
timestamp 1649977179
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_349
timestamp 1649977179
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_361
timestamp 1649977179
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_17_373
timestamp 1649977179
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1649977179
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1649977179
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_17_393
timestamp 1649977179
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_405
timestamp 1649977179
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_18_3
timestamp 1649977179
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_15
timestamp 1649977179
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1649977179
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_29
timestamp 1649977179
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_41
timestamp 1649977179
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_53
timestamp 1649977179
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_65
timestamp 1649977179
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1649977179
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1649977179
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_85
timestamp 1649977179
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_97
timestamp 1649977179
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_109
timestamp 1649977179
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_121
timestamp 1649977179
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1649977179
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1649977179
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_141
timestamp 1649977179
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_153
timestamp 1649977179
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_165
timestamp 1649977179
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_177
timestamp 1649977179
transform 1 0 17388 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_189
timestamp 1649977179
transform 1 0 18492 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_195
timestamp 1649977179
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_197
timestamp 1649977179
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_209
timestamp 1649977179
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_221
timestamp 1649977179
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_233
timestamp 1649977179
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_245
timestamp 1649977179
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_251
timestamp 1649977179
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_253
timestamp 1649977179
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_265
timestamp 1649977179
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_277
timestamp 1649977179
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_289
timestamp 1649977179
transform 1 0 27692 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_301
timestamp 1649977179
transform 1 0 28796 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_307
timestamp 1649977179
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_309
timestamp 1649977179
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_321
timestamp 1649977179
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_333
timestamp 1649977179
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_345
timestamp 1649977179
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_357
timestamp 1649977179
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_363
timestamp 1649977179
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_18_365
timestamp 1649977179
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_18_377
timestamp 1649977179
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_389
timestamp 1649977179
transform 1 0 36892 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_397
timestamp 1649977179
transform 1 0 37628 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_403
timestamp 1649977179
transform 1 0 38180 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_19_3
timestamp 1649977179
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_15
timestamp 1649977179
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_27
timestamp 1649977179
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_39
timestamp 1649977179
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_51
timestamp 1649977179
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1649977179
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_57
timestamp 1649977179
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_69
timestamp 1649977179
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_81
timestamp 1649977179
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_93
timestamp 1649977179
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1649977179
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1649977179
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_113
timestamp 1649977179
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_125
timestamp 1649977179
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_137
timestamp 1649977179
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_149
timestamp 1649977179
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1649977179
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1649977179
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_169
timestamp 1649977179
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_181
timestamp 1649977179
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_193
timestamp 1649977179
transform 1 0 18860 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_205
timestamp 1649977179
transform 1 0 19964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_217
timestamp 1649977179
transform 1 0 21068 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1649977179
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_225
timestamp 1649977179
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_237
timestamp 1649977179
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_249
timestamp 1649977179
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_261
timestamp 1649977179
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_273
timestamp 1649977179
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_279
timestamp 1649977179
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_281
timestamp 1649977179
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_293
timestamp 1649977179
transform 1 0 28060 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_305
timestamp 1649977179
transform 1 0 29164 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_317
timestamp 1649977179
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1649977179
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1649977179
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_19_337
timestamp 1649977179
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_349
timestamp 1649977179
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_361
timestamp 1649977179
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_19_373
timestamp 1649977179
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_385
timestamp 1649977179
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_391
timestamp 1649977179
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_395
timestamp 1649977179
transform 1 0 37444 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_402
timestamp 1649977179
transform 1 0 38088 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_406
timestamp 1649977179
transform 1 0 38456 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_3
timestamp 1649977179
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_15
timestamp 1649977179
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_27
timestamp 1649977179
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_29
timestamp 1649977179
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_41
timestamp 1649977179
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_53
timestamp 1649977179
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_65
timestamp 1649977179
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1649977179
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1649977179
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_85
timestamp 1649977179
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_97
timestamp 1649977179
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_109
timestamp 1649977179
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_121
timestamp 1649977179
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1649977179
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1649977179
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_141
timestamp 1649977179
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_153
timestamp 1649977179
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_165
timestamp 1649977179
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_177
timestamp 1649977179
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_189
timestamp 1649977179
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_195
timestamp 1649977179
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_197
timestamp 1649977179
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_209
timestamp 1649977179
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_221
timestamp 1649977179
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_233
timestamp 1649977179
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1649977179
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1649977179
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_253
timestamp 1649977179
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_265
timestamp 1649977179
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_277
timestamp 1649977179
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_289
timestamp 1649977179
transform 1 0 27692 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_301
timestamp 1649977179
transform 1 0 28796 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_307
timestamp 1649977179
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_309
timestamp 1649977179
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_321
timestamp 1649977179
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_333
timestamp 1649977179
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_345
timestamp 1649977179
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_357
timestamp 1649977179
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_363
timestamp 1649977179
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_20_365
timestamp 1649977179
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_377
timestamp 1649977179
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_20_389
timestamp 1649977179
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_401
timestamp 1649977179
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_21_3
timestamp 1649977179
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_15
timestamp 1649977179
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_27
timestamp 1649977179
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_39
timestamp 1649977179
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_51
timestamp 1649977179
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1649977179
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_57
timestamp 1649977179
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_69
timestamp 1649977179
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_81
timestamp 1649977179
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_93
timestamp 1649977179
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1649977179
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1649977179
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_113
timestamp 1649977179
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_125
timestamp 1649977179
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_137
timestamp 1649977179
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_149
timestamp 1649977179
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1649977179
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1649977179
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_169
timestamp 1649977179
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_181
timestamp 1649977179
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_193
timestamp 1649977179
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_205
timestamp 1649977179
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_217
timestamp 1649977179
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1649977179
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_225
timestamp 1649977179
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_237
timestamp 1649977179
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_249
timestamp 1649977179
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_261
timestamp 1649977179
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_273
timestamp 1649977179
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_279
timestamp 1649977179
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_281
timestamp 1649977179
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_293
timestamp 1649977179
transform 1 0 28060 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_305
timestamp 1649977179
transform 1 0 29164 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_317
timestamp 1649977179
transform 1 0 30268 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_329
timestamp 1649977179
transform 1 0 31372 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_335
timestamp 1649977179
transform 1 0 31924 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_337
timestamp 1649977179
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_349
timestamp 1649977179
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_361
timestamp 1649977179
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_21_373
timestamp 1649977179
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_385
timestamp 1649977179
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_391
timestamp 1649977179
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_21_393
timestamp 1649977179
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_405
timestamp 1649977179
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_22_3
timestamp 1649977179
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_15
timestamp 1649977179
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1649977179
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_29
timestamp 1649977179
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_41
timestamp 1649977179
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_53
timestamp 1649977179
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_65
timestamp 1649977179
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1649977179
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1649977179
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_85
timestamp 1649977179
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_97
timestamp 1649977179
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_109
timestamp 1649977179
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_121
timestamp 1649977179
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1649977179
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1649977179
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_141
timestamp 1649977179
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_153
timestamp 1649977179
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_165
timestamp 1649977179
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_177
timestamp 1649977179
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1649977179
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1649977179
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_197
timestamp 1649977179
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_209
timestamp 1649977179
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_221
timestamp 1649977179
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_233
timestamp 1649977179
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_245
timestamp 1649977179
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1649977179
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_253
timestamp 1649977179
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_265
timestamp 1649977179
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_277
timestamp 1649977179
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_289
timestamp 1649977179
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_301
timestamp 1649977179
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1649977179
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_309
timestamp 1649977179
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_321
timestamp 1649977179
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_333
timestamp 1649977179
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_345
timestamp 1649977179
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_357
timestamp 1649977179
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1649977179
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_22_365
timestamp 1649977179
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_377
timestamp 1649977179
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_22_389
timestamp 1649977179
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_401
timestamp 1649977179
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_23_3
timestamp 1649977179
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_15
timestamp 1649977179
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_27
timestamp 1649977179
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_39
timestamp 1649977179
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1649977179
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1649977179
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_57
timestamp 1649977179
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_69
timestamp 1649977179
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_81
timestamp 1649977179
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_93
timestamp 1649977179
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_105
timestamp 1649977179
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1649977179
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_113
timestamp 1649977179
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_125
timestamp 1649977179
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_137
timestamp 1649977179
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_149
timestamp 1649977179
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1649977179
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1649977179
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_169
timestamp 1649977179
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_181
timestamp 1649977179
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_193
timestamp 1649977179
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_205
timestamp 1649977179
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_217
timestamp 1649977179
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1649977179
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_225
timestamp 1649977179
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_237
timestamp 1649977179
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_249
timestamp 1649977179
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_261
timestamp 1649977179
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_273
timestamp 1649977179
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_279
timestamp 1649977179
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_281
timestamp 1649977179
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_293
timestamp 1649977179
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_305
timestamp 1649977179
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_317
timestamp 1649977179
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_329
timestamp 1649977179
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1649977179
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_337
timestamp 1649977179
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_349
timestamp 1649977179
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_361
timestamp 1649977179
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_23_373
timestamp 1649977179
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_385
timestamp 1649977179
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_391
timestamp 1649977179
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_23_393
timestamp 1649977179
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_405
timestamp 1649977179
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_24_3
timestamp 1649977179
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_15
timestamp 1649977179
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1649977179
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_29
timestamp 1649977179
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_41
timestamp 1649977179
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_53
timestamp 1649977179
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_65
timestamp 1649977179
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1649977179
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1649977179
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_85
timestamp 1649977179
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_97
timestamp 1649977179
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_109
timestamp 1649977179
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_121
timestamp 1649977179
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_133
timestamp 1649977179
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_139
timestamp 1649977179
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_141
timestamp 1649977179
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_153
timestamp 1649977179
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_165
timestamp 1649977179
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_177
timestamp 1649977179
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_189
timestamp 1649977179
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_195
timestamp 1649977179
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_197
timestamp 1649977179
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_209
timestamp 1649977179
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_221
timestamp 1649977179
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_233
timestamp 1649977179
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_245
timestamp 1649977179
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1649977179
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_253
timestamp 1649977179
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_265
timestamp 1649977179
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_277
timestamp 1649977179
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_289
timestamp 1649977179
transform 1 0 27692 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1649977179
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1649977179
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_309
timestamp 1649977179
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_321
timestamp 1649977179
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_333
timestamp 1649977179
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_345
timestamp 1649977179
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_357
timestamp 1649977179
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_363
timestamp 1649977179
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_24_365
timestamp 1649977179
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_377
timestamp 1649977179
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_24_389
timestamp 1649977179
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_401
timestamp 1649977179
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_25_3
timestamp 1649977179
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_15
timestamp 1649977179
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_27
timestamp 1649977179
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_39
timestamp 1649977179
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1649977179
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1649977179
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_57
timestamp 1649977179
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_69
timestamp 1649977179
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_81
timestamp 1649977179
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_93
timestamp 1649977179
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1649977179
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1649977179
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_113
timestamp 1649977179
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_125
timestamp 1649977179
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_137
timestamp 1649977179
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_149
timestamp 1649977179
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_161
timestamp 1649977179
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_167
timestamp 1649977179
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_169
timestamp 1649977179
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_181
timestamp 1649977179
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_193
timestamp 1649977179
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_205
timestamp 1649977179
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_217
timestamp 1649977179
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_223
timestamp 1649977179
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_225
timestamp 1649977179
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_237
timestamp 1649977179
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_249
timestamp 1649977179
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_261
timestamp 1649977179
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_273
timestamp 1649977179
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1649977179
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_281
timestamp 1649977179
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_293
timestamp 1649977179
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_305
timestamp 1649977179
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_317
timestamp 1649977179
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_329
timestamp 1649977179
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_335
timestamp 1649977179
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_337
timestamp 1649977179
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_349
timestamp 1649977179
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_361
timestamp 1649977179
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_25_373
timestamp 1649977179
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_385
timestamp 1649977179
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1649977179
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_25_393
timestamp 1649977179
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_405
timestamp 1649977179
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_26_3
timestamp 1649977179
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_15
timestamp 1649977179
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_26_27
timestamp 1649977179
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_29
timestamp 1649977179
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_41
timestamp 1649977179
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_53
timestamp 1649977179
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_65
timestamp 1649977179
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_77
timestamp 1649977179
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1649977179
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_85
timestamp 1649977179
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_97
timestamp 1649977179
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_109
timestamp 1649977179
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_121
timestamp 1649977179
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_133
timestamp 1649977179
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_139
timestamp 1649977179
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_141
timestamp 1649977179
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_153
timestamp 1649977179
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_165
timestamp 1649977179
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_177
timestamp 1649977179
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_189
timestamp 1649977179
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_195
timestamp 1649977179
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_197
timestamp 1649977179
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_209
timestamp 1649977179
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_221
timestamp 1649977179
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_233
timestamp 1649977179
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_245
timestamp 1649977179
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_251
timestamp 1649977179
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_253
timestamp 1649977179
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_265
timestamp 1649977179
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_277
timestamp 1649977179
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_289
timestamp 1649977179
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_301
timestamp 1649977179
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_307
timestamp 1649977179
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_309
timestamp 1649977179
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_321
timestamp 1649977179
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_333
timestamp 1649977179
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_345
timestamp 1649977179
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_357
timestamp 1649977179
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_363
timestamp 1649977179
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_26_365
timestamp 1649977179
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_377
timestamp 1649977179
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_26_389
timestamp 1649977179
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_401
timestamp 1649977179
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_27_3
timestamp 1649977179
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_15
timestamp 1649977179
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_27
timestamp 1649977179
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_39
timestamp 1649977179
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_51
timestamp 1649977179
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1649977179
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_57
timestamp 1649977179
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_69
timestamp 1649977179
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_81
timestamp 1649977179
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_93
timestamp 1649977179
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_105
timestamp 1649977179
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_111
timestamp 1649977179
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_113
timestamp 1649977179
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_125
timestamp 1649977179
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_137
timestamp 1649977179
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_149
timestamp 1649977179
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_161
timestamp 1649977179
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1649977179
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_169
timestamp 1649977179
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_181
timestamp 1649977179
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_193
timestamp 1649977179
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_205
timestamp 1649977179
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_217
timestamp 1649977179
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_223
timestamp 1649977179
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_225
timestamp 1649977179
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_237
timestamp 1649977179
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_249
timestamp 1649977179
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_261
timestamp 1649977179
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1649977179
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1649977179
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_281
timestamp 1649977179
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_293
timestamp 1649977179
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_305
timestamp 1649977179
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_317
timestamp 1649977179
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_329
timestamp 1649977179
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1649977179
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_337
timestamp 1649977179
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_349
timestamp 1649977179
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_361
timestamp 1649977179
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_27_373
timestamp 1649977179
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_385
timestamp 1649977179
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_391
timestamp 1649977179
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_27_393
timestamp 1649977179
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_405
timestamp 1649977179
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_28_3
timestamp 1649977179
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_15
timestamp 1649977179
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1649977179
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_29
timestamp 1649977179
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_41
timestamp 1649977179
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_53
timestamp 1649977179
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_65
timestamp 1649977179
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_77
timestamp 1649977179
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_83
timestamp 1649977179
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_85
timestamp 1649977179
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_97
timestamp 1649977179
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_109
timestamp 1649977179
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_121
timestamp 1649977179
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_133
timestamp 1649977179
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_139
timestamp 1649977179
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_141
timestamp 1649977179
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_153
timestamp 1649977179
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_165
timestamp 1649977179
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_177
timestamp 1649977179
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1649977179
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1649977179
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_197
timestamp 1649977179
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_209
timestamp 1649977179
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_221
timestamp 1649977179
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_233
timestamp 1649977179
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_245
timestamp 1649977179
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_251
timestamp 1649977179
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_253
timestamp 1649977179
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_265
timestamp 1649977179
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_277
timestamp 1649977179
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_289
timestamp 1649977179
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1649977179
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1649977179
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_309
timestamp 1649977179
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_321
timestamp 1649977179
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_333
timestamp 1649977179
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_345
timestamp 1649977179
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_357
timestamp 1649977179
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1649977179
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_28_365
timestamp 1649977179
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_377
timestamp 1649977179
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_28_389
timestamp 1649977179
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_401
timestamp 1649977179
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_6
timestamp 1649977179
transform 1 0 1656 0 -1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_29_12
timestamp 1649977179
transform 1 0 2208 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_24
timestamp 1649977179
transform 1 0 3312 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_36
timestamp 1649977179
transform 1 0 4416 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_48
timestamp 1649977179
transform 1 0 5520 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_29_57
timestamp 1649977179
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_69
timestamp 1649977179
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_81
timestamp 1649977179
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_93
timestamp 1649977179
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_105
timestamp 1649977179
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_111
timestamp 1649977179
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_113
timestamp 1649977179
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_125
timestamp 1649977179
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_137
timestamp 1649977179
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_149
timestamp 1649977179
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_161
timestamp 1649977179
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1649977179
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_169
timestamp 1649977179
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_181
timestamp 1649977179
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_193
timestamp 1649977179
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_205
timestamp 1649977179
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_217
timestamp 1649977179
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_223
timestamp 1649977179
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_225
timestamp 1649977179
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_237
timestamp 1649977179
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_249
timestamp 1649977179
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_261
timestamp 1649977179
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_273
timestamp 1649977179
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1649977179
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_281
timestamp 1649977179
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_293
timestamp 1649977179
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_305
timestamp 1649977179
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_317
timestamp 1649977179
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_329
timestamp 1649977179
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_335
timestamp 1649977179
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_337
timestamp 1649977179
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_349
timestamp 1649977179
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_361
timestamp 1649977179
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_29_373
timestamp 1649977179
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1649977179
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1649977179
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_29_393
timestamp 1649977179
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_405
timestamp 1649977179
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_30_3
timestamp 1649977179
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_15
timestamp 1649977179
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1649977179
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_29
timestamp 1649977179
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_41
timestamp 1649977179
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_53
timestamp 1649977179
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_65
timestamp 1649977179
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_77
timestamp 1649977179
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1649977179
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_85
timestamp 1649977179
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_97
timestamp 1649977179
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_109
timestamp 1649977179
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_121
timestamp 1649977179
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_133
timestamp 1649977179
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1649977179
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_141
timestamp 1649977179
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_153
timestamp 1649977179
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_165
timestamp 1649977179
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_177
timestamp 1649977179
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_189
timestamp 1649977179
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1649977179
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_197
timestamp 1649977179
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_209
timestamp 1649977179
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_221
timestamp 1649977179
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_233
timestamp 1649977179
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_245
timestamp 1649977179
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_251
timestamp 1649977179
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_253
timestamp 1649977179
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_265
timestamp 1649977179
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_277
timestamp 1649977179
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_289
timestamp 1649977179
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_301
timestamp 1649977179
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_307
timestamp 1649977179
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_309
timestamp 1649977179
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_321
timestamp 1649977179
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_333
timestamp 1649977179
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_345
timestamp 1649977179
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_357
timestamp 1649977179
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1649977179
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_30_365
timestamp 1649977179
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_377
timestamp 1649977179
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_30_389
timestamp 1649977179
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_401
timestamp 1649977179
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_31_3
timestamp 1649977179
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_15
timestamp 1649977179
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_27
timestamp 1649977179
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_39
timestamp 1649977179
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1649977179
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1649977179
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_57
timestamp 1649977179
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_69
timestamp 1649977179
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_81
timestamp 1649977179
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_93
timestamp 1649977179
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_105
timestamp 1649977179
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_111
timestamp 1649977179
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_113
timestamp 1649977179
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_125
timestamp 1649977179
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_137
timestamp 1649977179
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_149
timestamp 1649977179
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_161
timestamp 1649977179
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_167
timestamp 1649977179
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_169
timestamp 1649977179
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_181
timestamp 1649977179
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_193
timestamp 1649977179
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_205
timestamp 1649977179
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_217
timestamp 1649977179
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_223
timestamp 1649977179
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_225
timestamp 1649977179
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_237
timestamp 1649977179
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_249
timestamp 1649977179
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_261
timestamp 1649977179
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_273
timestamp 1649977179
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_279
timestamp 1649977179
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_281
timestamp 1649977179
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_293
timestamp 1649977179
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_305
timestamp 1649977179
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_317
timestamp 1649977179
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_329
timestamp 1649977179
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_335
timestamp 1649977179
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_337
timestamp 1649977179
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_349
timestamp 1649977179
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_361
timestamp 1649977179
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_31_373
timestamp 1649977179
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_385
timestamp 1649977179
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1649977179
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_31_393
timestamp 1649977179
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_405
timestamp 1649977179
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_32_3
timestamp 1649977179
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_15
timestamp 1649977179
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1649977179
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_29
timestamp 1649977179
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_41
timestamp 1649977179
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_53
timestamp 1649977179
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_65
timestamp 1649977179
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1649977179
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1649977179
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_85
timestamp 1649977179
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_97
timestamp 1649977179
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_109
timestamp 1649977179
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_121
timestamp 1649977179
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_133
timestamp 1649977179
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_139
timestamp 1649977179
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_141
timestamp 1649977179
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_153
timestamp 1649977179
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_165
timestamp 1649977179
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_177
timestamp 1649977179
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_189
timestamp 1649977179
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_195
timestamp 1649977179
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_197
timestamp 1649977179
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_209
timestamp 1649977179
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_221
timestamp 1649977179
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_233
timestamp 1649977179
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_245
timestamp 1649977179
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1649977179
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_253
timestamp 1649977179
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_265
timestamp 1649977179
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_277
timestamp 1649977179
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_289
timestamp 1649977179
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_301
timestamp 1649977179
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_307
timestamp 1649977179
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_309
timestamp 1649977179
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_321
timestamp 1649977179
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_333
timestamp 1649977179
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_345
timestamp 1649977179
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_357
timestamp 1649977179
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1649977179
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_32_365
timestamp 1649977179
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_377
timestamp 1649977179
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_32_389
timestamp 1649977179
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_401
timestamp 1649977179
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_33_3
timestamp 1649977179
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_15
timestamp 1649977179
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_27
timestamp 1649977179
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_39
timestamp 1649977179
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1649977179
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1649977179
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_57
timestamp 1649977179
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_69
timestamp 1649977179
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_81
timestamp 1649977179
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_93
timestamp 1649977179
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_105
timestamp 1649977179
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_111
timestamp 1649977179
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_113
timestamp 1649977179
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_125
timestamp 1649977179
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_137
timestamp 1649977179
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_149
timestamp 1649977179
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_161
timestamp 1649977179
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1649977179
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_169
timestamp 1649977179
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_181
timestamp 1649977179
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_193
timestamp 1649977179
transform 1 0 18860 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_198
timestamp 1649977179
transform 1 0 19320 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_206
timestamp 1649977179
transform 1 0 20056 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_211
timestamp 1649977179
transform 1 0 20516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_223
timestamp 1649977179
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_227
timestamp 1649977179
transform 1 0 21988 0 -1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_33_233
timestamp 1649977179
transform 1 0 22540 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_245
timestamp 1649977179
transform 1 0 23644 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_257
timestamp 1649977179
transform 1 0 24748 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_269
timestamp 1649977179
transform 1 0 25852 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_277
timestamp 1649977179
transform 1 0 26588 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_33_281
timestamp 1649977179
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_293
timestamp 1649977179
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_305
timestamp 1649977179
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_317
timestamp 1649977179
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_329
timestamp 1649977179
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_335
timestamp 1649977179
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_337
timestamp 1649977179
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_349
timestamp 1649977179
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_361
timestamp 1649977179
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_33_373
timestamp 1649977179
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_385
timestamp 1649977179
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_391
timestamp 1649977179
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_33_393
timestamp 1649977179
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_405
timestamp 1649977179
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_34_3
timestamp 1649977179
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_15
timestamp 1649977179
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1649977179
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_29
timestamp 1649977179
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_41
timestamp 1649977179
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_53
timestamp 1649977179
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_65
timestamp 1649977179
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1649977179
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1649977179
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_85
timestamp 1649977179
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_97
timestamp 1649977179
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_109
timestamp 1649977179
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_121
timestamp 1649977179
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1649977179
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1649977179
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_141
timestamp 1649977179
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_153
timestamp 1649977179
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_165
timestamp 1649977179
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_177
timestamp 1649977179
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_189
timestamp 1649977179
transform 1 0 18492 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1649977179
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_197
timestamp 1649977179
transform 1 0 19228 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_205
timestamp 1649977179
transform 1 0 19964 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_213
timestamp 1649977179
transform 1 0 20700 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_224
timestamp 1649977179
transform 1 0 21712 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_231
timestamp 1649977179
transform 1 0 22356 0 1 20672
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_34_237
timestamp 1649977179
transform 1 0 22908 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_249
timestamp 1649977179
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_34_253
timestamp 1649977179
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_265
timestamp 1649977179
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_277
timestamp 1649977179
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_289
timestamp 1649977179
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1649977179
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1649977179
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_309
timestamp 1649977179
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_321
timestamp 1649977179
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_333
timestamp 1649977179
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_345
timestamp 1649977179
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_357
timestamp 1649977179
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_363
timestamp 1649977179
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_34_365
timestamp 1649977179
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_377
timestamp 1649977179
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_34_389
timestamp 1649977179
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_401
timestamp 1649977179
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_35_3
timestamp 1649977179
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_15
timestamp 1649977179
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_27
timestamp 1649977179
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_39
timestamp 1649977179
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1649977179
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1649977179
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_57
timestamp 1649977179
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_69
timestamp 1649977179
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_81
timestamp 1649977179
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_93
timestamp 1649977179
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_105
timestamp 1649977179
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1649977179
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_113
timestamp 1649977179
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_125
timestamp 1649977179
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_137
timestamp 1649977179
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_149
timestamp 1649977179
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_161
timestamp 1649977179
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1649977179
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_169
timestamp 1649977179
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_181
timestamp 1649977179
transform 1 0 17756 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_187
timestamp 1649977179
transform 1 0 18308 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_193
timestamp 1649977179
transform 1 0 18860 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_201
timestamp 1649977179
transform 1 0 19596 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_209
timestamp 1649977179
transform 1 0 20332 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_219
timestamp 1649977179
transform 1 0 21252 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_223
timestamp 1649977179
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_242
timestamp 1649977179
transform 1 0 23368 0 -1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_35_248
timestamp 1649977179
transform 1 0 23920 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_260
timestamp 1649977179
transform 1 0 25024 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_272
timestamp 1649977179
transform 1 0 26128 0 -1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_35_281
timestamp 1649977179
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_293
timestamp 1649977179
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_305
timestamp 1649977179
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_317
timestamp 1649977179
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_329
timestamp 1649977179
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_335
timestamp 1649977179
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_337
timestamp 1649977179
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_349
timestamp 1649977179
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_361
timestamp 1649977179
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_35_373
timestamp 1649977179
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_385
timestamp 1649977179
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1649977179
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_35_393
timestamp 1649977179
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_405
timestamp 1649977179
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_36_3
timestamp 1649977179
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_15
timestamp 1649977179
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1649977179
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_29
timestamp 1649977179
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_41
timestamp 1649977179
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_53
timestamp 1649977179
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_65
timestamp 1649977179
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1649977179
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1649977179
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_85
timestamp 1649977179
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_97
timestamp 1649977179
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_109
timestamp 1649977179
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_121
timestamp 1649977179
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_133
timestamp 1649977179
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1649977179
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_141
timestamp 1649977179
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_153
timestamp 1649977179
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_165
timestamp 1649977179
transform 1 0 16284 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_36_170
timestamp 1649977179
transform 1 0 16744 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_36_185
timestamp 1649977179
transform 1 0 18124 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_189
timestamp 1649977179
transform 1 0 18492 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1649977179
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_197
timestamp 1649977179
transform 1 0 19228 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_201
timestamp 1649977179
transform 1 0 19596 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_216
timestamp 1649977179
transform 1 0 20976 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_222
timestamp 1649977179
transform 1 0 21528 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_230
timestamp 1649977179
transform 1 0 22264 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_237
timestamp 1649977179
transform 1 0 22908 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_244
timestamp 1649977179
transform 1 0 23552 0 1 21760
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_36_253
timestamp 1649977179
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_265
timestamp 1649977179
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_277
timestamp 1649977179
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_289
timestamp 1649977179
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_301
timestamp 1649977179
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_307
timestamp 1649977179
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_309
timestamp 1649977179
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_321
timestamp 1649977179
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_333
timestamp 1649977179
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_345
timestamp 1649977179
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_357
timestamp 1649977179
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_363
timestamp 1649977179
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_36_365
timestamp 1649977179
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_377
timestamp 1649977179
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_36_389
timestamp 1649977179
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_401
timestamp 1649977179
transform 1 0 37996 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_37_3
timestamp 1649977179
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_15
timestamp 1649977179
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_27
timestamp 1649977179
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_39
timestamp 1649977179
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_51
timestamp 1649977179
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_55
timestamp 1649977179
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_57
timestamp 1649977179
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_69
timestamp 1649977179
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_81
timestamp 1649977179
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_93
timestamp 1649977179
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1649977179
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1649977179
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_113
timestamp 1649977179
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_125
timestamp 1649977179
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_137
timestamp 1649977179
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_152
timestamp 1649977179
transform 1 0 15088 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_161
timestamp 1649977179
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_167
timestamp 1649977179
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_169
timestamp 1649977179
transform 1 0 16652 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_178
timestamp 1649977179
transform 1 0 17480 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_189
timestamp 1649977179
transform 1 0 18492 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_199
timestamp 1649977179
transform 1 0 19412 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_209
timestamp 1649977179
transform 1 0 20332 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1649977179
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_231
timestamp 1649977179
transform 1 0 22356 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_237
timestamp 1649977179
transform 1 0 22908 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_243
timestamp 1649977179
transform 1 0 23460 0 -1 22848
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_37_249
timestamp 1649977179
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_261
timestamp 1649977179
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_273
timestamp 1649977179
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1649977179
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_281
timestamp 1649977179
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_293
timestamp 1649977179
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_305
timestamp 1649977179
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_317
timestamp 1649977179
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_329
timestamp 1649977179
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1649977179
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_337
timestamp 1649977179
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_349
timestamp 1649977179
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_361
timestamp 1649977179
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_37_373
timestamp 1649977179
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_385
timestamp 1649977179
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1649977179
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_37_393
timestamp 1649977179
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_405
timestamp 1649977179
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_38_3
timestamp 1649977179
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_15
timestamp 1649977179
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1649977179
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_29
timestamp 1649977179
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_41
timestamp 1649977179
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_53
timestamp 1649977179
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_65
timestamp 1649977179
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_77
timestamp 1649977179
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1649977179
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_85
timestamp 1649977179
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_97
timestamp 1649977179
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_109
timestamp 1649977179
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_121
timestamp 1649977179
transform 1 0 12236 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_127
timestamp 1649977179
transform 1 0 12788 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_135
timestamp 1649977179
transform 1 0 13524 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_139
timestamp 1649977179
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_141
timestamp 1649977179
transform 1 0 14076 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_149
timestamp 1649977179
transform 1 0 14812 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_155
timestamp 1649977179
transform 1 0 15364 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_166
timestamp 1649977179
transform 1 0 16376 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_177
timestamp 1649977179
transform 1 0 17388 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_186
timestamp 1649977179
transform 1 0 18216 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_192
timestamp 1649977179
transform 1 0 18768 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_203
timestamp 1649977179
transform 1 0 19780 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_214
timestamp 1649977179
transform 1 0 20792 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_225
timestamp 1649977179
transform 1 0 21804 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_231
timestamp 1649977179
transform 1 0 22356 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_241
timestamp 1649977179
transform 1 0 23276 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_247
timestamp 1649977179
transform 1 0 23828 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_251
timestamp 1649977179
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_255
timestamp 1649977179
transform 1 0 24564 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_267
timestamp 1649977179
transform 1 0 25668 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_279
timestamp 1649977179
transform 1 0 26772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_291
timestamp 1649977179
transform 1 0 27876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_303
timestamp 1649977179
transform 1 0 28980 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_307
timestamp 1649977179
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_309
timestamp 1649977179
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_321
timestamp 1649977179
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_333
timestamp 1649977179
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_345
timestamp 1649977179
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_357
timestamp 1649977179
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_363
timestamp 1649977179
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_38_365
timestamp 1649977179
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_377
timestamp 1649977179
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_38_389
timestamp 1649977179
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_401
timestamp 1649977179
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_39_3
timestamp 1649977179
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_15
timestamp 1649977179
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_27
timestamp 1649977179
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_39
timestamp 1649977179
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_51
timestamp 1649977179
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1649977179
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_57
timestamp 1649977179
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_69
timestamp 1649977179
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_81
timestamp 1649977179
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_93
timestamp 1649977179
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_105
timestamp 1649977179
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1649977179
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_113
timestamp 1649977179
transform 1 0 11500 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_121
timestamp 1649977179
transform 1 0 12236 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_125
timestamp 1649977179
transform 1 0 12604 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_133
timestamp 1649977179
transform 1 0 13340 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_142
timestamp 1649977179
transform 1 0 14168 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_148
timestamp 1649977179
transform 1 0 14720 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_155
timestamp 1649977179
transform 1 0 15364 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1649977179
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1649977179
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_173
timestamp 1649977179
transform 1 0 17020 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_182
timestamp 1649977179
transform 1 0 17848 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_206
timestamp 1649977179
transform 1 0 20056 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_212
timestamp 1649977179
transform 1 0 20608 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_220
timestamp 1649977179
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_235
timestamp 1649977179
transform 1 0 22724 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_246
timestamp 1649977179
transform 1 0 23736 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_39_256
timestamp 1649977179
transform 1 0 24656 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_268
timestamp 1649977179
transform 1 0 25760 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_281
timestamp 1649977179
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_293
timestamp 1649977179
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_305
timestamp 1649977179
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_317
timestamp 1649977179
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1649977179
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1649977179
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_337
timestamp 1649977179
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_349
timestamp 1649977179
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_361
timestamp 1649977179
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_39_373
timestamp 1649977179
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_385
timestamp 1649977179
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_391
timestamp 1649977179
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_39_393
timestamp 1649977179
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_405
timestamp 1649977179
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_40_3
timestamp 1649977179
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_15
timestamp 1649977179
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1649977179
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_29
timestamp 1649977179
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_41
timestamp 1649977179
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_53
timestamp 1649977179
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_65
timestamp 1649977179
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1649977179
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1649977179
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_85
timestamp 1649977179
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_97
timestamp 1649977179
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_109
timestamp 1649977179
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_121
timestamp 1649977179
transform 1 0 12236 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_124
timestamp 1649977179
transform 1 0 12512 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1649977179
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_148
timestamp 1649977179
transform 1 0 14720 0 1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_40_154
timestamp 1649977179
transform 1 0 15272 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_166
timestamp 1649977179
transform 1 0 16376 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_170
timestamp 1649977179
transform 1 0 16744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_176
timestamp 1649977179
transform 1 0 17296 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_184
timestamp 1649977179
transform 1 0 18032 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_191
timestamp 1649977179
transform 1 0 18676 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1649977179
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_199
timestamp 1649977179
transform 1 0 19412 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_209
timestamp 1649977179
transform 1 0 20332 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_215
timestamp 1649977179
transform 1 0 20884 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_221
timestamp 1649977179
transform 1 0 21436 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_224
timestamp 1649977179
transform 1 0 21712 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_234
timestamp 1649977179
transform 1 0 22632 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_40_245
timestamp 1649977179
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1649977179
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_255
timestamp 1649977179
transform 1 0 24564 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_267
timestamp 1649977179
transform 1 0 25668 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_279
timestamp 1649977179
transform 1 0 26772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_291
timestamp 1649977179
transform 1 0 27876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_303
timestamp 1649977179
transform 1 0 28980 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_307
timestamp 1649977179
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_309
timestamp 1649977179
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_321
timestamp 1649977179
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_333
timestamp 1649977179
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_345
timestamp 1649977179
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1649977179
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1649977179
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_40_365
timestamp 1649977179
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_377
timestamp 1649977179
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_40_389
timestamp 1649977179
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_401
timestamp 1649977179
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_41_3
timestamp 1649977179
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_15
timestamp 1649977179
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_27
timestamp 1649977179
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_39
timestamp 1649977179
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1649977179
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1649977179
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_57
timestamp 1649977179
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_69
timestamp 1649977179
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_81
timestamp 1649977179
transform 1 0 8556 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_89
timestamp 1649977179
transform 1 0 9292 0 -1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_41_94
timestamp 1649977179
transform 1 0 9752 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_106
timestamp 1649977179
transform 1 0 10856 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_41_113
timestamp 1649977179
transform 1 0 11500 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_117
timestamp 1649977179
transform 1 0 11868 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_127
timestamp 1649977179
transform 1 0 12788 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_140
timestamp 1649977179
transform 1 0 13984 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_146
timestamp 1649977179
transform 1 0 14536 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_158
timestamp 1649977179
transform 1 0 15640 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_166
timestamp 1649977179
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_186
timestamp 1649977179
transform 1 0 18216 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_192
timestamp 1649977179
transform 1 0 18768 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_195
timestamp 1649977179
transform 1 0 19044 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_203
timestamp 1649977179
transform 1 0 19780 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_220
timestamp 1649977179
transform 1 0 21344 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_225
timestamp 1649977179
transform 1 0 21804 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_228
timestamp 1649977179
transform 1 0 22080 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_236
timestamp 1649977179
transform 1 0 22816 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_239
timestamp 1649977179
transform 1 0 23092 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_247
timestamp 1649977179
transform 1 0 23828 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_41_254
timestamp 1649977179
transform 1 0 24472 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_266
timestamp 1649977179
transform 1 0 25576 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_278
timestamp 1649977179
transform 1 0 26680 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_41_281
timestamp 1649977179
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_293
timestamp 1649977179
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_305
timestamp 1649977179
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_317
timestamp 1649977179
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_329
timestamp 1649977179
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_335
timestamp 1649977179
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_337
timestamp 1649977179
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_349
timestamp 1649977179
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_361
timestamp 1649977179
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_41_373
timestamp 1649977179
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_385
timestamp 1649977179
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_391
timestamp 1649977179
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_41_393
timestamp 1649977179
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_405
timestamp 1649977179
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_3
timestamp 1649977179
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_15
timestamp 1649977179
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1649977179
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_29
timestamp 1649977179
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_41
timestamp 1649977179
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_53
timestamp 1649977179
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_65
timestamp 1649977179
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_77
timestamp 1649977179
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_83
timestamp 1649977179
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_85
timestamp 1649977179
transform 1 0 8924 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_42_92
timestamp 1649977179
transform 1 0 9568 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_100
timestamp 1649977179
transform 1 0 10304 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_105
timestamp 1649977179
transform 1 0 10764 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_111
timestamp 1649977179
transform 1 0 11316 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_116
timestamp 1649977179
transform 1 0 11776 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_122
timestamp 1649977179
transform 1 0 12328 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_125
timestamp 1649977179
transform 1 0 12604 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_133
timestamp 1649977179
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_139
timestamp 1649977179
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_141
timestamp 1649977179
transform 1 0 14076 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_145
timestamp 1649977179
transform 1 0 14444 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_153
timestamp 1649977179
transform 1 0 15180 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_177
timestamp 1649977179
transform 1 0 17388 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_190
timestamp 1649977179
transform 1 0 18584 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_197
timestamp 1649977179
transform 1 0 19228 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_206
timestamp 1649977179
transform 1 0 20056 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_217
timestamp 1649977179
transform 1 0 21068 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_223
timestamp 1649977179
transform 1 0 21620 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_226
timestamp 1649977179
transform 1 0 21896 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_238
timestamp 1649977179
transform 1 0 23000 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_250
timestamp 1649977179
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_42_253
timestamp 1649977179
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_265
timestamp 1649977179
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_277
timestamp 1649977179
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_289
timestamp 1649977179
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_301
timestamp 1649977179
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_307
timestamp 1649977179
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_309
timestamp 1649977179
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_321
timestamp 1649977179
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_333
timestamp 1649977179
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_345
timestamp 1649977179
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1649977179
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1649977179
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_42_365
timestamp 1649977179
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_377
timestamp 1649977179
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_42_389
timestamp 1649977179
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_401
timestamp 1649977179
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_43_3
timestamp 1649977179
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_15
timestamp 1649977179
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_27
timestamp 1649977179
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_39
timestamp 1649977179
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1649977179
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1649977179
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_57
timestamp 1649977179
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_69
timestamp 1649977179
transform 1 0 7452 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_74
timestamp 1649977179
transform 1 0 7912 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_43_95
timestamp 1649977179
transform 1 0 9844 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_107
timestamp 1649977179
transform 1 0 10948 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1649977179
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_43_113
timestamp 1649977179
transform 1 0 11500 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_130
timestamp 1649977179
transform 1 0 13064 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_136
timestamp 1649977179
transform 1 0 13616 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_143
timestamp 1649977179
transform 1 0 14260 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_147
timestamp 1649977179
transform 1 0 14628 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_164
timestamp 1649977179
transform 1 0 16192 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_169
timestamp 1649977179
transform 1 0 16652 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_175
timestamp 1649977179
transform 1 0 17204 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_201
timestamp 1649977179
transform 1 0 19596 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_207
timestamp 1649977179
transform 1 0 20148 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_211
timestamp 1649977179
transform 1 0 20516 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_214
timestamp 1649977179
transform 1 0 20792 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1649977179
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_225
timestamp 1649977179
transform 1 0 21804 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_232
timestamp 1649977179
transform 1 0 22448 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_244
timestamp 1649977179
transform 1 0 23552 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_256
timestamp 1649977179
transform 1 0 24656 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_268
timestamp 1649977179
transform 1 0 25760 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_281
timestamp 1649977179
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_293
timestamp 1649977179
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_305
timestamp 1649977179
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_317
timestamp 1649977179
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1649977179
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1649977179
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_337
timestamp 1649977179
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_349
timestamp 1649977179
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_361
timestamp 1649977179
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_43_373
timestamp 1649977179
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1649977179
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1649977179
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_43_393
timestamp 1649977179
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_405
timestamp 1649977179
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_19
timestamp 1649977179
transform 1 0 2852 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1649977179
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_48
timestamp 1649977179
transform 1 0 5520 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_60
timestamp 1649977179
transform 1 0 6624 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_72
timestamp 1649977179
transform 1 0 7728 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_89
timestamp 1649977179
transform 1 0 9292 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_96
timestamp 1649977179
transform 1 0 9936 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_102
timestamp 1649977179
transform 1 0 10488 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_110
timestamp 1649977179
transform 1 0 11224 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_113
timestamp 1649977179
transform 1 0 11500 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_123
timestamp 1649977179
transform 1 0 12420 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_129
timestamp 1649977179
transform 1 0 12972 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_133
timestamp 1649977179
transform 1 0 13340 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_136
timestamp 1649977179
transform 1 0 13616 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_141
timestamp 1649977179
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_153
timestamp 1649977179
transform 1 0 15180 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_157
timestamp 1649977179
transform 1 0 15548 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_178
timestamp 1649977179
transform 1 0 17480 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_191
timestamp 1649977179
transform 1 0 18676 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_195
timestamp 1649977179
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_44_197
timestamp 1649977179
transform 1 0 19228 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_203
timestamp 1649977179
transform 1 0 19780 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_213
timestamp 1649977179
transform 1 0 20700 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_219
timestamp 1649977179
transform 1 0 21252 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_230
timestamp 1649977179
transform 1 0 22264 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_44_238
timestamp 1649977179
transform 1 0 23000 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_250
timestamp 1649977179
transform 1 0 24104 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_44_253
timestamp 1649977179
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_265
timestamp 1649977179
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_277
timestamp 1649977179
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_289
timestamp 1649977179
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_301
timestamp 1649977179
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_307
timestamp 1649977179
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_309
timestamp 1649977179
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_321
timestamp 1649977179
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_333
timestamp 1649977179
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_345
timestamp 1649977179
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_357
timestamp 1649977179
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_363
timestamp 1649977179
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_44_365
timestamp 1649977179
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_377
timestamp 1649977179
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_44_389
timestamp 1649977179
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_401
timestamp 1649977179
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_45_3
timestamp 1649977179
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_15
timestamp 1649977179
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_27
timestamp 1649977179
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_39
timestamp 1649977179
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_51
timestamp 1649977179
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_55
timestamp 1649977179
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_57
timestamp 1649977179
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_69
timestamp 1649977179
transform 1 0 7452 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_45_87
timestamp 1649977179
transform 1 0 9108 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_45_101
timestamp 1649977179
transform 1 0 10396 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_109
timestamp 1649977179
transform 1 0 11132 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_118
timestamp 1649977179
transform 1 0 11960 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_125
timestamp 1649977179
transform 1 0 12604 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_131
timestamp 1649977179
transform 1 0 13156 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_139
timestamp 1649977179
transform 1 0 13892 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_45_143
timestamp 1649977179
transform 1 0 14260 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_149
timestamp 1649977179
transform 1 0 14812 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_153
timestamp 1649977179
transform 1 0 15180 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_160
timestamp 1649977179
transform 1 0 15824 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_185
timestamp 1649977179
transform 1 0 18124 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_197
timestamp 1649977179
transform 1 0 19228 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_208
timestamp 1649977179
transform 1 0 20240 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_220
timestamp 1649977179
transform 1 0 21344 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_229
timestamp 1649977179
transform 1 0 22172 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_45_235
timestamp 1649977179
transform 1 0 22724 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_247
timestamp 1649977179
transform 1 0 23828 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_259
timestamp 1649977179
transform 1 0 24932 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_271
timestamp 1649977179
transform 1 0 26036 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_279
timestamp 1649977179
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_281
timestamp 1649977179
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_293
timestamp 1649977179
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_305
timestamp 1649977179
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_317
timestamp 1649977179
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_329
timestamp 1649977179
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1649977179
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_337
timestamp 1649977179
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_349
timestamp 1649977179
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_361
timestamp 1649977179
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_45_373
timestamp 1649977179
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1649977179
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1649977179
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_45_393
timestamp 1649977179
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1649977179
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_20
timestamp 1649977179
transform 1 0 2944 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_46_29
timestamp 1649977179
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_41
timestamp 1649977179
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_53
timestamp 1649977179
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_65
timestamp 1649977179
transform 1 0 7084 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_46_72
timestamp 1649977179
transform 1 0 7728 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_94
timestamp 1649977179
transform 1 0 9752 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_104
timestamp 1649977179
transform 1 0 10672 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_117
timestamp 1649977179
transform 1 0 11868 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_123
timestamp 1649977179
transform 1 0 12420 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_130
timestamp 1649977179
transform 1 0 13064 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1649977179
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_143
timestamp 1649977179
transform 1 0 14260 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_151
timestamp 1649977179
transform 1 0 14996 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_46_155
timestamp 1649977179
transform 1 0 15364 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_177
timestamp 1649977179
transform 1 0 17388 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_183
timestamp 1649977179
transform 1 0 17940 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1649977179
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_197
timestamp 1649977179
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_201
timestamp 1649977179
transform 1 0 19596 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_208
timestamp 1649977179
transform 1 0 20240 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_218
timestamp 1649977179
transform 1 0 21160 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_222
timestamp 1649977179
transform 1 0 21528 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_225
timestamp 1649977179
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_237
timestamp 1649977179
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_249
timestamp 1649977179
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_46_253
timestamp 1649977179
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_265
timestamp 1649977179
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_277
timestamp 1649977179
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_289
timestamp 1649977179
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1649977179
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1649977179
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_309
timestamp 1649977179
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_321
timestamp 1649977179
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_333
timestamp 1649977179
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_345
timestamp 1649977179
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_357
timestamp 1649977179
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_363
timestamp 1649977179
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_46_365
timestamp 1649977179
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_377
timestamp 1649977179
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_46_389
timestamp 1649977179
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_401
timestamp 1649977179
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_47_3
timestamp 1649977179
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_32
timestamp 1649977179
transform 1 0 4048 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_44
timestamp 1649977179
transform 1 0 5152 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_57
timestamp 1649977179
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_69
timestamp 1649977179
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_81
timestamp 1649977179
transform 1 0 8556 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_87
timestamp 1649977179
transform 1 0 9108 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_90
timestamp 1649977179
transform 1 0 9384 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_97
timestamp 1649977179
transform 1 0 10028 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1649977179
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_113
timestamp 1649977179
transform 1 0 11500 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_117
timestamp 1649977179
transform 1 0 11868 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_137
timestamp 1649977179
transform 1 0 13708 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_47_148
timestamp 1649977179
transform 1 0 14720 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_157
timestamp 1649977179
transform 1 0 15548 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_165
timestamp 1649977179
transform 1 0 16284 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_47_169
timestamp 1649977179
transform 1 0 16652 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_177
timestamp 1649977179
transform 1 0 17388 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_180
timestamp 1649977179
transform 1 0 17664 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_189
timestamp 1649977179
transform 1 0 18492 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_196
timestamp 1649977179
transform 1 0 19136 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_207
timestamp 1649977179
transform 1 0 20148 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_213
timestamp 1649977179
transform 1 0 20700 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_219
timestamp 1649977179
transform 1 0 21252 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1649977179
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_225
timestamp 1649977179
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_237
timestamp 1649977179
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_249
timestamp 1649977179
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_261
timestamp 1649977179
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_273
timestamp 1649977179
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_279
timestamp 1649977179
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_281
timestamp 1649977179
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_293
timestamp 1649977179
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_305
timestamp 1649977179
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_317
timestamp 1649977179
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_329
timestamp 1649977179
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_335
timestamp 1649977179
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_337
timestamp 1649977179
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_349
timestamp 1649977179
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_361
timestamp 1649977179
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_47_373
timestamp 1649977179
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_385
timestamp 1649977179
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_391
timestamp 1649977179
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_47_393
timestamp 1649977179
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_405
timestamp 1649977179
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_48_3
timestamp 1649977179
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_15
timestamp 1649977179
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1649977179
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_29
timestamp 1649977179
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_41
timestamp 1649977179
transform 1 0 4876 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_65
timestamp 1649977179
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_77
timestamp 1649977179
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_83
timestamp 1649977179
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_85
timestamp 1649977179
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_93
timestamp 1649977179
transform 1 0 9660 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_97
timestamp 1649977179
transform 1 0 10028 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_121
timestamp 1649977179
transform 1 0 12236 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_48_128
timestamp 1649977179
transform 1 0 12880 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_141
timestamp 1649977179
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_153
timestamp 1649977179
transform 1 0 15180 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_159
timestamp 1649977179
transform 1 0 15732 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_176
timestamp 1649977179
transform 1 0 17296 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_188
timestamp 1649977179
transform 1 0 18400 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1649977179
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_201
timestamp 1649977179
transform 1 0 19596 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_48_209
timestamp 1649977179
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_221
timestamp 1649977179
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_233
timestamp 1649977179
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_245
timestamp 1649977179
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_251
timestamp 1649977179
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_253
timestamp 1649977179
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_265
timestamp 1649977179
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_277
timestamp 1649977179
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_289
timestamp 1649977179
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_301
timestamp 1649977179
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1649977179
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_309
timestamp 1649977179
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_321
timestamp 1649977179
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_333
timestamp 1649977179
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_345
timestamp 1649977179
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_357
timestamp 1649977179
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_363
timestamp 1649977179
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_48_365
timestamp 1649977179
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_377
timestamp 1649977179
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_48_389
timestamp 1649977179
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1649977179
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_49_3
timestamp 1649977179
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_15
timestamp 1649977179
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_27
timestamp 1649977179
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_39
timestamp 1649977179
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_51
timestamp 1649977179
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1649977179
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_57
timestamp 1649977179
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_85
timestamp 1649977179
transform 1 0 8924 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_97
timestamp 1649977179
transform 1 0 10028 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_105
timestamp 1649977179
transform 1 0 10764 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_108
timestamp 1649977179
transform 1 0 11040 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_119
timestamp 1649977179
transform 1 0 12052 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_125
timestamp 1649977179
transform 1 0 12604 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_145
timestamp 1649977179
transform 1 0 14444 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_153
timestamp 1649977179
transform 1 0 15180 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_158
timestamp 1649977179
transform 1 0 15640 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1649977179
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_49_169
timestamp 1649977179
transform 1 0 16652 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_49_176
timestamp 1649977179
transform 1 0 17296 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_188
timestamp 1649977179
transform 1 0 18400 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_194
timestamp 1649977179
transform 1 0 18952 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_199
timestamp 1649977179
transform 1 0 19412 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_49_205
timestamp 1649977179
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_217
timestamp 1649977179
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1649977179
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_225
timestamp 1649977179
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_237
timestamp 1649977179
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_249
timestamp 1649977179
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_261
timestamp 1649977179
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_273
timestamp 1649977179
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_279
timestamp 1649977179
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_281
timestamp 1649977179
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_293
timestamp 1649977179
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_305
timestamp 1649977179
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_317
timestamp 1649977179
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_329
timestamp 1649977179
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1649977179
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_337
timestamp 1649977179
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_349
timestamp 1649977179
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_361
timestamp 1649977179
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_49_373
timestamp 1649977179
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_385
timestamp 1649977179
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_391
timestamp 1649977179
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_49_393
timestamp 1649977179
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_405
timestamp 1649977179
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_50_3
timestamp 1649977179
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_15
timestamp 1649977179
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_27
timestamp 1649977179
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_29
timestamp 1649977179
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_41
timestamp 1649977179
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_53
timestamp 1649977179
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_65
timestamp 1649977179
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1649977179
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1649977179
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_85
timestamp 1649977179
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_97
timestamp 1649977179
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_111
timestamp 1649977179
transform 1 0 11316 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_123
timestamp 1649977179
transform 1 0 12420 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_135
timestamp 1649977179
transform 1 0 13524 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1649977179
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_141
timestamp 1649977179
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_159
timestamp 1649977179
transform 1 0 15732 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_165
timestamp 1649977179
transform 1 0 16284 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_171
timestamp 1649977179
transform 1 0 16836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_183
timestamp 1649977179
transform 1 0 17940 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_186
timestamp 1649977179
transform 1 0 18216 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1649977179
transform 1 0 18768 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_204
timestamp 1649977179
transform 1 0 19872 0 1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_50_210
timestamp 1649977179
transform 1 0 20424 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_222
timestamp 1649977179
transform 1 0 21528 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_234
timestamp 1649977179
transform 1 0 22632 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_246
timestamp 1649977179
transform 1 0 23736 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_50_253
timestamp 1649977179
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_265
timestamp 1649977179
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_277
timestamp 1649977179
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_289
timestamp 1649977179
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_301
timestamp 1649977179
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1649977179
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_309
timestamp 1649977179
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_321
timestamp 1649977179
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_333
timestamp 1649977179
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_345
timestamp 1649977179
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_357
timestamp 1649977179
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1649977179
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_50_365
timestamp 1649977179
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_377
timestamp 1649977179
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_50_389
timestamp 1649977179
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_401
timestamp 1649977179
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_51_3
timestamp 1649977179
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_15
timestamp 1649977179
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_27
timestamp 1649977179
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_39
timestamp 1649977179
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1649977179
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1649977179
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_57
timestamp 1649977179
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_69
timestamp 1649977179
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_81
timestamp 1649977179
transform 1 0 8556 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_87
timestamp 1649977179
transform 1 0 9108 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_90
timestamp 1649977179
transform 1 0 9384 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_102
timestamp 1649977179
transform 1 0 10488 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_110
timestamp 1649977179
transform 1 0 11224 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_51_113
timestamp 1649977179
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_125
timestamp 1649977179
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_137
timestamp 1649977179
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_149
timestamp 1649977179
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_161
timestamp 1649977179
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_167
timestamp 1649977179
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_185
timestamp 1649977179
transform 1 0 18124 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_199
timestamp 1649977179
transform 1 0 19412 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_51_205
timestamp 1649977179
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1649977179
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1649977179
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_225
timestamp 1649977179
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_237
timestamp 1649977179
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_249
timestamp 1649977179
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_261
timestamp 1649977179
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1649977179
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1649977179
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_281
timestamp 1649977179
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_293
timestamp 1649977179
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_305
timestamp 1649977179
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_317
timestamp 1649977179
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_329
timestamp 1649977179
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_335
timestamp 1649977179
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_51_337
timestamp 1649977179
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_349
timestamp 1649977179
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_361
timestamp 1649977179
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_51_373
timestamp 1649977179
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1649977179
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1649977179
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_393
timestamp 1649977179
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_403
timestamp 1649977179
transform 1 0 38180 0 -1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_3
timestamp 1649977179
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_15
timestamp 1649977179
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1649977179
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_29
timestamp 1649977179
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_41
timestamp 1649977179
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_53
timestamp 1649977179
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_65
timestamp 1649977179
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1649977179
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1649977179
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_85
timestamp 1649977179
transform 1 0 8924 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_89
timestamp 1649977179
transform 1 0 9292 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_110
timestamp 1649977179
transform 1 0 11224 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_122
timestamp 1649977179
transform 1 0 12328 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_134
timestamp 1649977179
transform 1 0 13432 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_52_158
timestamp 1649977179
transform 1 0 15640 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_170
timestamp 1649977179
transform 1 0 16744 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_178
timestamp 1649977179
transform 1 0 17480 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_183
timestamp 1649977179
transform 1 0 17940 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_189
timestamp 1649977179
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1649977179
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_197
timestamp 1649977179
transform 1 0 19228 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_205
timestamp 1649977179
transform 1 0 19964 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_212
timestamp 1649977179
transform 1 0 20608 0 1 30464
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_52_218
timestamp 1649977179
transform 1 0 21160 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_230
timestamp 1649977179
transform 1 0 22264 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_242
timestamp 1649977179
transform 1 0 23368 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_250
timestamp 1649977179
transform 1 0 24104 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_52_253
timestamp 1649977179
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_265
timestamp 1649977179
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_277
timestamp 1649977179
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_289
timestamp 1649977179
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1649977179
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1649977179
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_309
timestamp 1649977179
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_321
timestamp 1649977179
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_333
timestamp 1649977179
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_345
timestamp 1649977179
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_357
timestamp 1649977179
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1649977179
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_52_365
timestamp 1649977179
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_52_377
timestamp 1649977179
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_389
timestamp 1649977179
transform 1 0 36892 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_403
timestamp 1649977179
transform 1 0 38180 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_19
timestamp 1649977179
transform 1 0 2852 0 -1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_53_25
timestamp 1649977179
transform 1 0 3404 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_37
timestamp 1649977179
transform 1 0 4508 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_49
timestamp 1649977179
transform 1 0 5612 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1649977179
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_57
timestamp 1649977179
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_69
timestamp 1649977179
transform 1 0 7452 0 -1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_53_92
timestamp 1649977179
transform 1 0 9568 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_104
timestamp 1649977179
transform 1 0 10672 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_53_113
timestamp 1649977179
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_125
timestamp 1649977179
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_137
timestamp 1649977179
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_149
timestamp 1649977179
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_161
timestamp 1649977179
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_167
timestamp 1649977179
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_53_169
timestamp 1649977179
transform 1 0 16652 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_176
timestamp 1649977179
transform 1 0 17296 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_182
timestamp 1649977179
transform 1 0 17848 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_190
timestamp 1649977179
transform 1 0 18584 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_196
timestamp 1649977179
transform 1 0 19136 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_200
timestamp 1649977179
transform 1 0 19504 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_203
timestamp 1649977179
transform 1 0 19780 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_215
timestamp 1649977179
transform 1 0 20884 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_53_223
timestamp 1649977179
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_225
timestamp 1649977179
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_237
timestamp 1649977179
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_249
timestamp 1649977179
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_261
timestamp 1649977179
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_273
timestamp 1649977179
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_279
timestamp 1649977179
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_281
timestamp 1649977179
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_293
timestamp 1649977179
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_305
timestamp 1649977179
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_317
timestamp 1649977179
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_329
timestamp 1649977179
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1649977179
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_337
timestamp 1649977179
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_349
timestamp 1649977179
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_361
timestamp 1649977179
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_53_373
timestamp 1649977179
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_385
timestamp 1649977179
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1649977179
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_53_393
timestamp 1649977179
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_405
timestamp 1649977179
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_54_3
timestamp 1649977179
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_15
timestamp 1649977179
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_27
timestamp 1649977179
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_29
timestamp 1649977179
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_41
timestamp 1649977179
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_53
timestamp 1649977179
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_65
timestamp 1649977179
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_77
timestamp 1649977179
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_83
timestamp 1649977179
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_85
timestamp 1649977179
transform 1 0 8924 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_91
timestamp 1649977179
transform 1 0 9476 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_109
timestamp 1649977179
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_121
timestamp 1649977179
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_133
timestamp 1649977179
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_139
timestamp 1649977179
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_141
timestamp 1649977179
transform 1 0 14076 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_147
timestamp 1649977179
transform 1 0 14628 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_155
timestamp 1649977179
transform 1 0 15364 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_161
timestamp 1649977179
transform 1 0 15916 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_173
timestamp 1649977179
transform 1 0 17020 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_178
timestamp 1649977179
transform 1 0 17480 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_185
timestamp 1649977179
transform 1 0 18124 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_191
timestamp 1649977179
transform 1 0 18676 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1649977179
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_54_197
timestamp 1649977179
transform 1 0 19228 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_201
timestamp 1649977179
transform 1 0 19596 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_211
timestamp 1649977179
transform 1 0 20516 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_54_217
timestamp 1649977179
transform 1 0 21068 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_229
timestamp 1649977179
transform 1 0 22172 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_241
timestamp 1649977179
transform 1 0 23276 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_249
timestamp 1649977179
transform 1 0 24012 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_54_253
timestamp 1649977179
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_265
timestamp 1649977179
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_277
timestamp 1649977179
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_289
timestamp 1649977179
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_301
timestamp 1649977179
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_307
timestamp 1649977179
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_309
timestamp 1649977179
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_321
timestamp 1649977179
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_333
timestamp 1649977179
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_345
timestamp 1649977179
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1649977179
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1649977179
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_54_365
timestamp 1649977179
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_377
timestamp 1649977179
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_54_389
timestamp 1649977179
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_401
timestamp 1649977179
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_55_3
timestamp 1649977179
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_15
timestamp 1649977179
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_27
timestamp 1649977179
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_39
timestamp 1649977179
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1649977179
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1649977179
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_57
timestamp 1649977179
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_69
timestamp 1649977179
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_81
timestamp 1649977179
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_93
timestamp 1649977179
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1649977179
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1649977179
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_113
timestamp 1649977179
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_125
timestamp 1649977179
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_137
timestamp 1649977179
transform 1 0 13708 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_145
timestamp 1649977179
transform 1 0 14444 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_150
timestamp 1649977179
transform 1 0 14904 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_156
timestamp 1649977179
transform 1 0 15456 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_172
timestamp 1649977179
transform 1 0 16928 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_184
timestamp 1649977179
transform 1 0 18032 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_196
timestamp 1649977179
transform 1 0 19136 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_208
timestamp 1649977179
transform 1 0 20240 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_220
timestamp 1649977179
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_55_225
timestamp 1649977179
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_237
timestamp 1649977179
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_249
timestamp 1649977179
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_261
timestamp 1649977179
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_273
timestamp 1649977179
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1649977179
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_281
timestamp 1649977179
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_293
timestamp 1649977179
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_305
timestamp 1649977179
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_317
timestamp 1649977179
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_329
timestamp 1649977179
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_335
timestamp 1649977179
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_337
timestamp 1649977179
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_349
timestamp 1649977179
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_361
timestamp 1649977179
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_55_373
timestamp 1649977179
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_385
timestamp 1649977179
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1649977179
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_55_393
timestamp 1649977179
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_405
timestamp 1649977179
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_56_3
timestamp 1649977179
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_15
timestamp 1649977179
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1649977179
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_29
timestamp 1649977179
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_41
timestamp 1649977179
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_53
timestamp 1649977179
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_65
timestamp 1649977179
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1649977179
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1649977179
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_85
timestamp 1649977179
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_97
timestamp 1649977179
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_109
timestamp 1649977179
transform 1 0 11132 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_56_129
timestamp 1649977179
transform 1 0 12972 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_137
timestamp 1649977179
transform 1 0 13708 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_56_150
timestamp 1649977179
transform 1 0 14904 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_56_158
timestamp 1649977179
transform 1 0 15640 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_56_180
timestamp 1649977179
transform 1 0 17664 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1649977179
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_56_197
timestamp 1649977179
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_209
timestamp 1649977179
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_221
timestamp 1649977179
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_233
timestamp 1649977179
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_245
timestamp 1649977179
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_251
timestamp 1649977179
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_253
timestamp 1649977179
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_265
timestamp 1649977179
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_277
timestamp 1649977179
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_289
timestamp 1649977179
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_301
timestamp 1649977179
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_307
timestamp 1649977179
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_309
timestamp 1649977179
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_321
timestamp 1649977179
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_333
timestamp 1649977179
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_345
timestamp 1649977179
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_357
timestamp 1649977179
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1649977179
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_56_365
timestamp 1649977179
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_377
timestamp 1649977179
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_56_389
timestamp 1649977179
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_401
timestamp 1649977179
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_57_3
timestamp 1649977179
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_15
timestamp 1649977179
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_27
timestamp 1649977179
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_39
timestamp 1649977179
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_51
timestamp 1649977179
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1649977179
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_57
timestamp 1649977179
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_69
timestamp 1649977179
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_81
timestamp 1649977179
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_93
timestamp 1649977179
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1649977179
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1649977179
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_113
timestamp 1649977179
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_125
timestamp 1649977179
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_137
timestamp 1649977179
transform 1 0 13708 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_145
timestamp 1649977179
transform 1 0 14444 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_57_156
timestamp 1649977179
transform 1 0 15456 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_164
timestamp 1649977179
transform 1 0 16192 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_175
timestamp 1649977179
transform 1 0 17204 0 -1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_57_181
timestamp 1649977179
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_193
timestamp 1649977179
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_205
timestamp 1649977179
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1649977179
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1649977179
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_225
timestamp 1649977179
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_237
timestamp 1649977179
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_249
timestamp 1649977179
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_261
timestamp 1649977179
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_273
timestamp 1649977179
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1649977179
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_281
timestamp 1649977179
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_293
timestamp 1649977179
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_305
timestamp 1649977179
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_317
timestamp 1649977179
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_329
timestamp 1649977179
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1649977179
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_337
timestamp 1649977179
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_349
timestamp 1649977179
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_361
timestamp 1649977179
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_57_373
timestamp 1649977179
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_385
timestamp 1649977179
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_391
timestamp 1649977179
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_57_393
timestamp 1649977179
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_405
timestamp 1649977179
transform 1 0 38364 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_58_3
timestamp 1649977179
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_15
timestamp 1649977179
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1649977179
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_29
timestamp 1649977179
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_41
timestamp 1649977179
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_53
timestamp 1649977179
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_65
timestamp 1649977179
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1649977179
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1649977179
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_85
timestamp 1649977179
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_97
timestamp 1649977179
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_109
timestamp 1649977179
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_121
timestamp 1649977179
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1649977179
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1649977179
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_141
timestamp 1649977179
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_153
timestamp 1649977179
transform 1 0 15180 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_157
timestamp 1649977179
transform 1 0 15548 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_175
timestamp 1649977179
transform 1 0 17204 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_187
timestamp 1649977179
transform 1 0 18308 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_195
timestamp 1649977179
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_197
timestamp 1649977179
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_209
timestamp 1649977179
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_221
timestamp 1649977179
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_233
timestamp 1649977179
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_245
timestamp 1649977179
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_251
timestamp 1649977179
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_253
timestamp 1649977179
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_265
timestamp 1649977179
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_277
timestamp 1649977179
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_289
timestamp 1649977179
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_301
timestamp 1649977179
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1649977179
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_309
timestamp 1649977179
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_321
timestamp 1649977179
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_333
timestamp 1649977179
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_345
timestamp 1649977179
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1649977179
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1649977179
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_58_365
timestamp 1649977179
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_377
timestamp 1649977179
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_58_389
timestamp 1649977179
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_401
timestamp 1649977179
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_59_3
timestamp 1649977179
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_15
timestamp 1649977179
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_27
timestamp 1649977179
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_39
timestamp 1649977179
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1649977179
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1649977179
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_57
timestamp 1649977179
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_69
timestamp 1649977179
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_81
timestamp 1649977179
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_93
timestamp 1649977179
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1649977179
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1649977179
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_113
timestamp 1649977179
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_125
timestamp 1649977179
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_137
timestamp 1649977179
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_149
timestamp 1649977179
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_161
timestamp 1649977179
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_167
timestamp 1649977179
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_185
timestamp 1649977179
transform 1 0 18124 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_197
timestamp 1649977179
transform 1 0 19228 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_209
timestamp 1649977179
transform 1 0 20332 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_221
timestamp 1649977179
transform 1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_59_225
timestamp 1649977179
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_237
timestamp 1649977179
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_249
timestamp 1649977179
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_261
timestamp 1649977179
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_273
timestamp 1649977179
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_279
timestamp 1649977179
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_281
timestamp 1649977179
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_293
timestamp 1649977179
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_305
timestamp 1649977179
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_317
timestamp 1649977179
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_329
timestamp 1649977179
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1649977179
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_337
timestamp 1649977179
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_349
timestamp 1649977179
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_361
timestamp 1649977179
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_59_373
timestamp 1649977179
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_385
timestamp 1649977179
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_391
timestamp 1649977179
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_59_393
timestamp 1649977179
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_405
timestamp 1649977179
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_60_3
timestamp 1649977179
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_15
timestamp 1649977179
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1649977179
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_29
timestamp 1649977179
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_41
timestamp 1649977179
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_53
timestamp 1649977179
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_65
timestamp 1649977179
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1649977179
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1649977179
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_85
timestamp 1649977179
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_97
timestamp 1649977179
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_109
timestamp 1649977179
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_121
timestamp 1649977179
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1649977179
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1649977179
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_141
timestamp 1649977179
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_153
timestamp 1649977179
transform 1 0 15180 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_60_176
timestamp 1649977179
transform 1 0 17296 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_188
timestamp 1649977179
transform 1 0 18400 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_60_197
timestamp 1649977179
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_209
timestamp 1649977179
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_221
timestamp 1649977179
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_233
timestamp 1649977179
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_245
timestamp 1649977179
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_251
timestamp 1649977179
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_253
timestamp 1649977179
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_265
timestamp 1649977179
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_277
timestamp 1649977179
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_289
timestamp 1649977179
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_301
timestamp 1649977179
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1649977179
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_309
timestamp 1649977179
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_321
timestamp 1649977179
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_333
timestamp 1649977179
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_345
timestamp 1649977179
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1649977179
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1649977179
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_60_365
timestamp 1649977179
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_377
timestamp 1649977179
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_60_389
timestamp 1649977179
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_401
timestamp 1649977179
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_61_3
timestamp 1649977179
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_15
timestamp 1649977179
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_27
timestamp 1649977179
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_39
timestamp 1649977179
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1649977179
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1649977179
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_74
timestamp 1649977179
transform 1 0 7912 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_82
timestamp 1649977179
transform 1 0 8648 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_100
timestamp 1649977179
transform 1 0 10304 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_113
timestamp 1649977179
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_125
timestamp 1649977179
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_137
timestamp 1649977179
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_149
timestamp 1649977179
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1649977179
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1649977179
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_169
timestamp 1649977179
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_181
timestamp 1649977179
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_193
timestamp 1649977179
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_205
timestamp 1649977179
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_217
timestamp 1649977179
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1649977179
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_225
timestamp 1649977179
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_237
timestamp 1649977179
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_249
timestamp 1649977179
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_261
timestamp 1649977179
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_273
timestamp 1649977179
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1649977179
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_281
timestamp 1649977179
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_293
timestamp 1649977179
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_305
timestamp 1649977179
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_317
timestamp 1649977179
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1649977179
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1649977179
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_337
timestamp 1649977179
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_349
timestamp 1649977179
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_361
timestamp 1649977179
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_61_373
timestamp 1649977179
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1649977179
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1649977179
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_61_393
timestamp 1649977179
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_405
timestamp 1649977179
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_62_3
timestamp 1649977179
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_15
timestamp 1649977179
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1649977179
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_29
timestamp 1649977179
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_41
timestamp 1649977179
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_53
timestamp 1649977179
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_65
timestamp 1649977179
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_77
timestamp 1649977179
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_83
timestamp 1649977179
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_85
timestamp 1649977179
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_97
timestamp 1649977179
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_109
timestamp 1649977179
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_121
timestamp 1649977179
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1649977179
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1649977179
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_141
timestamp 1649977179
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_153
timestamp 1649977179
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_165
timestamp 1649977179
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_177
timestamp 1649977179
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1649977179
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1649977179
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_197
timestamp 1649977179
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_209
timestamp 1649977179
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_221
timestamp 1649977179
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_233
timestamp 1649977179
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_245
timestamp 1649977179
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1649977179
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_253
timestamp 1649977179
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_265
timestamp 1649977179
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_277
timestamp 1649977179
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_289
timestamp 1649977179
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_301
timestamp 1649977179
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_307
timestamp 1649977179
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_309
timestamp 1649977179
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_321
timestamp 1649977179
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_333
timestamp 1649977179
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_345
timestamp 1649977179
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1649977179
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1649977179
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_62_365
timestamp 1649977179
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_377
timestamp 1649977179
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_62_389
timestamp 1649977179
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_401
timestamp 1649977179
transform 1 0 37996 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_3
timestamp 1649977179
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_15
timestamp 1649977179
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_27
timestamp 1649977179
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_39
timestamp 1649977179
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_51
timestamp 1649977179
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_55
timestamp 1649977179
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_57
timestamp 1649977179
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_69
timestamp 1649977179
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_81
timestamp 1649977179
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_93
timestamp 1649977179
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_105
timestamp 1649977179
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1649977179
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_113
timestamp 1649977179
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_125
timestamp 1649977179
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_137
timestamp 1649977179
transform 1 0 13708 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_63_145
timestamp 1649977179
transform 1 0 14444 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_157
timestamp 1649977179
transform 1 0 15548 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_165
timestamp 1649977179
transform 1 0 16284 0 -1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_63_169
timestamp 1649977179
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_181
timestamp 1649977179
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_193
timestamp 1649977179
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_205
timestamp 1649977179
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_217
timestamp 1649977179
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1649977179
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_225
timestamp 1649977179
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_237
timestamp 1649977179
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_249
timestamp 1649977179
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_261
timestamp 1649977179
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_273
timestamp 1649977179
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1649977179
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_281
timestamp 1649977179
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_293
timestamp 1649977179
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_305
timestamp 1649977179
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_317
timestamp 1649977179
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_329
timestamp 1649977179
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_335
timestamp 1649977179
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_337
timestamp 1649977179
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_349
timestamp 1649977179
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_361
timestamp 1649977179
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_63_373
timestamp 1649977179
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1649977179
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1649977179
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_63_393
timestamp 1649977179
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_405
timestamp 1649977179
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_64_3
timestamp 1649977179
transform 1 0 1380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_15
timestamp 1649977179
transform 1 0 2484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1649977179
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_29
timestamp 1649977179
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_41
timestamp 1649977179
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_53
timestamp 1649977179
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_57
timestamp 1649977179
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_69
timestamp 1649977179
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_81
timestamp 1649977179
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_85
timestamp 1649977179
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_97
timestamp 1649977179
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_109
timestamp 1649977179
transform 1 0 11132 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_113
timestamp 1649977179
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_125
timestamp 1649977179
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_137
timestamp 1649977179
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_141
timestamp 1649977179
transform 1 0 14076 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_64_149
timestamp 1649977179
transform 1 0 14812 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_161
timestamp 1649977179
transform 1 0 15916 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_167
timestamp 1649977179
transform 1 0 16468 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_64_169
timestamp 1649977179
transform 1 0 16652 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_181
timestamp 1649977179
transform 1 0 17756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_193
timestamp 1649977179
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_197
timestamp 1649977179
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_209
timestamp 1649977179
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_221
timestamp 1649977179
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_225
timestamp 1649977179
transform 1 0 21804 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_237
timestamp 1649977179
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_249
timestamp 1649977179
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_253
timestamp 1649977179
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_265
timestamp 1649977179
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_277
timestamp 1649977179
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_281
timestamp 1649977179
transform 1 0 26956 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_293
timestamp 1649977179
transform 1 0 28060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_305
timestamp 1649977179
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_309
timestamp 1649977179
transform 1 0 29532 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_317
timestamp 1649977179
transform 1 0 30268 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_321
timestamp 1649977179
transform 1 0 30636 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_328
timestamp 1649977179
transform 1 0 31280 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_64_337
timestamp 1649977179
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_349
timestamp 1649977179
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_361
timestamp 1649977179
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_365
timestamp 1649977179
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_64_377
timestamp 1649977179
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_389
timestamp 1649977179
transform 1 0 36892 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_64_393
timestamp 1649977179
transform 1 0 37260 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_405
timestamp 1649977179
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1649977179
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1649977179
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1649977179
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1649977179
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1649977179
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1649977179
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1649977179
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1649977179
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1649977179
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1649977179
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1649977179
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1649977179
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1649977179
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1649977179
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1649977179
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1649977179
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1649977179
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1649977179
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1649977179
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1649977179
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1649977179
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1649977179
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1649977179
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1649977179
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1649977179
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1649977179
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1649977179
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1649977179
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1649977179
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1649977179
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1649977179
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1649977179
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1649977179
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1649977179
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1649977179
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1649977179
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1649977179
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1649977179
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1649977179
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1649977179
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1649977179
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1649977179
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1649977179
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1649977179
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1649977179
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1649977179
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1649977179
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1649977179
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1649977179
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1649977179
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1649977179
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1649977179
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1649977179
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1649977179
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1649977179
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1649977179
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1649977179
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1649977179
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1649977179
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1649977179
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1649977179
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1649977179
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1649977179
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1649977179
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1649977179
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1649977179
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1649977179
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1649977179
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1649977179
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1649977179
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1649977179
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1649977179
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1649977179
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1649977179
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1649977179
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1649977179
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1649977179
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1649977179
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1649977179
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1649977179
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1649977179
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1649977179
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1649977179
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1649977179
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1649977179
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1649977179
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1649977179
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1649977179
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1649977179
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1649977179
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1649977179
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1649977179
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1649977179
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1649977179
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1649977179
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1649977179
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1649977179
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1649977179
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1649977179
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1649977179
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1649977179
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1649977179
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1649977179
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1649977179
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1649977179
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1649977179
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1649977179
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1649977179
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1649977179
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1649977179
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1649977179
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1649977179
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1649977179
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1649977179
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1649977179
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1649977179
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1649977179
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1649977179
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1649977179
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1649977179
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1649977179
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1649977179
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1649977179
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1649977179
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1649977179
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1649977179
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1649977179
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1649977179
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1649977179
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1649977179
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1649977179
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1649977179
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1649977179
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1649977179
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1649977179
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1649977179
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1649977179
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1649977179
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1649977179
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1649977179
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1649977179
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1649977179
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1649977179
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1649977179
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1649977179
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1649977179
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1649977179
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1649977179
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1649977179
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1649977179
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1649977179
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1649977179
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1649977179
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1649977179
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1649977179
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1649977179
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1649977179
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1649977179
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1649977179
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1649977179
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1649977179
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1649977179
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1649977179
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1649977179
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1649977179
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1649977179
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1649977179
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1649977179
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1649977179
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1649977179
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1649977179
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1649977179
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1649977179
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1649977179
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1649977179
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1649977179
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1649977179
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1649977179
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1649977179
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1649977179
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1649977179
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1649977179
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1649977179
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1649977179
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1649977179
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1649977179
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1649977179
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1649977179
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1649977179
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1649977179
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1649977179
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1649977179
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1649977179
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1649977179
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1649977179
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1649977179
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1649977179
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1649977179
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1649977179
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1649977179
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1649977179
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1649977179
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1649977179
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1649977179
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1649977179
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1649977179
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1649977179
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1649977179
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1649977179
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1649977179
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1649977179
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1649977179
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1649977179
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1649977179
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1649977179
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1649977179
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1649977179
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1649977179
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1649977179
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1649977179
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1649977179
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1649977179
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1649977179
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1649977179
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1649977179
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1649977179
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1649977179
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1649977179
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1649977179
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1649977179
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1649977179
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1649977179
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1649977179
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1649977179
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1649977179
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1649977179
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1649977179
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1649977179
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1649977179
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1649977179
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1649977179
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1649977179
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1649977179
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1649977179
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1649977179
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1649977179
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1649977179
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1649977179
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1649977179
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1649977179
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1649977179
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1649977179
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1649977179
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1649977179
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1649977179
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1649977179
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1649977179
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1649977179
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1649977179
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1649977179
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1649977179
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1649977179
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1649977179
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1649977179
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1649977179
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1649977179
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1649977179
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1649977179
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1649977179
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1649977179
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1649977179
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1649977179
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1649977179
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1649977179
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1649977179
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1649977179
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1649977179
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1649977179
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1649977179
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1649977179
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1649977179
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1649977179
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1649977179
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1649977179
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1649977179
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1649977179
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1649977179
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1649977179
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1649977179
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1649977179
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1649977179
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1649977179
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1649977179
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1649977179
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1649977179
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1649977179
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1649977179
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1649977179
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1649977179
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1649977179
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1649977179
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1649977179
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1649977179
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1649977179
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1649977179
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1649977179
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1649977179
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1649977179
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1649977179
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1649977179
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1649977179
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1649977179
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1649977179
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1649977179
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1649977179
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1649977179
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1649977179
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1649977179
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1649977179
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1649977179
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1649977179
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1649977179
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1649977179
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1649977179
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1649977179
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1649977179
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1649977179
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1649977179
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1649977179
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1649977179
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1649977179
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1649977179
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1649977179
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1649977179
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1649977179
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1649977179
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1649977179
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1649977179
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1649977179
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1649977179
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1649977179
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1649977179
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1649977179
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1649977179
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1649977179
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1649977179
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1649977179
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1649977179
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1649977179
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1649977179
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1649977179
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1649977179
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1649977179
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1649977179
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1649977179
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1649977179
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1649977179
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1649977179
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1649977179
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1649977179
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1649977179
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1649977179
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1649977179
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1649977179
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1649977179
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1649977179
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1649977179
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1649977179
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1649977179
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1649977179
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1649977179
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1649977179
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1649977179
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1649977179
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1649977179
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1649977179
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1649977179
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1649977179
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1649977179
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1649977179
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1649977179
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1649977179
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1649977179
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1649977179
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1649977179
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1649977179
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1649977179
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1649977179
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1649977179
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1649977179
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1649977179
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1649977179
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1649977179
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1649977179
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1649977179
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1649977179
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1649977179
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1649977179
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1649977179
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1649977179
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1649977179
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1649977179
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1649977179
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1649977179
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1649977179
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1649977179
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1649977179
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1649977179
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1649977179
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1649977179
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1649977179
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1649977179
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1649977179
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1649977179
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1649977179
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1649977179
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1649977179
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1649977179
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1649977179
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1649977179
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1649977179
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1649977179
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1649977179
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1649977179
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1649977179
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1649977179
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1649977179
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1649977179
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1649977179
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1649977179
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1649977179
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1649977179
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1649977179
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1649977179
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1649977179
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1649977179
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1649977179
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1649977179
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1649977179
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1649977179
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1649977179
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1649977179
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1649977179
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1649977179
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1649977179
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1649977179
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1649977179
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1649977179
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1649977179
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1649977179
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1649977179
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1649977179
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1649977179
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1649977179
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1649977179
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1649977179
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1649977179
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1649977179
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1649977179
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1649977179
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1649977179
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1649977179
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1649977179
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1649977179
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1649977179
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1649977179
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1649977179
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1649977179
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1649977179
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1649977179
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1649977179
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1649977179
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1649977179
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1649977179
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1649977179
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1649977179
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1649977179
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1649977179
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1649977179
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1649977179
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1649977179
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1649977179
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1649977179
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1649977179
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1649977179
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1649977179
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1649977179
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1649977179
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1649977179
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1649977179
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1649977179
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1649977179
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1649977179
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1649977179
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1649977179
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1649977179
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1649977179
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1649977179
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1649977179
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1649977179
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1649977179
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1649977179
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1649977179
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1649977179
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1649977179
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1649977179
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1649977179
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1649977179
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1649977179
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1649977179
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1649977179
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1649977179
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1649977179
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1649977179
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1649977179
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1649977179
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1649977179
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1649977179
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1649977179
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1649977179
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1649977179
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1649977179
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1649977179
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1649977179
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1649977179
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1649977179
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1649977179
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1649977179
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1649977179
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1649977179
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1649977179
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1649977179
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1649977179
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1649977179
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1649977179
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1649977179
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1649977179
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1649977179
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1649977179
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1649977179
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1649977179
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1649977179
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1649977179
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1649977179
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1649977179
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1649977179
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1649977179
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1649977179
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1649977179
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1649977179
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1649977179
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1649977179
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1649977179
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1649977179
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1649977179
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1649977179
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1649977179
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1649977179
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1649977179
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1649977179
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1649977179
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1649977179
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1649977179
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1649977179
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1649977179
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1649977179
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1649977179
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1649977179
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1649977179
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1649977179
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1649977179
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1649977179
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1649977179
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1649977179
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1649977179
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1649977179
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1649977179
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1649977179
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1649977179
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1649977179
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1649977179
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1649977179
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1649977179
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1649977179
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1649977179
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1649977179
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1649977179
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1649977179
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1649977179
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1649977179
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1649977179
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1649977179
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1649977179
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1649977179
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1649977179
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1649977179
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1649977179
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1649977179
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_2  _114_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18676 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__buf_1  _115_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 37812 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _116_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13064 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _117_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 22632 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _118_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20332 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _119_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 19780 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _120_
timestamp 1649977179
transform 1 0 21528 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _121_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20516 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_2  _122_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21804 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_4  _123_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21344 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _124_
timestamp 1649977179
transform 1 0 23276 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _125_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 22448 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _126_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20608 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _127_
timestamp 1649977179
transform 1 0 20792 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _128_
timestamp 1649977179
transform -1 0 22172 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__o22ai_2  _129_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 21344 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _130_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21344 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_4  _131_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20976 0 1 21760
box -38 -48 1326 592
use sky130_fd_sc_hd__o21bai_1  _132_
timestamp 1649977179
transform -1 0 24656 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _133_
timestamp 1649977179
transform 1 0 22080 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _134_
timestamp 1649977179
transform 1 0 22724 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _135_
timestamp 1649977179
transform -1 0 23828 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _136_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 23092 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _137_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19228 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _138_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19780 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_1  _139_
timestamp 1649977179
transform 1 0 21804 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _140_
timestamp 1649977179
transform 1 0 18860 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2ai_1  _141_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 19688 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _142_
timestamp 1649977179
transform -1 0 22356 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _143_
timestamp 1649977179
transform 1 0 21436 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_4  _144_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 23368 0 -1 21760
box -38 -48 1602 592
use sky130_fd_sc_hd__a21oi_1  _145_
timestamp 1649977179
transform 1 0 14996 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_1  _146_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20516 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _147_
timestamp 1649977179
transform 1 0 16652 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _148_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 22264 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _149_
timestamp 1649977179
transform -1 0 22908 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _150_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20700 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__o2bb2ai_1  _151_
timestamp 1649977179
transform 1 0 17480 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _152_
timestamp 1649977179
transform -1 0 17020 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _153_
timestamp 1649977179
transform 1 0 11868 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _154_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12972 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _155_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 11960 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _156_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 9936 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _157_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17296 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and4_2  _158_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14444 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _159_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 15732 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _160_
timestamp 1649977179
transform 1 0 9200 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _161_
timestamp 1649977179
transform 1 0 8924 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _162_
timestamp 1649977179
transform 1 0 12972 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _163_
timestamp 1649977179
transform -1 0 12788 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _164_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 13616 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _165_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14076 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _166_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 13708 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _167_
timestamp 1649977179
transform -1 0 15088 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _168_
timestamp 1649977179
transform -1 0 13984 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _169_
timestamp 1649977179
transform -1 0 7912 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _170_
timestamp 1649977179
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _171_
timestamp 1649977179
transform 1 0 19320 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _172_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 20148 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_2  _173_
timestamp 1649977179
transform 1 0 18492 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__a22oi_1  _174_
timestamp 1649977179
transform 1 0 20056 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _175_
timestamp 1649977179
transform 1 0 16744 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a41o_1  _176_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18492 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _177_
timestamp 1649977179
transform -1 0 14260 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a31oi_1  _178_
timestamp 1649977179
transform -1 0 14720 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _179_
timestamp 1649977179
transform 1 0 19596 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _180_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 18032 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _181_
timestamp 1649977179
transform -1 0 18768 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _182_
timestamp 1649977179
transform -1 0 15548 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _183_
timestamp 1649977179
transform 1 0 19320 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _184_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 21068 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _185_
timestamp 1649977179
transform 1 0 17572 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _186_
timestamp 1649977179
transform -1 0 18676 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _187_
timestamp 1649977179
transform 1 0 12328 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _188_
timestamp 1649977179
transform -1 0 17388 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _189_
timestamp 1649977179
transform -1 0 10764 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _190_
timestamp 1649977179
transform 1 0 11408 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand4_1  _191_
timestamp 1649977179
transform 1 0 17020 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _192_
timestamp 1649977179
transform 1 0 17848 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _193_
timestamp 1649977179
transform -1 0 18216 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _194_
timestamp 1649977179
transform -1 0 15180 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _195_
timestamp 1649977179
transform 1 0 15732 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand4_1  _196_
timestamp 1649977179
transform -1 0 15916 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _197_
timestamp 1649977179
transform 1 0 14904 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _198_
timestamp 1649977179
transform -1 0 15824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _199_
timestamp 1649977179
transform -1 0 14260 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _200_
timestamp 1649977179
transform -1 0 19964 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_1  _201_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 23184 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _202_
timestamp 1649977179
transform -1 0 24472 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _203_
timestamp 1649977179
transform -1 0 11868 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_4  _204_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 15456 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  _205_
timestamp 1649977179
transform 1 0 18860 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a41oi_1  _206_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 20148 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _207_
timestamp 1649977179
transform 1 0 19688 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _208_
timestamp 1649977179
transform -1 0 18124 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a41oi_1  _209_
timestamp 1649977179
transform 1 0 17940 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _210_
timestamp 1649977179
transform -1 0 17480 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__a41oi_1  _211_
timestamp 1649977179
transform 1 0 19228 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _212_
timestamp 1649977179
transform -1 0 19412 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _213_
timestamp 1649977179
transform 1 0 11500 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _214_
timestamp 1649977179
transform 1 0 9752 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_1  _215_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9660 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__and2_2  _216_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 14812 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _217_
timestamp 1649977179
transform 1 0 10396 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _218_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 11868 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _219_
timestamp 1649977179
transform -1 0 12880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _220_
timestamp 1649977179
transform -1 0 15456 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _221_
timestamp 1649977179
transform -1 0 16928 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _222_
timestamp 1649977179
transform -1 0 14904 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _223_
timestamp 1649977179
transform -1 0 14904 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _224_
timestamp 1649977179
transform 1 0 8924 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _225_
timestamp 1649977179
transform 1 0 7452 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _226_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 18584 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _227_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 17204 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _228_
timestamp 1649977179
transform 1 0 16836 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__dfxtp_2  _229_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 12972 0 1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _230_
timestamp 1649977179
transform -1 0 17204 0 1 33728
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _231_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 12236 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _232_
timestamp 1649977179
transform 1 0 7452 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _233_
timestamp 1649977179
transform 1 0 8004 0 -1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _234_
timestamp 1649977179
transform 1 0 16652 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _235_
timestamp 1649977179
transform 1 0 8280 0 -1 26112
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _236_
timestamp 1649977179
transform 1 0 6348 0 -1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _237_
timestamp 1649977179
transform -1 0 17296 0 1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _238_
timestamp 1649977179
transform 1 0 16652 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _239_
timestamp 1649977179
transform 1 0 15916 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _240_
timestamp 1649977179
transform 1 0 7636 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _241_
timestamp 1649977179
transform 1 0 14076 0 1 30464
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _242_
timestamp 1649977179
transform 1 0 16652 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _243_
timestamp 1649977179
transform 1 0 16192 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _244_
timestamp 1649977179
transform 1 0 11592 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _245_
timestamp 1649977179
transform 1 0 1380 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _246_
timestamp 1649977179
transform 1 0 2484 0 -1 28288
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _247_
timestamp 1649977179
transform 1 0 8740 0 -1 35904
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_4  _248_ opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 3772 0 1 26112
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_2  _249_
timestamp 1649977179
transform 1 0 9568 0 1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_2  _250_
timestamp 1649977179
transform 1 0 1380 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _251_
timestamp 1649977179
transform 1 0 12972 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _252_
timestamp 1649977179
transform -1 0 17296 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _253_
timestamp 1649977179
transform 1 0 14720 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _254_
timestamp 1649977179
transform 1 0 1380 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _255_
timestamp 1649977179
transform 1 0 16652 0 -1 25024
box -38 -48 1602 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_i_clk opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 9384 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_res_clk
timestamp 1649977179
transform 1 0 17756 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_i_clk
timestamp 1649977179
transform -1 0 7084 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f_res_clk
timestamp 1649977179
transform -1 0 17480 0 1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_i_clk
timestamp 1649977179
transform 1 0 10396 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f_res_clk
timestamp 1649977179
transform 1 0 18216 0 -1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input2 opt/silicon/pdk/sky130B/libs.ref/sky130_fd_sc_hd/mag
timestamp 1649977179
transform -1 0 35420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1649977179
transform 1 0 31004 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1649977179
transform -1 0 38180 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1649977179
transform -1 0 1656 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1649977179
transform 1 0 16836 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1649977179
transform 1 0 14444 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  output8
timestamp 1649977179
transform -1 0 38180 0 1 11968
box -38 -48 314 592
<< labels >>
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 clock_sel
port 0 nsew signal input
flabel metal2 s 34150 0 34206 800 0 FreeSans 224 90 0 0 div[0]
port 1 nsew signal input
flabel metal2 s 30930 39200 30986 40000 0 FreeSans 224 90 0 0 div[1]
port 2 nsew signal input
flabel metal3 s 39200 30608 40000 30728 0 FreeSans 480 0 0 0 div[2]
port 3 nsew signal input
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 div[3]
port 4 nsew signal input
flabel metal2 s 16762 0 16818 800 0 FreeSans 224 90 0 0 div_we
port 5 nsew signal input
flabel metal3 s 0 36048 800 36168 0 FreeSans 480 0 0 0 i_clk
port 6 nsew signal input
flabel metal2 s 13542 39200 13598 40000 0 FreeSans 224 90 0 0 i_rst
port 7 nsew signal input
flabel metal3 s 39200 12248 40000 12368 0 FreeSans 480 0 0 0 o_clk
port 8 nsew signal tristate
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 1920 90 0 0 vccd1
port 9 nsew power bidirectional
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 1920 90 0 0 vccd1
port 9 nsew power bidirectional
flabel metal4 s 19568 2128 19888 37584 0 FreeSans 1920 90 0 0 vssd1
port 10 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
