* NGSPICE file created from alu.ext - technology: sky130B

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_2 abstract view
.subckt sky130_fd_sc_hd__o32a_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

.subckt alu i_carry i_l[0] i_l[10] i_l[11] i_l[12] i_l[13] i_l[14] i_l[15] i_l[1]
+ i_l[2] i_l[3] i_l[4] i_l[5] i_l[6] i_l[7] i_l[8] i_l[9] i_mode[0] i_mode[1] i_mode[2]
+ i_mode[3] i_r[0] i_r[10] i_r[11] i_r[12] i_r[13] i_r[14] i_r[15] i_r[1] i_r[2] i_r[3]
+ i_r[4] i_r[5] i_r[6] i_r[7] i_r[8] i_r[9] o_flags[0] o_flags[1] o_flags[2] o_flags[3]
+ o_flags[4] o_out[0] o_out[10] o_out[11] o_out[12] o_out[13] o_out[14] o_out[15]
+ o_out[1] o_out[2] o_out[3] o_out[4] o_out[5] o_out[6] o_out[7] o_out[8] o_out[9]
+ vccd1 vssd1
XFILLER_39_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0703__A _0738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0708__B1 _0729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0985_ _0808_/X _0948_/C _0985_/S vssd1 vssd1 vccd1 vccd1 _0985_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0947__B1 _0808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0770_ _0770_/A _0858_/S _0770_/C _0669_/A vssd1 vssd1 vccd1 vccd1 _0770_/X sky130_fd_sc_hd__or4b_1
XANTENNA__1174__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0632__A2 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0968_ _0975_/A _0965_/Y _1014_/A vssd1 vssd1 vccd1 vccd1 _1043_/A sky130_fd_sc_hd__a21o_1
X_0899_ _0954_/A _0952_/A vssd1 vssd1 vccd1 vccd1 _0901_/A sky130_fd_sc_hd__or2_1
XFILLER_23_75 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0822_ _0800_/A _0798_/B _0805_/A vssd1 vssd1 vccd1 vccd1 _0823_/B sky130_fd_sc_hd__a21oi_1
XANTENNA__1169__A _1169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0753_ _0759_/A _0796_/B vssd1 vssd1 vccd1 vccd1 _0754_/B sky130_fd_sc_hd__or2_1
X_0684_ _0684_/A _0684_/B vssd1 vssd1 vccd1 vccd1 _0684_/Y sky130_fd_sc_hd__nand2_1
X_1167_ _1167_/A _1167_/B _1167_/C _1167_/D vssd1 vssd1 vccd1 vccd1 _1168_/C sky130_fd_sc_hd__or4_1
XFILLER_44_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1098_ _0861_/X _0923_/Y _1096_/X _1097_/X vssd1 vssd1 vccd1 vccd1 _1098_/X sky130_fd_sc_hd__o211a_1
XANTENNA__1079__A _1108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_172 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1021_ _1019_/X _1021_/B vssd1 vssd1 vccd1 vccd1 _1021_/X sky130_fd_sc_hd__and2b_1
X_0805_ _0805_/A _0805_/B vssd1 vssd1 vccd1 vccd1 _0805_/Y sky130_fd_sc_hd__nor2_1
X_0736_ _0738_/S _0736_/B vssd1 vssd1 vccd1 vccd1 _0736_/Y sky130_fd_sc_hd__nor2_1
X_0667_ _1155_/A input7/X vssd1 vssd1 vccd1 vccd1 _0669_/B sky130_fd_sc_hd__or2_1
X_0598_ _0843_/A _0598_/B vssd1 vssd1 vccd1 vccd1 _1126_/A sky130_fd_sc_hd__nor2_1
XFILLER_37_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0677__S _0738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0762__A1 _0796_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input18_A i_mode[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1166__B _1166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1004_ _1004_/A vssd1 vssd1 vccd1 vccd1 _1004_/Y sky130_fd_sc_hd__inv_2
X_0719_ _0719_/A _0719_/B vssd1 vssd1 vccd1 vccd1 _1167_/B sky130_fd_sc_hd__nand2_2
XFILLER_25_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0680__A0 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput53 _1168_/A vssd1 vssd1 vccd1 vccd1 o_out[4] sky130_fd_sc_hd__buf_2
Xoutput42 _1150_/Y vssd1 vssd1 vccd1 vccd1 o_flags[4] sky130_fd_sc_hd__buf_2
XANTENNA__0602__C _0975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0983__A1 _1003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1160__A1 _1131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0726__A1 _0738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0708__A1 _0733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0984_ _1097_/B _0984_/B vssd1 vssd1 vccd1 vccd1 _0984_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__0947__A1 _0975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0865__B1 _0729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0967_ _0966_/Y _0975_/B _0992_/A vssd1 vssd1 vccd1 vccd1 _1014_/A sky130_fd_sc_hd__o21a_1
X_0898_ _0748_/X _0877_/X _0891_/X _0897_/X vssd1 vssd1 vccd1 vccd1 _1165_/B sky130_fd_sc_hd__o211ai_2
XANTENNA__0709__A _0733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0619__A _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0752_ _0759_/A _0796_/B vssd1 vssd1 vccd1 vccd1 _0754_/A sky130_fd_sc_hd__nand2_1
X_0821_ _0821_/A _0821_/B vssd1 vssd1 vccd1 vccd1 _0913_/B sky130_fd_sc_hd__nand2_1
XFILLER_9_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1169__B _1169_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0683_ _0848_/B _0892_/A _0925_/A _0952_/A _0858_/S _0733_/A vssd1 vssd1 vccd1 vccd1
+ _0684_/B sky130_fd_sc_hd__mux4_1
X_1166_ _1166_/A _1166_/B vssd1 vssd1 vccd1 vccd1 _1171_/B sky130_fd_sc_hd__or2_1
X_1097_ _1097_/A _1097_/B _1097_/C vssd1 vssd1 vccd1 vccd1 _1097_/X sky130_fd_sc_hd__or3_1
XFILLER_50_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0902__A _0905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1020_ _1014_/Y _0974_/B _0974_/C _1043_/C vssd1 vssd1 vccd1 vccd1 _1021_/B sky130_fd_sc_hd__a31o_1
XFILLER_15_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_184 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0804_ _0805_/A _0805_/B vssd1 vssd1 vccd1 vccd1 _0831_/B sky130_fd_sc_hd__and2_1
X_0735_ _1097_/C _0734_/X _1007_/A vssd1 vssd1 vccd1 vccd1 _0984_/B sky130_fd_sc_hd__mux2_1
X_0666_ _0759_/A vssd1 vssd1 vccd1 vccd1 _1006_/A sky130_fd_sc_hd__buf_2
X_0597_ _1131_/A _0597_/B vssd1 vssd1 vccd1 vccd1 _0598_/B sky130_fd_sc_hd__xnor2_1
X_1149_ _1149_/A _1149_/B vssd1 vssd1 vccd1 vccd1 _1150_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__0706__B input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0762__A2 _0657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1003_ _1003_/A _1003_/B vssd1 vssd1 vccd1 vccd1 _1003_/Y sky130_fd_sc_hd__nand2_1
XFILLER_19_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0718_ _0692_/X _1103_/A _1003_/A _0717_/Y vssd1 vssd1 vccd1 vccd1 _0719_/B sky130_fd_sc_hd__o31a_1
X_0649_ _0747_/A _0653_/B _0653_/A _0720_/A vssd1 vssd1 vccd1 vccd1 _0808_/A sky130_fd_sc_hd__and4bb_2
XANTENNA__0680__A1 _0763_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0983__A2 _0744_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput54 _1168_/B vssd1 vssd1 vccd1 vccd1 o_out[5] sky130_fd_sc_hd__buf_2
Xoutput43 _1167_/A vssd1 vssd1 vccd1 vccd1 o_out[0] sky130_fd_sc_hd__buf_2
XFILLER_0_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input30_A i_r[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1127__C1 _0866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0708__A2 _0834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0947__A2 _0834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0983_ _1003_/A _0744_/X _1125_/A vssd1 vssd1 vccd1 vccd1 _0983_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_37_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0905__A _0905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0865__A1 _0894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0815__A _0815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0897_ _0910_/A _0853_/Y _0912_/B _0896_/Y _0824_/A vssd1 vssd1 vccd1 vccd1 _0897_/X
+ sky130_fd_sc_hd__a311o_1
X_0966_ _0975_/A vssd1 vssd1 vccd1 vccd1 _0966_/Y sky130_fd_sc_hd__inv_2
XANTENNA__0709__B input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0725__A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0847__A1 _0848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0751_ _0751_/A vssd1 vssd1 vccd1 vccd1 _1119_/A sky130_fd_sc_hd__clkbuf_4
X_0820_ _0820_/A _1131_/A _0820_/C vssd1 vssd1 vccd1 vccd1 _0821_/B sky130_fd_sc_hd__nand3_1
XFILLER_14_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0682_ _0874_/B vssd1 vssd1 vccd1 vccd1 _0925_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_49_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1096_ _1081_/A _1094_/Y _1095_/X vssd1 vssd1 vccd1 vccd1 _1096_/X sky130_fd_sc_hd__o21ba_1
X_1165_ _1165_/A _1165_/B vssd1 vssd1 vccd1 vccd1 _1171_/A sky130_fd_sc_hd__or2_1
XFILLER_20_222 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0774__A0 _0874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0949_ _0975_/B _0656_/B _1132_/A _0948_/X vssd1 vssd1 vccd1 vccd1 _0949_/X sky130_fd_sc_hd__a211o_1
XFILLER_47_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0902__B _0925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0803_ _0757_/A _0754_/B _0757_/B _0759_/X vssd1 vssd1 vccd1 vccd1 _0805_/B sky130_fd_sc_hd__a31o_1
X_0734_ _0608_/Y _0613_/Y _0781_/A vssd1 vssd1 vccd1 vccd1 _0734_/X sky130_fd_sc_hd__mux2_1
X_0665_ _0665_/A _0665_/B vssd1 vssd1 vccd1 vccd1 _1167_/A sky130_fd_sc_hd__nand2_2
X_0596_ _1130_/A _1131_/B vssd1 vssd1 vccd1 vccd1 _0597_/B sky130_fd_sc_hd__or2_1
XFILLER_37_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1079_ _1108_/A input7/X vssd1 vssd1 vccd1 vccd1 _1081_/A sky130_fd_sc_hd__nor2_1
X_1148_ _1148_/A _1148_/B vssd1 vssd1 vccd1 vccd1 _1149_/B sky130_fd_sc_hd__xnor2_1
XFILLER_4_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1163__B1 _0748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1002_ _1102_/S _1002_/B vssd1 vssd1 vccd1 vccd1 _1002_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_199 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0717_ _0703_/Y _0705_/X _0716_/X vssd1 vssd1 vccd1 vccd1 _0717_/Y sky130_fd_sc_hd__a21oi_1
X_0648_ _0653_/B _0653_/C _0653_/A vssd1 vssd1 vccd1 vccd1 _0729_/A sky130_fd_sc_hd__and3b_2
X_0579_ _0759_/A _0771_/S _0770_/A _0693_/B vssd1 vssd1 vccd1 vccd1 _1131_/B sky130_fd_sc_hd__or4_2
XFILLER_40_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0680__A2 _0796_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0733__A _0733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0879__S _1099_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput44 _1166_/A vssd1 vssd1 vccd1 vccd1 o_out[10] sky130_fd_sc_hd__buf_2
XFILLER_48_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput55 _1165_/A vssd1 vssd1 vccd1 vccd1 o_out[6] sky130_fd_sc_hd__buf_2
XANTENNA_input23_A i_r[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1127__B1 _0808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0728__A _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0810__C1 _0866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_272 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0982_ _1124_/A _0982_/B vssd1 vssd1 vccd1 vccd1 _0982_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__0820__B _1131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1060__A2 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0865__A2 _0834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0896_ _0910_/A _0853_/Y _0912_/B vssd1 vssd1 vccd1 vccd1 _0896_/Y sky130_fd_sc_hd__a21oi_1
X_0965_ _0975_/B _0992_/A vssd1 vssd1 vccd1 vccd1 _0965_/Y sky130_fd_sc_hd__nor2_1
XFILLER_23_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0847__A2 _0848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0916__A _1173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0750_ _0750_/A _0750_/B vssd1 vssd1 vccd1 vccd1 _1167_/C sky130_fd_sc_hd__nand2_2
X_0681_ _0684_/A _0681_/B vssd1 vssd1 vccd1 vccd1 _0681_/Y sky130_fd_sc_hd__nand2_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1095_ input7/X _0656_/B _1118_/A _0948_/C _1132_/A vssd1 vssd1 vccd1 vccd1 _1095_/X
+ sky130_fd_sc_hd__a221o_1
X_1164_ _1173_/A _1154_/X _1162_/X _1163_/Y vssd1 vssd1 vccd1 vccd1 _1164_/X sky130_fd_sc_hd__a211o_1
X_0948_ _0975_/A _0975_/B _0948_/C vssd1 vssd1 vccd1 vccd1 _0948_/X sky130_fd_sc_hd__and3_1
XFILLER_20_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0774__A1 _0952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0879_ _0925_/A _0892_/A _1099_/S vssd1 vssd1 vccd1 vccd1 _0879_/X sky130_fd_sc_hd__mux2_1
XFILLER_28_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0736__A _0738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0765__A1 _0781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0802_ _1173_/A _0802_/B vssd1 vssd1 vccd1 vccd1 _0802_/Y sky130_fd_sc_hd__nand2_1
X_0733_ _0733_/A _0733_/B vssd1 vssd1 vccd1 vccd1 _1097_/C sky130_fd_sc_hd__or2_1
X_0664_ _0886_/A _0621_/X _1006_/B _0663_/X vssd1 vssd1 vccd1 vccd1 _0665_/B sky130_fd_sc_hd__o31a_1
XFILLER_6_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0595_ _0653_/A _0653_/B _0595_/C _0595_/D vssd1 vssd1 vccd1 vccd1 _1130_/A sky130_fd_sc_hd__nand4b_2
XFILLER_37_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_81 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1078_ _1078_/A vssd1 vssd1 vccd1 vccd1 _1170_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_1147_ _1166_/A _1166_/B vssd1 vssd1 vccd1 vccd1 _1148_/B sky130_fd_sc_hd__xor2_1
XFILLER_20_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_20_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0683__A0 _0848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0986__A1 _0866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1001_ _0941_/Y _1000_/Y _1101_/S vssd1 vssd1 vccd1 vccd1 _1002_/B sky130_fd_sc_hd__mux2_1
XFILLER_19_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0716_ _0711_/B _0708_/X _0714_/X _0715_/X vssd1 vssd1 vccd1 vccd1 _0716_/X sky130_fd_sc_hd__a211o_1
X_0647_ _0720_/A _0747_/A vssd1 vssd1 vccd1 vccd1 _0653_/C sky130_fd_sc_hd__nor2_1
X_0578_ _0631_/B vssd1 vssd1 vccd1 vccd1 _0693_/B sky130_fd_sc_hd__clkbuf_4
XANTENNA__1154__B2 _1110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0680__A3 _0815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_156 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0968__A1 _0975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_266 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput56 _1165_/B vssd1 vssd1 vccd1 vccd1 o_out[7] sky130_fd_sc_hd__buf_2
Xoutput45 _1166_/B vssd1 vssd1 vccd1 vccd1 o_out[11] sky130_fd_sc_hd__buf_2
XANTENNA_input16_A i_l[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0834__A _0834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input8_A i_l[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1127__A1 _1110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_45 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0810__B1 _0729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_181 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0629__A0 _0763_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0981_ _0860_/X _0980_/X _1102_/S vssd1 vssd1 vccd1 vccd1 _0982_/B sky130_fd_sc_hd__mux2_1
XFILLER_8_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0964_ _0964_/A _0985_/S vssd1 vssd1 vccd1 vccd1 _0992_/A sky130_fd_sc_hd__nor2_2
X_0895_ _0895_/A _0895_/B vssd1 vssd1 vccd1 vccd1 _0912_/B sky130_fd_sc_hd__nand2_1
XFILLER_4_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1009__B1 _0808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0680_ input9/X _0763_/B _0796_/B _0815_/A _0858_/S _0733_/A vssd1 vssd1 vccd1 vccd1
+ _0681_/B sky130_fd_sc_hd__mux4_1
XFILLER_49_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1003__A _1003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1094_ _1108_/A _0834_/X _0808_/X _1093_/Y _0866_/X vssd1 vssd1 vccd1 vccd1 _1094_/Y
+ sky130_fd_sc_hd__a221oi_1
X_1163_ _1111_/A _1119_/B _0748_/X vssd1 vssd1 vccd1 vccd1 _1163_/Y sky130_fd_sc_hd__a21oi_1
X_0947_ _0975_/A _0834_/X _0808_/X _0935_/A _0866_/X vssd1 vssd1 vccd1 vccd1 _0947_/X
+ sky130_fd_sc_hd__a221o_1
X_0878_ _0878_/A vssd1 vssd1 vccd1 vccd1 _0878_/X sky130_fd_sc_hd__buf_2
XFILLER_18_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0752__A _0759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_246 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0646__B _0693_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0801_ _0800_/A _0913_/A _0800_/Y vssd1 vssd1 vccd1 vccd1 _0802_/B sky130_fd_sc_hd__a21o_1
X_0732_ _0757_/A _0730_/X _0731_/X vssd1 vssd1 vccd1 vccd1 _0732_/Y sky130_fd_sc_hd__a21oi_1
X_0594_ _0653_/B _0653_/A _0747_/A _0720_/A vssd1 vssd1 vccd1 vccd1 _1161_/A sky130_fd_sc_hd__and4b_1
X_0663_ _1097_/B _0640_/X _0652_/Y _0662_/X vssd1 vssd1 vccd1 vccd1 _0663_/X sky130_fd_sc_hd__o211a_1
XFILLER_37_154 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1146_ _1146_/A _1146_/B vssd1 vssd1 vccd1 vccd1 _1148_/A sky130_fd_sc_hd__xnor2_1
XFILLER_1_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1077_ _1077_/A _1077_/B _1077_/C _1077_/D vssd1 vssd1 vccd1 vccd1 _1078_/A sky130_fd_sc_hd__or4_1
XFILLER_20_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0683__A1 _0892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1000_ _0878_/X _0999_/X _1073_/A vssd1 vssd1 vccd1 vccd1 _1000_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_42_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0674__A1 _0779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0715_ _0808_/A _0711_/B _0711_/C _0657_/X input9/X vssd1 vssd1 vccd1 vccd1 _0715_/X
+ sky130_fd_sc_hd__a32o_1
X_0646_ input2/X _0693_/B vssd1 vssd1 vccd1 vccd1 _0646_/X sky130_fd_sc_hd__and2_1
XFILLER_25_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1129_ _1110_/A input8/X _0948_/C _0656_/B vssd1 vssd1 vccd1 vccd1 _1132_/B sky130_fd_sc_hd__a31o_1
Xoutput57 _1169_/A vssd1 vssd1 vccd1 vccd1 o_out[8] sky130_fd_sc_hd__buf_2
XFILLER_31_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput46 _1170_/A vssd1 vssd1 vccd1 vccd1 o_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_47_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0629_ _0763_/B _0796_/B _0779_/S vssd1 vssd1 vccd1 vccd1 _0629_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1127__A2 _0834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0810__A1 _1131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0629__A1 _0796_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_260 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0980_ _0918_/Y _0979_/Y _1101_/S vssd1 vssd1 vccd1 vccd1 _0980_/X sky130_fd_sc_hd__mux2_1
XFILLER_12_160 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0670__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0845__A _0894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0786__A0 _0815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0894_ _0894_/A _0894_/B _0894_/C vssd1 vssd1 vccd1 vccd1 _0895_/B sky130_fd_sc_hd__nand3_1
X_0963_ _1015_/A input3/X vssd1 vssd1 vccd1 vccd1 _0985_/S sky130_fd_sc_hd__and2_2
XANTENNA__0710__B1 input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1009__A1 _1039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0940__A0 _0975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1162_ _0598_/B _1158_/Y _1161_/X vssd1 vssd1 vccd1 vccd1 _1162_/X sky130_fd_sc_hd__o21a_1
X_1093_ _1118_/A vssd1 vssd1 vccd1 vccd1 _1093_/Y sky130_fd_sc_hd__inv_2
X_0877_ _0894_/C _0877_/B vssd1 vssd1 vccd1 vccd1 _0877_/X sky130_fd_sc_hd__xor2_1
XFILLER_20_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0946_ _1124_/A _0939_/Y _0943_/Y _0944_/Y _0945_/Y vssd1 vssd1 vccd1 vccd1 _0946_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_18_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0752__B _0796_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0998__B1 _1119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0731_ _0763_/B _0657_/X _0746_/A _0808_/A vssd1 vssd1 vccd1 vccd1 _0731_/X sky130_fd_sc_hd__a22o_1
X_0800_ _0800_/A _0805_/A vssd1 vssd1 vccd1 vccd1 _0800_/Y sky130_fd_sc_hd__nor2_1
XFILLER_6_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0662_ input2/X _0657_/X _0660_/X _0661_/Y vssd1 vssd1 vccd1 vccd1 _0662_/X sky130_fd_sc_hd__o2bb2a_1
X_0593_ _0595_/C vssd1 vssd1 vccd1 vccd1 _0720_/A sky130_fd_sc_hd__buf_2
XFILLER_34_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1145_ _1169_/A _1145_/B vssd1 vssd1 vccd1 vccd1 _1146_/B sky130_fd_sc_hd__xnor2_1
X_1076_ _1103_/A _1076_/B vssd1 vssd1 vccd1 vccd1 _1077_/D sky130_fd_sc_hd__nor2_1
X_0929_ _0886_/B _0600_/B _0923_/Y _0928_/Y vssd1 vssd1 vccd1 vccd1 _0929_/X sky130_fd_sc_hd__o31a_1
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0683__A2 _0925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0674__A2 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0673__A _1155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0714_ _0745_/B _0751_/A _0714_/C vssd1 vssd1 vccd1 vccd1 _0714_/X sky130_fd_sc_hd__and3b_1
X_0645_ _0720_/A _0747_/A _0720_/C vssd1 vssd1 vccd1 vccd1 _0834_/A sky130_fd_sc_hd__and3b_2
XANTENNA__0612__S _0693_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0848__A _0848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0583__A _1015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1059_ _1059_/A vssd1 vssd1 vccd1 vccd1 _1061_/A sky130_fd_sc_hd__inv_2
X_1128_ _1128_/A _1128_/B vssd1 vssd1 vccd1 vccd1 _1133_/B sky130_fd_sc_hd__and2_1
XFILLER_31_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_59 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput47 _1170_/B vssd1 vssd1 vccd1 vccd1 o_out[13] sky130_fd_sc_hd__buf_2
XFILLER_0_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput58 _1169_/B vssd1 vssd1 vccd1 vccd1 o_out[9] sky130_fd_sc_hd__buf_2
XFILLER_16_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1066__C1 _0866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0668__A _0693_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0607__S _0693_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0628_ _0770_/A vssd1 vssd1 vccd1 vccd1 _0733_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0578__A _0631_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_46 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0810__A2 _0834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input21_A i_mode[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0845__B _0892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_16 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_35 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0786__A1 _0796_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0893_ _0894_/A _0894_/B _0894_/C vssd1 vssd1 vccd1 vccd1 _0895_/A sky130_fd_sc_hd__a21o_1
X_0962_ _1015_/A input3/X vssd1 vssd1 vccd1 vccd1 _0964_/A sky130_fd_sc_hd__nor2_1
XFILLER_4_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_3_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0701__A1 _0693_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0768__A1 _1119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1009__A2 _0834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0940__A1 _0952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output52_A _1167_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1161_ _1161_/A _1161_/B _1161_/C vssd1 vssd1 vccd1 vccd1 _1161_/X sky130_fd_sc_hd__and3_1
X_1092_ _1151_/A _1092_/B vssd1 vssd1 vccd1 vccd1 _1092_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_20_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0876_ _0876_/A _0876_/B vssd1 vssd1 vccd1 vccd1 _0877_/B sky130_fd_sc_hd__nand2_1
X_0945_ _1124_/A _1003_/A vssd1 vssd1 vccd1 vccd1 _0945_/Y sky130_fd_sc_hd__nor2_1
XFILLER_9_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0931__A1 _1119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0586__A _0695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1175__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0989__A1 _1119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0661_ _1099_/S _0661_/B vssd1 vssd1 vccd1 vccd1 _0661_/Y sky130_fd_sc_hd__nor2_1
X_0730_ _1097_/A _0834_/A _0948_/C _0724_/B _0866_/A vssd1 vssd1 vccd1 vccd1 _0730_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_10_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0592_ _0595_/D vssd1 vssd1 vccd1 vccd1 _0747_/A sky130_fd_sc_hd__buf_2
XANTENNA__0868__A1_N _0892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1144_ _1144_/A _1144_/B vssd1 vssd1 vccd1 vccd1 _1146_/A sky130_fd_sc_hd__xnor2_1
X_1075_ _0943_/B _1074_/X _1102_/S vssd1 vssd1 vccd1 vccd1 _1076_/B sky130_fd_sc_hd__mux2_1
XANTENNA__1030__A _1059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0859_ _0878_/A _0858_/X _1073_/A vssd1 vssd1 vccd1 vccd1 _0859_/Y sky130_fd_sc_hd__o21ai_1
X_0928_ _0901_/A _0924_/X _0927_/X vssd1 vssd1 vccd1 vccd1 _0928_/Y sky130_fd_sc_hd__a21oi_1
XANTENNA__1157__A1 _1003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0763__B _0763_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0683__A3 _0952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0954__A _0954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1084__B1 _1119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0673__B input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0644_ _0653_/A _0653_/B vssd1 vssd1 vccd1 vccd1 _0720_/C sky130_fd_sc_hd__nor2_2
X_0713_ _0711_/B _0711_/C _0711_/D _0711_/A vssd1 vssd1 vccd1 vccd1 _0714_/C sky130_fd_sc_hd__a22o_1
XANTENNA__0848__B _0848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0864__A _0894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0583__B _1059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1127_ _1110_/A _0834_/X _0808_/X _1111_/A _0866_/X vssd1 vssd1 vccd1 vccd1 _1128_/B
+ sky130_fd_sc_hd__a221o_1
X_1058_ _1119_/A _1058_/B _1058_/C vssd1 vssd1 vccd1 vccd1 _1077_/A sky130_fd_sc_hd__and3_1
XFILLER_15_16 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xoutput48 _1170_/C vssd1 vssd1 vccd1 vccd1 o_out[14] sky130_fd_sc_hd__buf_2
XFILLER_0_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_148 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1066__B1 _0808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0668__B input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_262 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0627_ _1007_/A _0684_/A vssd1 vssd1 vccd1 vccd1 _0627_/X sky130_fd_sc_hd__and2_1
XFILLER_38_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input14_A i_l[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0679__A _0759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0618__S _0738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0580__C _0595_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input6_A i_l[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0962__A _1015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0961_ _1145_/B vssd1 vssd1 vccd1 vccd1 _1169_/B sky130_fd_sc_hd__inv_2
X_0892_ _0892_/A vssd1 vssd1 vccd1 vccd1 _0894_/B sky130_fd_sc_hd__inv_2
XANTENNA__1017__B input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0710__A2 _0631_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1160_ _1131_/A _0878_/X _1131_/B _0848_/A vssd1 vssd1 vccd1 vccd1 _1161_/C sky130_fd_sc_hd__a31o_1
X_1091_ _1091_/A _1091_/B _1091_/C vssd1 vssd1 vccd1 vccd1 _1092_/B sky130_fd_sc_hd__and3_1
XANTENNA_output45_A _1166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0944_ _1155_/C _0944_/B vssd1 vssd1 vccd1 vccd1 _0944_/Y sky130_fd_sc_hd__nor2_1
X_0875_ _0875_/A _0875_/B vssd1 vssd1 vccd1 vccd1 _0894_/C sky130_fd_sc_hd__nand2_1
XFILLER_18_16 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1175__A2 _1176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0660_ _1099_/S _0661_/B _0747_/B vssd1 vssd1 vccd1 vccd1 _0660_/X sky130_fd_sc_hd__a21o_1
X_0591_ input2/X _0878_/A _0787_/A vssd1 vssd1 vccd1 vccd1 _0600_/B sky130_fd_sc_hd__o21ai_4
XFILLER_6_253 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1143_ _1143_/A _1143_/B vssd1 vssd1 vccd1 vccd1 _1144_/B sky130_fd_sc_hd__xnor2_1
X_1074_ _1000_/Y _1073_/Y _1101_/S vssd1 vssd1 vccd1 vccd1 _1074_/X sky130_fd_sc_hd__mux2_1
X_0927_ _0952_/A _0656_/B _1132_/A _0926_/X vssd1 vssd1 vccd1 vccd1 _0927_/X sky130_fd_sc_hd__a211o_1
XANTENNA__1030__B input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0858_ _0892_/A _0848_/B _0858_/S vssd1 vssd1 vccd1 vccd1 _0858_/X sky130_fd_sc_hd__mux2_1
X_0789_ _0743_/Y _0788_/Y _0919_/A vssd1 vssd1 vccd1 vccd1 _0789_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0597__A _1131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_25 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0840__A1 _0848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1131__A _1131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0712_ _0747_/A _0747_/B vssd1 vssd1 vccd1 vccd1 _0751_/A sky130_fd_sc_hd__nor2_1
X_0643_ _0858_/S vssd1 vssd1 vccd1 vccd1 _1099_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__0898__A1 _0748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1126_ _1126_/A _1161_/A _1126_/C _1126_/D vssd1 vssd1 vccd1 vccd1 _1133_/A sky130_fd_sc_hd__and4_1
XFILLER_40_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0864__B _0892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0583__C _1039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1057_ _1057_/A _1057_/B _1061_/C vssd1 vssd1 vccd1 vccd1 _1058_/C sky130_fd_sc_hd__or3_1
XFILLER_15_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0889__A1 _0925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput49 _1176_/X vssd1 vssd1 vccd1 vccd1 o_out[15] sky130_fd_sc_hd__buf_2
XFILLER_0_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput38 _1171_/Y vssd1 vssd1 vccd1 vccd1 o_flags[0] sky130_fd_sc_hd__buf_2
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0813__A1 _0748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1066__A1 _1086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_71 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0965__A _0975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0626_ _0626_/A vssd1 vssd1 vccd1 vccd1 _1097_/B sky130_fd_sc_hd__buf_2
X_1109_ _1110_/A input8/X vssd1 vssd1 vccd1 vccd1 _1111_/A sky130_fd_sc_hd__nand2_1
XFILLER_42_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0679__B _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0695__A _0695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0634__S _0779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0580__D _0595_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0609_ _0770_/A vssd1 vssd1 vccd1 vccd1 _0781_/A sky130_fd_sc_hd__clkinv_4
XFILLER_26_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0962__B input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0960_ _1119_/A _0938_/Y _0959_/X vssd1 vssd1 vccd1 vccd1 _1145_/B sky130_fd_sc_hd__a21oi_2
X_0891_ _1103_/A _1125_/B _0890_/X vssd1 vssd1 vccd1 vccd1 _0891_/X sky130_fd_sc_hd__o21a_1
XANTENNA__0629__S _0779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_133 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_100 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1090_ _1064_/A _1061_/X _1062_/A vssd1 vssd1 vccd1 vccd1 _1091_/C sky130_fd_sc_hd__a21oi_1
X_0874_ _0905_/A _0874_/B vssd1 vssd1 vccd1 vccd1 _0875_/B sky130_fd_sc_hd__or2_1
XFILLER_13_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0943_ _1102_/S _0943_/B vssd1 vssd1 vccd1 vccd1 _0943_/Y sky130_fd_sc_hd__nand2_1
XFILLER_18_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0793__A _0815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0590_ _0590_/A _1155_/B vssd1 vssd1 vccd1 vccd1 _0787_/A sky130_fd_sc_hd__nand2_2
X_1142_ _1142_/A _1142_/B vssd1 vssd1 vccd1 vccd1 _1143_/B sky130_fd_sc_hd__xnor2_1
XFILLER_1_31 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1073_ _1073_/A _1073_/B vssd1 vssd1 vccd1 vccd1 _1073_/Y sky130_fd_sc_hd__nand2_1
X_0857_ _1119_/A _0876_/B _0857_/C vssd1 vssd1 vccd1 vccd1 _0857_/X sky130_fd_sc_hd__and3_1
X_0926_ _0954_/A _0834_/X _0808_/X _0907_/C vssd1 vssd1 vccd1 vccd1 _0926_/X sky130_fd_sc_hd__a22o_1
XANTENNA__1039__A _1039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0788_ _0878_/A _0786_/X _1073_/A vssd1 vssd1 vccd1 vccd1 _0788_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_45_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0840__A2 _0657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input37_A i_r[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_91 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0711_ _0711_/A _0711_/B _0711_/C _0711_/D vssd1 vssd1 vccd1 vccd1 _0745_/B sky130_fd_sc_hd__and4_1
X_0642_ _0693_/B vssd1 vssd1 vccd1 vccd1 _0858_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__0637__S _0779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1125_ _1125_/A _1125_/B vssd1 vssd1 vccd1 vccd1 _1126_/D sky130_fd_sc_hd__nand2_1
XANTENNA__0583__D _1086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1056_ _1057_/A _1057_/B _1061_/C vssd1 vssd1 vccd1 vccd1 _1058_/B sky130_fd_sc_hd__o21ai_1
XFILLER_21_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0909_ _0909_/A vssd1 vssd1 vccd1 vccd1 _0909_/Y sky130_fd_sc_hd__inv_2
Xoutput39 _1164_/X vssd1 vssd1 vccd1 vccd1 o_flags[1] sky130_fd_sc_hd__buf_2
XFILLER_48_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0889__A2 _0657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1066__A2 _0834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0625_ _0759_/A _0625_/B vssd1 vssd1 vccd1 vccd1 _0626_/A sky130_fd_sc_hd__or2_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1039_ _1039_/A vssd1 vssd1 vccd1 vccd1 _1039_/Y sky130_fd_sc_hd__inv_2
X_1108_ _1108_/A vssd1 vssd1 vccd1 vccd1 _1113_/A sky130_fd_sc_hd__inv_2
XFILLER_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0731__A1 _0763_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0731__B2 _0808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_197 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0608_ _0669_/A _0608_/B vssd1 vssd1 vccd1 vccd1 _0608_/Y sky130_fd_sc_hd__nand2_1
XFILLER_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0890_ _1006_/B _0885_/X _0886_/X _0889_/Y vssd1 vssd1 vccd1 vccd1 _0890_/X sky130_fd_sc_hd__o211a_1
XFILLER_4_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_237 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1120__A1 _1155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0861__A0 _0744_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0873_ _0905_/A _0874_/B vssd1 vssd1 vccd1 vccd1 _0875_/A sky130_fd_sc_hd__nand2_1
XFILLER_9_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0942_ _0880_/Y _0941_/Y _1101_/S vssd1 vssd1 vccd1 vccd1 _0943_/B sky130_fd_sc_hd__mux2_1
XFILLER_18_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0793__B _1131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_277 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1141_ _1167_/A _1167_/B vssd1 vssd1 vccd1 vccd1 _1142_/B sky130_fd_sc_hd__xor2_1
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_43 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_output50_A _1167_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1072_ _0669_/C _0673_/X _0878_/X vssd1 vssd1 vccd1 vccd1 _1073_/B sky130_fd_sc_hd__a21o_1
XANTENNA__1145__A _1169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0856_ _0855_/C _0855_/B _0846_/X vssd1 vssd1 vccd1 vccd1 _0857_/C sky130_fd_sc_hd__a21bo_1
X_0925_ _0925_/A _0925_/B vssd1 vssd1 vccd1 vccd1 _1132_/A sky130_fd_sc_hd__and2_2
X_0787_ _0787_/A vssd1 vssd1 vccd1 vccd1 _1073_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_43_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0894__A _0894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0825__A0 _0848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0761__C1 _0866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0641_ _0720_/A _0653_/B _0653_/A _0747_/A vssd1 vssd1 vccd1 vccd1 _0866_/A sky130_fd_sc_hd__and4bb_2
X_0710_ input2/X _0631_/B input1/X vssd1 vssd1 vccd1 vccd1 _0711_/D sky130_fd_sc_hd__a21o_1
X_1055_ _1055_/A _1055_/B vssd1 vssd1 vccd1 vccd1 _1061_/C sky130_fd_sc_hd__and2_1
XFILLER_18_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1124_ _1124_/A _1124_/B vssd1 vssd1 vccd1 vccd1 _1126_/C sky130_fd_sc_hd__nand2_1
XFILLER_31_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0839_ _0839_/A _0839_/B vssd1 vssd1 vccd1 vccd1 _0839_/Y sky130_fd_sc_hd__nor2_1
X_0908_ _0957_/A _0908_/B vssd1 vssd1 vccd1 vccd1 _0914_/A sky130_fd_sc_hd__nand2_1
XFILLER_0_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0738__S _0738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0624_ _0625_/B vssd1 vssd1 vccd1 vccd1 _1006_/B sky130_fd_sc_hd__buf_2
XFILLER_7_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1038_ input4/X _1038_/B vssd1 vssd1 vccd1 vccd1 _1038_/Y sky130_fd_sc_hd__nor2_1
X_1107_ _1091_/A _1091_/B _1091_/C _1151_/A vssd1 vssd1 vccd1 vccd1 _1115_/B sky130_fd_sc_hd__a31o_1
XFILLER_21_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0731__A2 _0657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_110 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_238 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0607_ input5/X input6/X _0693_/B vssd1 vssd1 vccd1 vccd1 _0608_/B sky130_fd_sc_hd__mux2_1
XFILLER_26_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0796__B _0796_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input12_A i_l[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1058__A _1119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input4_A i_l[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0870__A1 _1103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0941_ _0878_/X _0940_/X _1073_/A vssd1 vssd1 vccd1 vccd1 _0941_/Y sky130_fd_sc_hd__o21ai_1
X_0872_ _0872_/A vssd1 vssd1 vccd1 vccd1 _1165_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1140_ _1167_/C _1167_/D vssd1 vssd1 vccd1 vccd1 _1142_/A sky130_fd_sc_hd__xor2_1
XFILLER_45_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_output43_A _1167_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1071_ _0830_/B _0923_/Y _1070_/X vssd1 vssd1 vccd1 vccd1 _1077_/C sky130_fd_sc_hd__o21ai_1
XFILLER_45_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0924_ _0954_/A _0952_/A _0948_/C _0866_/X vssd1 vssd1 vccd1 vccd1 _0924_/X sky130_fd_sc_hd__a31o_1
X_0786_ _0815_/A _0796_/B _0858_/S vssd1 vssd1 vccd1 vccd1 _0786_/X sky130_fd_sc_hd__mux2_1
X_0855_ _0846_/X _0855_/B _0855_/C vssd1 vssd1 vccd1 vccd1 _0876_/B sky130_fd_sc_hd__nand3b_1
XANTENNA__1011__A1 _0866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0825__A1 _0815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0640_ _0627_/X _0633_/X _1007_/A _0639_/X vssd1 vssd1 vccd1 vccd1 _0640_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__0995__A _1039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1054_ _1086_/A input6/X vssd1 vssd1 vccd1 vccd1 _1055_/B sky130_fd_sc_hd__or2_1
X_1123_ _1003_/A _1002_/B _1122_/X vssd1 vssd1 vccd1 vccd1 _1124_/B sky130_fd_sc_hd__a21o_1
XFILLER_33_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0907_ _0907_/A _0925_/A _0907_/C vssd1 vssd1 vccd1 vccd1 _0908_/B sky130_fd_sc_hd__or3_1
X_0838_ _0884_/A _0684_/Y _0685_/Y _0677_/X _1006_/B vssd1 vssd1 vccd1 vccd1 _0839_/B
+ sky130_fd_sc_hd__a221o_1
X_0769_ _0669_/Y _0674_/Y _0781_/A vssd1 vssd1 vccd1 vccd1 _0769_/X sky130_fd_sc_hd__mux2_1
XFILLER_0_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_144 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0623_ _1130_/A _1131_/C _1131_/A vssd1 vssd1 vccd1 vccd1 _0625_/B sky130_fd_sc_hd__a21o_1
XFILLER_7_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1106_ _1106_/A vssd1 vssd1 vccd1 vccd1 _1115_/A sky130_fd_sc_hd__inv_2
XFILLER_42_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1037_ _1059_/A _0834_/X _0808_/X _1038_/B _1036_/Y vssd1 vssd1 vccd1 vccd1 _1048_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_21_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_206 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0606_ _0669_/A _0606_/B vssd1 vssd1 vccd1 vccd1 _0733_/B sky130_fd_sc_hd__nand2_1
XFILLER_43_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_261 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_13_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0940_ _0975_/B _0952_/A _1099_/S vssd1 vssd1 vccd1 vccd1 _0940_/X sky130_fd_sc_hd__mux2_1
XFILLER_20_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0871_ _1173_/A _0853_/Y _0857_/X _0870_/Y vssd1 vssd1 vccd1 vccd1 _0872_/A sky130_fd_sc_hd__a211o_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_51 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_235 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1087__A2 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1070_ _1097_/A _1097_/B _0672_/X _1069_/Y vssd1 vssd1 vccd1 vccd1 _1070_/X sky130_fd_sc_hd__o31a_1
X_0854_ _0843_/A _0848_/B _0805_/A _0805_/B _0831_/A vssd1 vssd1 vccd1 vccd1 _0855_/B
+ sky130_fd_sc_hd__a221o_1
X_0923_ _0923_/A _1125_/A vssd1 vssd1 vccd1 vccd1 _0923_/Y sky130_fd_sc_hd__nand2_1
X_0785_ _0785_/A vssd1 vssd1 vccd1 vccd1 _1167_/D sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_28_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0589__A1 _0695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0761__A1 _0729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_183 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_72 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0995__B input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1172__A _1173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1122_ _1101_/S _1073_/Y _1120_/X _1121_/Y _1102_/S vssd1 vssd1 vccd1 vccd1 _1122_/X
+ sky130_fd_sc_hd__o221a_1
XFILLER_33_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1053_ _1086_/A input6/X vssd1 vssd1 vccd1 vccd1 _1055_/A sky130_fd_sc_hd__nand2_1
XFILLER_18_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0837_ _1097_/A _0672_/X _1006_/A vssd1 vssd1 vccd1 vccd1 _0839_/A sky130_fd_sc_hd__o21a_1
X_0906_ _0907_/A _0925_/A _0907_/C vssd1 vssd1 vccd1 vccd1 _0957_/A sky130_fd_sc_hd__o21ai_1
X_0768_ _1119_/A _0758_/Y _0762_/X _0767_/Y vssd1 vssd1 vccd1 vccd1 _0784_/A sky130_fd_sc_hd__a211o_1
X_0699_ _0771_/S _0828_/B vssd1 vssd1 vccd1 vccd1 _1003_/A sky130_fd_sc_hd__xnor2_4
XFILLER_24_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input35_A i_r[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_30_101 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1167__A _1167_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0622_ _0720_/A _0747_/A _0653_/A _0653_/B vssd1 vssd1 vccd1 vccd1 _1131_/C sky130_fd_sc_hd__or4b_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1105_ _1118_/B _1084_/Y _1104_/X vssd1 vssd1 vccd1 vccd1 _1170_/C sky130_fd_sc_hd__o21ai_4
X_1036_ _1036_/A _1036_/B vssd1 vssd1 vccd1 vccd1 _1036_/Y sky130_fd_sc_hd__nor2_1
XFILLER_21_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_8_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0605_ input7/X input8/X _0779_/S vssd1 vssd1 vccd1 vccd1 _0606_/B sky130_fd_sc_hd__mux2_1
XFILLER_41_207 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1019_ _1014_/Y _0974_/B _0974_/C _1043_/C _0824_/A vssd1 vssd1 vccd1 vccd1 _1019_/X
+ sky130_fd_sc_hd__a41o_1
XANTENNA__1123__A1 _1003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0634__A0 _0892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0616__A0 _0952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0607__A0 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0870_ _1103_/A _0861_/X _0869_/X vssd1 vssd1 vccd1 vccd1 _0870_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_9_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0999_ _1099_/S input4/X _0675_/X vssd1 vssd1 vccd1 vccd1 _0999_/X sky130_fd_sc_hd__o21a_1
XANTENNA__1085__A input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0802__A _1173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0853_ _0912_/A _0853_/B vssd1 vssd1 vccd1 vccd1 _0853_/Y sky130_fd_sc_hd__xnor2_1
X_0922_ _1124_/A vssd1 vssd1 vccd1 vccd1 _1125_/A sky130_fd_sc_hd__inv_2
X_0784_ _0784_/A _0784_/B _0783_/X vssd1 vssd1 vccd1 vccd1 _0785_/A sky130_fd_sc_hd__or3b_1
XFILLER_36_151 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput1 i_carry vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_2
XFILLER_36_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0737__C1 _0759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1052_ _0985_/S _0993_/Y _0996_/A _0995_/X _1038_/B vssd1 vssd1 vccd1 vccd1 _1057_/B
+ sky130_fd_sc_hd__o311a_1
X_1121_ _0878_/X _0669_/B _1101_/S vssd1 vssd1 vccd1 vccd1 _1121_/Y sky130_fd_sc_hd__o21ai_1
X_0767_ _0824_/A _0767_/B vssd1 vssd1 vccd1 vccd1 _0767_/Y sky130_fd_sc_hd__nor2_1
X_0836_ _0843_/A _0834_/X _0866_/A _0835_/X vssd1 vssd1 vccd1 vccd1 _0836_/X sky130_fd_sc_hd__a211o_1
X_0905_ _0905_/A vssd1 vssd1 vccd1 vccd1 _0907_/A sky130_fd_sc_hd__inv_2
X_0698_ _0878_/A _1007_/B vssd1 vssd1 vccd1 vccd1 _0828_/B sky130_fd_sc_hd__nand2_2
XFILLER_24_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input28_A i_r[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1167__B _1167_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0621_ _0611_/X _0618_/X _1007_/A vssd1 vssd1 vccd1 vccd1 _0621_/X sky130_fd_sc_hd__mux2_1
XFILLER_23_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1035_ _0948_/C _1057_/A _0866_/X vssd1 vssd1 vccd1 vccd1 _1036_/B sky130_fd_sc_hd__a21oi_1
X_1104_ _0824_/A _1092_/Y _1098_/X _1103_/X vssd1 vssd1 vccd1 vccd1 _1104_/X sky130_fd_sc_hd__o211a_1
X_0819_ _0820_/A _1131_/A _0820_/C vssd1 vssd1 vccd1 vccd1 _0821_/A sky130_fd_sc_hd__a21o_1
XFILLER_44_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0652__A1 _0866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0900__A _0954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0891__A1 _1103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0662__A2_N _0657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0604_ _0693_/B vssd1 vssd1 vccd1 vccd1 _0779_/S sky130_fd_sc_hd__buf_4
XFILLER_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0634__A1 _0874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_26_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1018_ _1018_/A _1018_/B vssd1 vssd1 vccd1 vccd1 _1043_/C sky130_fd_sc_hd__nand2_1
XFILLER_43_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0630__A _0693_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_13 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0616__A1 _0975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1041__A1 _1039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0607__A1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input10_A i_l[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1099__A1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0625__A _0759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0773__A0 _0796_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0998_ _0985_/S _0993_/Y _1017_/C _1119_/A vssd1 vssd1 vccd1 vccd1 _0998_/X sky130_fd_sc_hd__o31a_1
XANTENNA_input2_A i_l[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_18_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0921_ _0789_/X _0920_/X _1102_/S vssd1 vssd1 vccd1 vccd1 _0921_/X sky130_fd_sc_hd__mux2_1
X_0783_ _1103_/A _1003_/A _1004_/A vssd1 vssd1 vccd1 vccd1 _0783_/X sky130_fd_sc_hd__or3_1
X_0852_ _0800_/A _0850_/Y _0909_/A vssd1 vssd1 vccd1 vccd1 _0853_/B sky130_fd_sc_hd__a21o_1
XFILLER_5_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput2 i_l[0] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_2
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_163 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_56 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0985__A0 _0808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0737__B1 _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1051_ _1051_/A vssd1 vssd1 vccd1 vccd1 _1170_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1120_ _1155_/A _0590_/A _1155_/B vssd1 vssd1 vccd1 vccd1 _1120_/X sky130_fd_sc_hd__o21a_1
XFILLER_33_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0904_ _0907_/C _0936_/A vssd1 vssd1 vccd1 vccd1 _0904_/Y sky130_fd_sc_hd__xnor2_1
X_0766_ _0764_/A _0764_/X _0766_/S vssd1 vssd1 vccd1 vccd1 _0767_/B sky130_fd_sc_hd__mux2_1
X_0835_ _0729_/A _0808_/A _0835_/S vssd1 vssd1 vccd1 vccd1 _0835_/X sky130_fd_sc_hd__mux2_1
X_0697_ _0923_/A _1124_/A vssd1 vssd1 vccd1 vccd1 _1103_/A sky130_fd_sc_hd__nand2_4
XANTENNA__0707__B input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0723__A _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_46_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_125 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1167__C _1167_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0779__S _0779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0620_ _0763_/A vssd1 vssd1 vccd1 vccd1 _1007_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0808__A _0808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1034_ _1038_/B _1034_/B vssd1 vssd1 vccd1 vccd1 _1034_/X sky130_fd_sc_hd__xor2_1
X_1103_ _1103_/A _1103_/B vssd1 vssd1 vccd1 vccd1 _1103_/X sky130_fd_sc_hd__or2_1
XANTENNA__0949__B1 _1132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0749_ _1103_/A _1003_/A _0744_/X _0746_/Y _0748_/X vssd1 vssd1 vccd1 vccd1 _0750_/B
+ sky130_fd_sc_hd__o32a_1
X_0818_ _0855_/C _0835_/S vssd1 vssd1 vccd1 vccd1 _0820_/C sky130_fd_sc_hd__nand2_1
XFILLER_44_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0900__B _0952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0603_ _0603_/A _0603_/B _0603_/C vssd1 vssd1 vccd1 vccd1 _0669_/A sky130_fd_sc_hd__nor3_4
XANTENNA__0867__C1 _0866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1017_ _1017_/A input3/X _1017_/C vssd1 vssd1 vccd1 vccd1 _1018_/B sky130_fd_sc_hd__or3_1
XFILLER_32_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_246 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_9_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0816__A _0843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0773__A1 _0815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0997_ _0985_/S _0993_/Y _1017_/C vssd1 vssd1 vccd1 vccd1 _0997_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0819__A2 _1131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0636__A _0816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0920_ _0859_/Y _0918_/Y _1101_/S vssd1 vssd1 vccd1 vccd1 _0920_/X sky130_fd_sc_hd__mux2_1
X_0851_ _0799_/B _0821_/A _0821_/B vssd1 vssd1 vccd1 vccd1 _0909_/A sky130_fd_sc_hd__a21boi_1
X_0782_ _0944_/B _0780_/Y _0919_/A vssd1 vssd1 vccd1 vccd1 _1004_/A sky130_fd_sc_hd__mux2_1
XFILLER_46_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput3 i_l[10] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__buf_2
XFILLER_51_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_68 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0737__A1 _0738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0985__A1 _0948_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1050_ _0923_/A _1024_/Y _1029_/Y _1049_/X vssd1 vssd1 vccd1 vccd1 _1051_/A sky130_fd_sc_hd__a31o_1
X_0834_ _0834_/A vssd1 vssd1 vccd1 vccd1 _0834_/X sky130_fd_sc_hd__clkbuf_4
X_0903_ _0876_/A _0876_/B _0875_/A _0902_/Y vssd1 vssd1 vccd1 vccd1 _0936_/A sky130_fd_sc_hd__a31o_1
X_0765_ _0781_/A _0703_/B _0746_/A _0725_/X vssd1 vssd1 vccd1 vccd1 _0766_/S sky130_fd_sc_hd__a211o_1
X_0696_ _0886_/A _0696_/B vssd1 vssd1 vccd1 vccd1 _1124_/A sky130_fd_sc_hd__xnor2_4
XFILLER_24_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0723__B _0763_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1167__D _1167_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1102_ _0980_/X _1101_/X _1102_/S vssd1 vssd1 vccd1 vccd1 _1103_/B sky130_fd_sc_hd__mux2_1
XANTENNA__0824__A _0824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1033_ _0985_/S _0993_/Y _0996_/A _0995_/X vssd1 vssd1 vccd1 vccd1 _1034_/B sky130_fd_sc_hd__o31a_1
XFILLER_21_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0817_ _0843_/A _0848_/B vssd1 vssd1 vccd1 vccd1 _0835_/S sky130_fd_sc_hd__nand2_1
XANTENNA__0949__A1 _0975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0748_ _0748_/A vssd1 vssd1 vccd1 vccd1 _0748_/X sky130_fd_sc_hd__buf_2
X_0679_ _0759_/A _0771_/S vssd1 vssd1 vccd1 vccd1 _0884_/A sky130_fd_sc_hd__nor2_1
XFILLER_44_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0637__A0 _0815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_248 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_input33_A i_r[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0602_ _0843_/A _0954_/A _0975_/A vssd1 vssd1 vccd1 vccd1 _0603_/C sky130_fd_sc_hd__or3_1
XFILLER_26_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1016_ _1017_/A input3/X _1017_/C vssd1 vssd1 vccd1 vccd1 _1018_/A sky130_fd_sc_hd__o21ai_1
XANTENNA__0729__A _0729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0858__A0 _0892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1035__B1 _0866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_166 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0816__B _0816_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0996_ _0996_/A _0995_/X vssd1 vssd1 vccd1 vccd1 _1017_/C sky130_fd_sc_hd__nor2b_1
XANTENNA__0773__A2 _0848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0978__S _1099_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0850_ _0913_/A _0913_/B vssd1 vssd1 vccd1 vccd1 _0850_/Y sky130_fd_sc_hd__nor2_1
X_0781_ _0781_/A _0781_/B vssd1 vssd1 vccd1 vccd1 _0919_/A sky130_fd_sc_hd__xnor2_4
XFILLER_39_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput4 i_l[11] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_4
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0979_ _0878_/X _0978_/X _1073_/A vssd1 vssd1 vccd1 vccd1 _0979_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_10_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_146 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0833_ _0820_/C _0831_/Y _0832_/Y vssd1 vssd1 vccd1 vccd1 _0841_/C sky130_fd_sc_hd__o21a_1
X_0902_ _0905_/A _0925_/A vssd1 vssd1 vccd1 vccd1 _0902_/Y sky130_fd_sc_hd__nor2_1
X_0764_ _0764_/A _0764_/B vssd1 vssd1 vccd1 vccd1 _0764_/X sky130_fd_sc_hd__xor2_1
X_0695_ _0695_/A _0886_/B vssd1 vssd1 vccd1 vccd1 _0696_/B sky130_fd_sc_hd__nand2_1
XANTENNA__0967__A2 _0975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1135__A2 _0656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1032_ _1036_/A _1057_/A vssd1 vssd1 vccd1 vccd1 _1038_/B sky130_fd_sc_hd__nor2_2
X_1101_ _1026_/Y _1100_/Y _1101_/S vssd1 vssd1 vccd1 vccd1 _1101_/X sky130_fd_sc_hd__mux2_1
XFILLER_21_127 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0747_ _0747_/A _0747_/B vssd1 vssd1 vccd1 vccd1 _0748_/A sky130_fd_sc_hd__or2_1
X_0816_ _0843_/A _0816_/B vssd1 vssd1 vccd1 vccd1 _0855_/C sky130_fd_sc_hd__or2_1
XANTENNA__0949__A2 _0656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1071__A1 _0830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0678_ _0672_/X _0677_/X _1007_/A vssd1 vssd1 vccd1 vccd1 _0950_/B sky130_fd_sc_hd__mux2_1
XANTENNA__0637__A1 _0848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input26_A i_r[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0925__A _0925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0601_ _0759_/A vssd1 vssd1 vccd1 vccd1 _0886_/A sky130_fd_sc_hd__clkinv_2
XFILLER_7_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0867__A1 _0808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1015_ _1015_/A vssd1 vssd1 vccd1 vccd1 _1017_/A sky130_fd_sc_hd__inv_2
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0858__A1 _0848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1035__A1 _0948_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output57_A _1169_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0995_ _1039_/A input4/X vssd1 vssd1 vccd1 vccd1 _0995_/X sky130_fd_sc_hd__or2_1
XANTENNA__0773__A3 _0892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0930__B1 _1103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0780_ _0878_/A _0779_/X _0787_/A vssd1 vssd1 vccd1 vccd1 _0780_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__0933__A _0975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_111 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput5 i_l[12] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__buf_2
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0843__A _0843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0978_ input3/X _0975_/B _1099_/S vssd1 vssd1 vccd1 vccd1 _0978_/X sky130_fd_sc_hd__mux2_1
XFILLER_10_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0753__A _0759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0763_ _0763_/A _0763_/B vssd1 vssd1 vccd1 vccd1 _0764_/B sky130_fd_sc_hd__or2_1
X_0832_ _0820_/C _0831_/Y _0748_/X vssd1 vssd1 vccd1 vccd1 _0832_/Y sky130_fd_sc_hd__a21oi_1
X_0901_ _0901_/A _0937_/A vssd1 vssd1 vccd1 vccd1 _0907_/C sky130_fd_sc_hd__and2_1
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0897__C1 _0824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0694_ _0771_/S _1007_/B vssd1 vssd1 vccd1 vccd1 _0886_/B sky130_fd_sc_hd__or2_1
XANTENNA__1129__B1 _0656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_14 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_21_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1031_ _1059_/A input5/X vssd1 vssd1 vccd1 vccd1 _1057_/A sky130_fd_sc_hd__and2_1
X_1100_ _0878_/X _1099_/X _1073_/A vssd1 vssd1 vccd1 vccd1 _1100_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_21_139 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput30 i_r[2] vssd1 vssd1 vccd1 vccd1 _0771_/S sky130_fd_sc_hd__buf_4
X_0746_ _0746_/A _0746_/B vssd1 vssd1 vccd1 vccd1 _0746_/Y sky130_fd_sc_hd__xnor2_1
X_0815_ _0815_/A vssd1 vssd1 vccd1 vccd1 _0820_/A sky130_fd_sc_hd__inv_2
X_0677_ _0674_/Y _0676_/Y _0738_/S vssd1 vssd1 vccd1 vccd1 _0677_/X sky130_fd_sc_hd__mux2_1
XFILLER_37_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_161 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input19_A i_mode[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0600_ _1131_/B _0600_/B _0923_/A vssd1 vssd1 vccd1 vccd1 _0665_/A sky130_fd_sc_hd__or3b_1
XFILLER_14_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_34_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1014_ _1014_/A vssd1 vssd1 vccd1 vccd1 _1014_/Y sky130_fd_sc_hd__inv_2
X_0729_ _0729_/A vssd1 vssd1 vccd1 vccd1 _0948_/C sky130_fd_sc_hd__clkbuf_4
XFILLER_43_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0671__A _0733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0776__A1 _0781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0666__A _0759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0994_ _1039_/A input4/X vssd1 vssd1 vccd1 vccd1 _0996_/A sky130_fd_sc_hd__and2_1
XANTENNA__0605__S _0779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0749__A1 _1103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0749__B2 _0748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1110__A _1110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput6 i_l[13] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__clkbuf_4
X_0977_ _0992_/A _0977_/B vssd1 vssd1 vccd1 vccd1 _0977_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_19_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0753__B _0796_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0900_ _0954_/A _0952_/A vssd1 vssd1 vccd1 vccd1 _0937_/A sky130_fd_sc_hd__nand2_2
X_0762_ _0796_/B _0657_/X _0754_/B _0761_/X vssd1 vssd1 vccd1 vccd1 _0762_/X sky130_fd_sc_hd__a22o_1
X_0831_ _0831_/A _0831_/B vssd1 vssd1 vccd1 vccd1 _0831_/Y sky130_fd_sc_hd__nor2_1
X_0693_ _0770_/A _0693_/B vssd1 vssd1 vccd1 vccd1 _1007_/B sky130_fd_sc_hd__or2_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1015__A _1015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1176_ _1176_/A vssd1 vssd1 vccd1 vccd1 _1176_/X sky130_fd_sc_hd__clkbuf_1
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1129__A1 _1110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0658__B input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0939__A _1003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0879__A0 _0925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1030_ _1059_/A input5/X vssd1 vssd1 vccd1 vccd1 _1036_/A sky130_fd_sc_hd__nor2_1
Xinput31 i_r[3] vssd1 vssd1 vccd1 vccd1 _0759_/A sky130_fd_sc_hd__buf_2
Xinput20 i_mode[2] vssd1 vssd1 vccd1 vccd1 _0653_/A sky130_fd_sc_hd__clkbuf_2
X_0814_ _1103_/A _1024_/B _0802_/Y _0813_/X vssd1 vssd1 vccd1 vccd1 _1168_/A sky130_fd_sc_hd__o211ai_2
XFILLER_14_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0745_ _0745_/A _0745_/B vssd1 vssd1 vccd1 vccd1 _0746_/B sky130_fd_sc_hd__or2_1
X_0676_ _0858_/S _0975_/B _0684_/A _0675_/X vssd1 vssd1 vccd1 vccd1 _0676_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_37_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1159_ _1131_/B _0600_/B _0598_/B vssd1 vssd1 vccd1 vccd1 _1161_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__0584__A _0894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1047__B1 _0824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_173 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0759__A _0759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0730__C1 _0866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1013_ _0923_/A _1005_/X _1012_/X vssd1 vssd1 vccd1 vccd1 _1013_/X sky130_fd_sc_hd__a21o_1
XFILLER_19_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0659_ _0720_/A _0720_/C vssd1 vssd1 vccd1 vccd1 _0747_/B sky130_fd_sc_hd__nand2_1
X_0728_ _0771_/S vssd1 vssd1 vccd1 vccd1 _1097_/A sky130_fd_sc_hd__clkbuf_4
XANTENNA__0579__A _0759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_14 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input31_A i_r[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0952__A _0952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0671__B _1155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_38 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1108__A _1108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0682__A _0874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0993_ _0937_/A _0937_/B _0935_/A _0975_/Y _0992_/Y vssd1 vssd1 vccd1 vccd1 _0993_/Y
+ sky130_fd_sc_hd__a311oi_4
XFILLER_39_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0857__A _1119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0749__A2 _1003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0592__A _0595_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0767__A _0824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1110__B input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput7 i_l[14] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__0616__S _0779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0976_ _0937_/A _0937_/B _0935_/A _0975_/Y vssd1 vssd1 vccd1 vccd1 _0977_/B sky130_fd_sc_hd__a31o_1
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_19_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_69 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0830_ _1103_/A _0830_/B vssd1 vssd1 vccd1 vccd1 _0841_/B sky130_fd_sc_hd__nor2_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0761_ _0729_/A _0759_/X _0760_/X _0866_/A vssd1 vssd1 vccd1 vccd1 _0761_/X sky130_fd_sc_hd__a211o_1
XFILLER_41_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0692_ _1155_/C _0944_/B vssd1 vssd1 vccd1 vccd1 _0692_/X sky130_fd_sc_hd__or2_1
XFILLER_49_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_260 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1175_ input8/X _1176_/A _1172_/Y _1173_/X _1174_/Y vssd1 vssd1 vccd1 vccd1 _1175_/X
+ sky130_fd_sc_hd__o2111a_1
XANTENNA__1031__A _1059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0959_ _0923_/A _0946_/X _0951_/X _0958_/X vssd1 vssd1 vccd1 vccd1 _0959_/X sky130_fd_sc_hd__a211o_1
XFILLER_21_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1129__A2 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0879__A1 _0892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0813_ _0748_/X _0831_/B _0805_/Y _0812_/X vssd1 vssd1 vccd1 vccd1 _0813_/X sky130_fd_sc_hd__o31a_1
Xinput21 i_mode[3] vssd1 vssd1 vccd1 vccd1 _0653_/B sky130_fd_sc_hd__buf_2
Xinput32 i_r[4] vssd1 vssd1 vccd1 vccd1 _1131_/A sky130_fd_sc_hd__clkbuf_4
Xinput10 i_l[2] vssd1 vssd1 vccd1 vccd1 _0763_/B sky130_fd_sc_hd__buf_2
X_0744_ _0600_/B _0671_/Y _1155_/C _0743_/Y vssd1 vssd1 vccd1 vccd1 _0744_/X sky130_fd_sc_hd__o22a_1
X_0675_ _1155_/A input3/X vssd1 vssd1 vccd1 vccd1 _0675_/X sky130_fd_sc_hd__or2_1
XFILLER_37_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0584__B _0905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1158_ _1124_/A _0921_/X _1157_/X vssd1 vssd1 vccd1 vccd1 _1158_/Y sky130_fd_sc_hd__o21ai_1
X_1089_ _1089_/A vssd1 vssd1 vccd1 vccd1 _1151_/A sky130_fd_sc_hd__inv_2
XFILLER_20_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0759__B _0796_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0730__B1 _0948_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_233 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1012_ _1006_/Y _1008_/Y _1011_/X vssd1 vssd1 vccd1 vccd1 _1012_/X sky130_fd_sc_hd__a21o_1
XFILLER_34_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0727_ _0746_/A _0727_/B vssd1 vssd1 vccd1 vccd1 _0727_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_8_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0658_ input2/X input1/X vssd1 vssd1 vccd1 vccd1 _0661_/B sky130_fd_sc_hd__xor2_1
XANTENNA__0579__B _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0589_ _0695_/A _0587_/X _0586_/B _0770_/C vssd1 vssd1 vccd1 vccd1 _1155_/B sky130_fd_sc_hd__a211o_1
XFILLER_27_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_26 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_25_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0779__A0 _0796_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input24_A i_r[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_38_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0924__B1 _0866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0963__A _1015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0992_ _0992_/A vssd1 vssd1 vccd1 vccd1 _0992_/Y sky130_fd_sc_hd__inv_2
XFILLER_39_177 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0873__A _0905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0749__A3 _0744_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0783__A _1103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1095__C1 _1132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1119__A _1119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput8 i_l[15] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_output55_A _1165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0958__A _1173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0676__A2 _0975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0975_ _0975_/A _0975_/B vssd1 vssd1 vccd1 vccd1 _0975_/Y sky130_fd_sc_hd__nor2_1
XFILLER_10_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1010__C1 _1132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_279 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1068__C1 _1132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0760_ _0759_/A _0834_/A _0808_/A _0754_/A vssd1 vssd1 vccd1 vccd1 _0760_/X sky130_fd_sc_hd__a22o_1
XFILLER_41_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0688__A _0779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0691_ _0787_/A _0691_/B vssd1 vssd1 vccd1 vccd1 _0944_/B sky130_fd_sc_hd__nand2_1
XFILLER_49_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1174_ input8/X _1174_/B vssd1 vssd1 vccd1 vccd1 _1174_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_85 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1031__B input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0889_ _0925_/A _0657_/X _0875_/B _0887_/X _0888_/X vssd1 vssd1 vccd1 vccd1 _0889_/Y
+ sky130_fd_sc_hd__a221oi_1
X_0958_ _1173_/A _0972_/A _0972_/B vssd1 vssd1 vccd1 vccd1 _0958_/X sky130_fd_sc_hd__and3_1
XANTENNA__0680__S1 _0733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1129__A3 _0948_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0598__A _0843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1132__A _1132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0812_ _1006_/B _0806_/X _0807_/X _0809_/Y _0811_/X vssd1 vssd1 vccd1 vccd1 _0812_/X
+ sky130_fd_sc_hd__o311a_1
Xinput11 i_l[3] vssd1 vssd1 vccd1 vccd1 _0796_/B sky130_fd_sc_hd__buf_2
X_0743_ _0878_/A _0742_/X _0787_/A vssd1 vssd1 vccd1 vccd1 _0743_/Y sky130_fd_sc_hd__o21ai_1
Xinput33 i_r[5] vssd1 vssd1 vccd1 vccd1 _0843_/A sky130_fd_sc_hd__clkbuf_4
Xinput22 i_r[0] vssd1 vssd1 vccd1 vccd1 _0631_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_0674_ _0779_/S input4/X _0669_/A _0673_/X vssd1 vssd1 vccd1 vccd1 _0674_/Y sky130_fd_sc_hd__o211ai_1
XFILLER_37_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0584__C _1108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1157_ _1003_/A _1027_/X _1156_/X _1125_/A vssd1 vssd1 vccd1 vccd1 _1157_/X sky130_fd_sc_hd__a211o_1
XFILLER_32_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1088_ _1086_/A _1085_/Y _1106_/A vssd1 vssd1 vccd1 vccd1 _1089_/A sky130_fd_sc_hd__a21oi_1
XFILLER_20_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_186 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_22_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0966__A _0975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1011_ _0866_/X _0995_/X _1009_/X _1010_/X vssd1 vssd1 vccd1 vccd1 _1011_/X sky130_fd_sc_hd__a211o_1
XFILLER_34_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0726_ _0738_/S _0703_/B _0725_/X vssd1 vssd1 vccd1 vccd1 _0727_/B sky130_fd_sc_hd__a21oi_1
XFILLER_8_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0657_ _0657_/A vssd1 vssd1 vccd1 vccd1 _0657_/X sky130_fd_sc_hd__buf_2
X_0588_ input8/X vssd1 vssd1 vccd1 vccd1 _0770_/C sky130_fd_sc_hd__clkinv_2
XANTENNA__0960__A1 _1119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0779__A1 _0763_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input17_A i_l[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0709_ _0733_/A input9/X vssd1 vssd1 vccd1 vccd1 _0711_/C sky130_fd_sc_hd__nand2_1
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_input9_A i_l[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0924__A1 _0954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0963__B input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1140__A _1167_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0991_ _0991_/A vssd1 vssd1 vccd1 vccd1 _1166_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__0612__A0 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0873__B _0874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0783__B _1003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput9 i_l[1] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_4
XANTENNA_output48_A _1170_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0974__A _1173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0693__B _0693_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0974_ _1173_/A _0974_/B _0974_/C vssd1 vssd1 vccd1 vccd1 _0974_/X sky130_fd_sc_hd__and3_1
XFILLER_35_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_137 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0794__A _0815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_151 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0690_ _1155_/A input9/X _0878_/A _0646_/X vssd1 vssd1 vccd1 vccd1 _0691_/B sky130_fd_sc_hd__a211o_1
XANTENNA__0688__B _0695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1173_ _1173_/A _1173_/B vssd1 vssd1 vccd1 vccd1 _1173_/X sky130_fd_sc_hd__or2_1
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_24_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0888_ _0905_/A _0925_/A _0948_/C vssd1 vssd1 vccd1 vccd1 _0888_/X sky130_fd_sc_hd__and3_1
X_0957_ _0957_/A _0957_/B _0957_/C _1042_/A vssd1 vssd1 vccd1 vccd1 _0972_/B sky130_fd_sc_hd__nand4_1
XFILLER_21_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput23 i_r[10] vssd1 vssd1 vccd1 vccd1 _1015_/A sky130_fd_sc_hd__buf_2
X_0811_ _0811_/A _0810_/X vssd1 vssd1 vccd1 vccd1 _0811_/X sky130_fd_sc_hd__or2b_1
X_0742_ _0763_/B input9/X _0858_/S vssd1 vssd1 vccd1 vccd1 _0742_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0699__A _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput12 i_l[4] vssd1 vssd1 vccd1 vccd1 _0815_/A sky130_fd_sc_hd__clkbuf_4
Xinput34 i_r[6] vssd1 vssd1 vccd1 vccd1 _0894_/A sky130_fd_sc_hd__buf_2
X_0673_ _1155_/A input5/X vssd1 vssd1 vccd1 vccd1 _0673_/X sky130_fd_sc_hd__or2_1
XFILLER_42_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1087_ _1086_/Y input6/X _1085_/B vssd1 vssd1 vccd1 vccd1 _1106_/A sky130_fd_sc_hd__o21a_1
XANTENNA__0584__D _1110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1156_ _1101_/S _1100_/Y _1155_/X _1102_/S vssd1 vssd1 vccd1 vccd1 _1156_/X sky130_fd_sc_hd__o211a_1
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0730__A2 _0834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_232 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1010_ input4/X _0656_/B _0996_/A _0948_/C _1132_/A vssd1 vssd1 vccd1 vccd1 _1010_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_19_265 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0725_ input9/X _0725_/B vssd1 vssd1 vccd1 vccd1 _0725_/X sky130_fd_sc_hd__and2_1
X_0656_ _0925_/B _0656_/B vssd1 vssd1 vccd1 vccd1 _0657_/A sky130_fd_sc_hd__or2_1
XANTENNA__0579__D _0693_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0595__C _0595_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1053__A _1086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0587_ _1131_/A _1131_/B _0843_/A _0975_/A vssd1 vssd1 vccd1 vccd1 _0587_/X sky130_fd_sc_hd__a211o_1
X_1139_ _1168_/A _1168_/B vssd1 vssd1 vccd1 vccd1 _1143_/A sky130_fd_sc_hd__xor2_1
XFILLER_43_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0892__A _0892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1138__A _1165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0708_ _0733_/A _0834_/A _0729_/A _0745_/A _0866_/A vssd1 vssd1 vccd1 vccd1 _0708_/X
+ sky130_fd_sc_hd__a221o_1
X_0639_ _0635_/Y _0736_/B _0738_/S vssd1 vssd1 vccd1 vccd1 _0639_/X sky130_fd_sc_hd__mux2_1
XANTENNA__1048__A _1132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0924__A2 _0952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1140__B _1167_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0990_ input3/X _0656_/B _0974_/X _0989_/X vssd1 vssd1 vccd1 vccd1 _0991_/A sky130_fd_sc_hd__a211o_1
XFILLER_12_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0612__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0906__A2 _0925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1095__B2 _0948_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0973_ _0972_/A _0972_/B _1043_/B _1043_/A vssd1 vssd1 vccd1 vccd1 _0974_/C sky130_fd_sc_hd__a31o_1
XANTENNA__1010__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1010__B2 _0948_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0760__B1 _0808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0794__B _1131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1068__B2 _0948_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1068__A1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1172_ _1173_/A _1173_/B vssd1 vssd1 vccd1 vccd1 _1172_/Y sky130_fd_sc_hd__nand2_1
XFILLER_2_65 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0956_ _0957_/A _0957_/B _0957_/C _1042_/A vssd1 vssd1 vccd1 vccd1 _0972_/A sky130_fd_sc_hd__a31o_1
X_0887_ _0905_/A _0834_/X _0808_/X _0875_/A _0866_/X vssd1 vssd1 vccd1 vccd1 _0887_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_46_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0742__A0 _0763_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0810_ _1131_/A _0834_/A _0729_/A _0831_/A _0866_/A vssd1 vssd1 vccd1 vccd1 _0810_/X
+ sky130_fd_sc_hd__a221o_1
Xinput13 i_l[5] vssd1 vssd1 vccd1 vccd1 _0816_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_14_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput35 i_r[7] vssd1 vssd1 vccd1 vccd1 _0905_/A sky130_fd_sc_hd__clkbuf_4
X_0741_ _0824_/A _0727_/Y _0732_/Y _0740_/X vssd1 vssd1 vccd1 vccd1 _0750_/A sky130_fd_sc_hd__o211a_1
X_0672_ _0733_/A _0669_/Y _1131_/D _0671_/Y vssd1 vssd1 vccd1 vccd1 _0672_/X sky130_fd_sc_hd__o22a_1
Xinput24 i_r[11] vssd1 vssd1 vccd1 vccd1 _1039_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1086_ _1086_/A vssd1 vssd1 vccd1 vccd1 _1086_/Y sky130_fd_sc_hd__inv_2
X_1155_ _1155_/A _1155_/B _1155_/C vssd1 vssd1 vccd1 vccd1 _1155_/X sky130_fd_sc_hd__or3_1
XFILLER_32_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0939_ _1003_/A _0939_/B vssd1 vssd1 vccd1 vccd1 _0939_/Y sky130_fd_sc_hd__nand2_1
XFILLER_20_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0715__B1 _0657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_247 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0724_ _0724_/A _0724_/B vssd1 vssd1 vccd1 vccd1 _0746_/A sky130_fd_sc_hd__nor2_2
X_0655_ _0653_/C _0720_/C _0654_/X vssd1 vssd1 vccd1 vccd1 _0656_/B sky130_fd_sc_hd__a21o_4
XFILLER_6_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0586_ _0695_/A _0586_/B vssd1 vssd1 vccd1 vccd1 _0590_/A sky130_fd_sc_hd__or2_1
XANTENNA__0595__D _0595_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1053__B input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1138_ _1165_/A _1165_/B vssd1 vssd1 vccd1 vccd1 _1144_/A sky130_fd_sc_hd__xor2_1
X_1069_ _1055_/B _1066_/X _1068_/X vssd1 vssd1 vccd1 vccd1 _1069_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0927__B1 _1132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0707_ _0770_/A input9/X vssd1 vssd1 vccd1 vccd1 _0745_/A sky130_fd_sc_hd__and2_1
XFILLER_30_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0638_ _0684_/A _0638_/B vssd1 vssd1 vccd1 vccd1 _0736_/B sky130_fd_sc_hd__nand2_1
XFILLER_13_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0924__A3 _0948_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input22_A i_r[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1059__A _1059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1095__A2 _0656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0601__A _0759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0972_ _0972_/A _0972_/B _1043_/A _1043_/B vssd1 vssd1 vccd1 vccd1 _0974_/B sky130_fd_sc_hd__nand4_1
XANTENNA__1010__A2 _0656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1061__B input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0683__S1 _0733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0760__A1 _0759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1068__A2 _0656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1171_ _1171_/A _1171_/B _1171_/C _1171_/D vssd1 vssd1 vccd1 vccd1 _1171_/Y sky130_fd_sc_hd__nor4_1
XFILLER_49_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0886_ _0886_/A _0886_/B _1006_/B _1131_/D vssd1 vssd1 vccd1 vccd1 _0886_/X sky130_fd_sc_hd__or4_1
X_0955_ _0955_/A _0954_/Y vssd1 vssd1 vccd1 vccd1 _1042_/A sky130_fd_sc_hd__or2b_1
XANTENNA__0940__S _1099_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0742__A1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0990__A1 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_153 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
Xinput36 i_r[8] vssd1 vssd1 vccd1 vccd1 _0954_/A sky130_fd_sc_hd__buf_2
Xinput14 i_l[6] vssd1 vssd1 vccd1 vccd1 _0892_/A sky130_fd_sc_hd__clkbuf_4
X_0740_ _1006_/A _0984_/B _0739_/X _1006_/B vssd1 vssd1 vccd1 vccd1 _0740_/X sky130_fd_sc_hd__a211o_1
Xinput25 i_r[12] vssd1 vssd1 vccd1 vccd1 _1059_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0868__A2_N _0657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0671_ _0733_/A _1155_/A vssd1 vssd1 vccd1 vccd1 _0671_/Y sky130_fd_sc_hd__nand2_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1154_ _1114_/A _1152_/X _1153_/X _0770_/C _1110_/A vssd1 vssd1 vccd1 vccd1 _1154_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_37_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1085_ input6/X _1085_/B vssd1 vssd1 vccd1 vccd1 _1085_/Y sky130_fd_sc_hd__nor2_1
XFILLER_20_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0869_ _1006_/B _0862_/X _0863_/X _0868_/X vssd1 vssd1 vccd1 vccd1 _0869_/X sky130_fd_sc_hd__o31a_1
XANTENNA__1067__A _1086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0938_ _0954_/C _0938_/B vssd1 vssd1 vccd1 vccd1 _0938_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__0715__A1 _0808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0715__B2 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0723_ _0771_/S _0763_/B vssd1 vssd1 vccd1 vccd1 _0724_/B sky130_fd_sc_hd__and2_1
X_0654_ _0720_/A _0595_/D _0653_/A _0653_/B vssd1 vssd1 vccd1 vccd1 _0654_/X sky130_fd_sc_hd__o211a_1
XFILLER_6_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0585_ _0954_/A _0975_/A _0603_/A _0603_/B vssd1 vssd1 vccd1 vccd1 _0586_/B sky130_fd_sc_hd__or4_1
X_1137_ _1170_/A _1170_/B vssd1 vssd1 vccd1 vccd1 _1149_/A sky130_fd_sc_hd__xor2_1
XFILLER_40_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1068_ input6/X _0656_/B _1067_/X _0948_/C _1132_/A vssd1 vssd1 vccd1 vccd1 _1068_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_16_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0604__A _0693_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0927__A1 _0952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1104__A1 _0824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_292 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0706_ _0770_/A input9/X vssd1 vssd1 vccd1 vccd1 _0711_/B sky130_fd_sc_hd__or2_1
XFILLER_38_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0637_ _0815_/A _0848_/B _0779_/S vssd1 vssd1 vccd1 vccd1 _0638_/B sky130_fd_sc_hd__mux2_1
XANTENNA__1080__A _1108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input15_A i_l[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_77 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1165__A _1165_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0836__B1 _0866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_17 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input7_A i_l[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_258 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0971_ _0971_/A vssd1 vssd1 vccd1 vccd1 _1043_/B sky130_fd_sc_hd__inv_2
XFILLER_4_291 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_50_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0702__A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0760__A2 _0834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1170_ _1170_/A _1170_/B _1170_/C _1176_/A vssd1 vssd1 vccd1 vccd1 _1171_/D sky130_fd_sc_hd__or4_1
X_0885_ _1006_/A _1007_/A _0769_/X _0884_/Y vssd1 vssd1 vccd1 vccd1 _0885_/X sky130_fd_sc_hd__o31a_1
X_0954_ _0954_/A _0954_/B _0954_/C vssd1 vssd1 vccd1 vccd1 _0954_/Y sky130_fd_sc_hd__nand3_1
XANTENNA__0990__A2 _0656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_279 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput15 i_l[7] vssd1 vssd1 vccd1 vccd1 _0874_/B sky130_fd_sc_hd__clkbuf_2
Xinput26 i_r[13] vssd1 vssd1 vccd1 vccd1 _1086_/A sky130_fd_sc_hd__buf_2
X_0670_ input8/X _0684_/A vssd1 vssd1 vccd1 vccd1 _1131_/D sky130_fd_sc_hd__nand2_1
Xinput37 i_r[9] vssd1 vssd1 vccd1 vccd1 _0975_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1153_ _1106_/A _1114_/B _1152_/D _1091_/C vssd1 vssd1 vccd1 vccd1 _1153_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__1173__A _1173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1084_ _1085_/B _1083_/X _1119_/A vssd1 vssd1 vccd1 vccd1 _1084_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__0660__A1 _1099_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_113 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0799_ _0799_/A _0799_/B vssd1 vssd1 vccd1 vccd1 _0913_/A sky130_fd_sc_hd__nand2_1
X_0868_ _0892_/A _0657_/X _0846_/A _0867_/Y vssd1 vssd1 vccd1 vccd1 _0868_/X sky130_fd_sc_hd__o2bb2a_1
XANTENNA__1067__B input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0937_ _0937_/A _0937_/B vssd1 vssd1 vccd1 vccd1 _0938_/B sky130_fd_sc_hd__nand2_1
XFILLER_43_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0651__B2 _0729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0651__A1 _1099_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0771__S _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0722_ _0757_/A vssd1 vssd1 vccd1 vccd1 _0724_/A sky130_fd_sc_hd__inv_2
X_0653_ _0653_/A _0653_/B _0653_/C vssd1 vssd1 vccd1 vccd1 _0925_/B sky130_fd_sc_hd__and3_1
XFILLER_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0584_ _0894_/A _0905_/A _1108_/A _1110_/A vssd1 vssd1 vccd1 vccd1 _0603_/B sky130_fd_sc_hd__or4_1
X_1136_ _1170_/C _1176_/A vssd1 vssd1 vccd1 vccd1 _1150_/A sky130_fd_sc_hd__xnor2_1
XFILLER_25_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1067_ _1086_/A input6/X vssd1 vssd1 vccd1 vccd1 _1067_/X sky130_fd_sc_hd__and2_1
XFILLER_40_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0633__A1 _0733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_109 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_271 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_16_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0927__A2 _0656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_0705_ _0738_/S _0703_/B _0791_/A vssd1 vssd1 vccd1 vccd1 _0705_/X sky130_fd_sc_hd__o21a_1
X_0636_ _0816_/B vssd1 vssd1 vccd1 vccd1 _0848_/B sky130_fd_sc_hd__buf_2
XANTENNA__0854__A1 _0843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1119_ _1119_/A _1119_/B _1119_/C vssd1 vssd1 vccd1 vccd1 _1119_/X sky130_fd_sc_hd__and3_1
XFILLER_21_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0790__B1 _1003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_171 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0836__A1 _0843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0619_ _0771_/S vssd1 vssd1 vccd1 vccd1 _0763_/A sky130_fd_sc_hd__inv_2
XFILLER_45_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_204 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0970_ _0969_/X _0954_/Y _0955_/A vssd1 vssd1 vccd1 vccd1 _0971_/A sky130_fd_sc_hd__a21o_1
XANTENNA__1176__A _1176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0809__A1 _0815_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0809__B2 _0808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1086__A _1086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1025__S _1099_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_152 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0774__S _0779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output39_A _1164_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0884_ _0884_/A _0884_/B vssd1 vssd1 vccd1 vccd1 _0884_/Y sky130_fd_sc_hd__nand2_1
X_0953_ _0954_/A _0954_/B _0954_/C vssd1 vssd1 vccd1 vccd1 _0955_/A sky130_fd_sc_hd__a21oi_1
XFILLER_23_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_99 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput16 i_l[8] vssd1 vssd1 vccd1 vccd1 _0952_/A sky130_fd_sc_hd__clkbuf_4
Xinput27 i_r[14] vssd1 vssd1 vccd1 vccd1 _1108_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_14_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0769__S _0781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1152_ _1152_/A _1152_/B _1152_/C _1152_/D vssd1 vssd1 vccd1 vccd1 _1152_/X sky130_fd_sc_hd__or4_1
X_1083_ _1057_/A _1057_/B _1067_/X _1055_/B vssd1 vssd1 vccd1 vccd1 _1083_/X sky130_fd_sc_hd__o31a_1
X_0936_ _0936_/A _0907_/C vssd1 vssd1 vccd1 vccd1 _0937_/B sky130_fd_sc_hd__or2b_1
X_0798_ _0805_/A _0798_/B vssd1 vssd1 vccd1 vccd1 _0799_/B sky130_fd_sc_hd__nand2_1
X_0867_ _0808_/A _0876_/A _0865_/X _0866_/X vssd1 vssd1 vccd1 vccd1 _0867_/Y sky130_fd_sc_hd__a211oi_1
XANTENNA__0651__A2 _0834_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0721_ _0771_/S _0763_/B vssd1 vssd1 vccd1 vccd1 _0757_/A sky130_fd_sc_hd__or2_1
X_0652_ _0866_/A _0651_/X _0711_/A vssd1 vssd1 vccd1 vccd1 _0652_/Y sky130_fd_sc_hd__o21ai_1
X_0583_ _1015_/A _1059_/A _1039_/A _1086_/A vssd1 vssd1 vccd1 vccd1 _0603_/A sky130_fd_sc_hd__or4_2
XFILLER_10_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1135_ _0770_/C _0656_/B _1174_/B vssd1 vssd1 vccd1 vccd1 _1176_/A sky130_fd_sc_hd__a21boi_4
X_1066_ _1086_/A _0834_/X _0808_/X _1055_/A _0866_/X vssd1 vssd1 vccd1 vccd1 _1066_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_33_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0919_ _0919_/A vssd1 vssd1 vccd1 vccd1 _1101_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_17_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1170__C _1170_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0704_ _0720_/A _0747_/A _0720_/C vssd1 vssd1 vccd1 vccd1 _0791_/A sky130_fd_sc_hd__and3_1
X_0635_ _0684_/A _0635_/B vssd1 vssd1 vccd1 vccd1 _0635_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__1040__A2 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0854__A2 _0848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1118_ _1118_/A _1118_/B _1173_/B vssd1 vssd1 vccd1 vccd1 _1119_/C sky130_fd_sc_hd__or3_1
X_1049_ input5/X _0656_/B _1119_/A _1034_/X _1048_/X vssd1 vssd1 vccd1 vccd1 _1049_/X
+ sky130_fd_sc_hd__a221o_1
XANTENNA__0721__A _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_220 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0836__A2 _0834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0618_ _0613_/Y _0617_/Y _0738_/S vssd1 vssd1 vccd1 vccd1 _0618_/X sky130_fd_sc_hd__mux2_1
XFILLER_41_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_88 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input20_A i_mode[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0809__A2 _0657_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_164 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_26_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_42 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_98 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0952_ _0952_/A vssd1 vssd1 vccd1 vccd1 _0954_/B sky130_fd_sc_hd__inv_2
X_0883_ _1004_/A _1003_/B _1102_/S vssd1 vssd1 vccd1 vccd1 _1125_/B sky130_fd_sc_hd__mux2_1
XFILLER_2_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput28 i_r[15] vssd1 vssd1 vccd1 vccd1 _1110_/A sky130_fd_sc_hd__buf_2
Xinput17 i_l[9] vssd1 vssd1 vccd1 vccd1 _0934_/B sky130_fd_sc_hd__clkbuf_1
XANTENNA_output51_A _1167_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1151_ _1151_/A _1151_/B vssd1 vssd1 vccd1 vccd1 _1152_/D sky130_fd_sc_hd__or2_1
XANTENNA__1134__A1 _1173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1082_ _1057_/A _1057_/B _1067_/X _1055_/B _1085_/B vssd1 vssd1 vccd1 vccd1 _1118_/B
+ sky130_fd_sc_hd__o311a_1
X_0866_ _0866_/A vssd1 vssd1 vccd1 vccd1 _0866_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_9_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0935_ _0935_/A _0935_/B vssd1 vssd1 vccd1 vccd1 _0954_/C sky130_fd_sc_hd__nand2_1
X_0797_ _0805_/A _0798_/B vssd1 vssd1 vccd1 vccd1 _0799_/A sky130_fd_sc_hd__or2_1
XFILLER_28_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_115 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0720_ _0720_/A _0747_/A _0720_/C vssd1 vssd1 vccd1 vccd1 _0824_/A sky130_fd_sc_hd__nand3_4
XFILLER_42_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0651_ _1099_/S _0834_/A _0646_/X _0729_/A _0650_/X vssd1 vssd1 vccd1 vccd1 _0651_/X
+ sky130_fd_sc_hd__a221o_1
XFILLER_40_5 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0582_ _0695_/A vssd1 vssd1 vccd1 vccd1 _0878_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_10_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1134_ _1173_/A _1115_/Y _1116_/X _1119_/X _1133_/X vssd1 vssd1 vccd1 vccd1 _1174_/B
+ sky130_fd_sc_hd__a311o_1
XFILLER_33_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1065_ _1173_/A _1091_/A _1091_/B vssd1 vssd1 vccd1 vccd1 _1077_/B sky130_fd_sc_hd__and3_1
XFILLER_18_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0849_ _0910_/A _0849_/B vssd1 vssd1 vccd1 vccd1 _0912_/A sky130_fd_sc_hd__nand2_1
X_0918_ _0878_/X _0917_/X _1073_/A vssd1 vssd1 vccd1 vccd1 _0918_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1170__D _1176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0703_ _0738_/S _0703_/B vssd1 vssd1 vccd1 vccd1 _0703_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__1025__A0 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0634_ _0892_/A _0874_/B _0779_/S vssd1 vssd1 vccd1 vccd1 _0635_/B sky130_fd_sc_hd__mux2_1
X_1117_ _1118_/A _1118_/B _1173_/B vssd1 vssd1 vccd1 vccd1 _1119_/B sky130_fd_sc_hd__o21ai_1
X_1048_ _1132_/A _1048_/B _1047_/X vssd1 vssd1 vccd1 vccd1 _1048_/X sky130_fd_sc_hd__or3b_1
XANTENNA__0721__B _0763_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0631__B _0631_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0617_ _0684_/A _0617_/B vssd1 vssd1 vccd1 vccd1 _0617_/Y sky130_fd_sc_hd__nand2_1
XANTENNA_input13_A i_l[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0642__A _0693_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0817__A _0843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0690__A1 _1155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input5_A i_l[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_33 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_1_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0882_ _0882_/A vssd1 vssd1 vccd1 vccd1 _1102_/S sky130_fd_sc_hd__clkbuf_4
XANTENNA__0672__A1 _0733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0951_ _0935_/B _0947_/X _0949_/X _0950_/Y vssd1 vssd1 vccd1 vccd1 _0951_/X sky130_fd_sc_hd__a211o_1
XFILLER_23_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0718__A2 _1103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_32 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput18 i_mode[0] vssd1 vssd1 vccd1 vccd1 _0595_/D sky130_fd_sc_hd__clkbuf_2
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput29 i_r[1] vssd1 vssd1 vccd1 vccd1 _0770_/A sky130_fd_sc_hd__buf_2
XANTENNA_output44_A _1166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1150_ _1150_/A _1150_/B vssd1 vssd1 vccd1 vccd1 _1150_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_28_7 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_45_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0893__A1 _0894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1081_ _1081_/A _1118_/A vssd1 vssd1 vccd1 vccd1 _1085_/B sky130_fd_sc_hd__nor2_1
XANTENNA__0830__A _1103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0865_ _0894_/A _0834_/A _0729_/A _0846_/B vssd1 vssd1 vccd1 vccd1 _0865_/X sky130_fd_sc_hd__a22o_1
X_0934_ _0975_/A _0934_/B vssd1 vssd1 vccd1 vccd1 _0935_/B sky130_fd_sc_hd__or2_1
X_0796_ _0886_/A _0796_/B vssd1 vssd1 vccd1 vccd1 _0798_/B sky130_fd_sc_hd__or2_1
XFILLER_51_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0650_ _0646_/X _0808_/A vssd1 vssd1 vccd1 vccd1 _0650_/X sky130_fd_sc_hd__and2b_1
X_0581_ _0581_/A vssd1 vssd1 vccd1 vccd1 _0695_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1064_ _1064_/A _1064_/B _1152_/C vssd1 vssd1 vccd1 vccd1 _1091_/B sky130_fd_sc_hd__or3b_1
X_1133_ _1133_/A _1133_/B _1133_/C vssd1 vssd1 vccd1 vccd1 _1133_/X sky130_fd_sc_hd__or3_1
XFILLER_19_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0779_ _0796_/B _0763_/B _0779_/S vssd1 vssd1 vccd1 vccd1 _0779_/X sky130_fd_sc_hd__mux2_1
X_0848_ _0848_/A _0848_/B _0846_/X vssd1 vssd1 vccd1 vccd1 _0849_/B sky130_fd_sc_hd__or3b_1
X_0917_ _0952_/A _0925_/A _1099_/S vssd1 vssd1 vccd1 vccd1 _0917_/X sky130_fd_sc_hd__mux2_1
XFILLER_24_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_23 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0702_ input9/X _0725_/B vssd1 vssd1 vccd1 vccd1 _0703_/B sky130_fd_sc_hd__xor2_2
X_0633_ _0733_/A _0629_/X _0632_/X vssd1 vssd1 vccd1 vccd1 _0633_/X sky130_fd_sc_hd__a21o_1
XANTENNA__1025__A1 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1116_ _1115_/A _1115_/B _1151_/B vssd1 vssd1 vccd1 vccd1 _1116_/X sky130_fd_sc_hd__a21o_1
XFILLER_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1047_ _1097_/A _0611_/X _1097_/B _0824_/A _1064_/B vssd1 vssd1 vccd1 vccd1 _1047_/X
+ sky130_fd_sc_hd__o32a_1
XFILLER_5_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_8_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0616_ _0952_/A _0975_/B _0779_/S vssd1 vssd1 vccd1 vccd1 _0617_/B sky130_fd_sc_hd__mux2_1
XFILLER_7_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_174 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0907__B _0925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0987__B1 _1132_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0690__A2 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0817__B _0848_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0978__A0 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_12 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_169 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0881_ _0826_/Y _0880_/Y _0919_/A vssd1 vssd1 vccd1 vccd1 _1003_/B sky130_fd_sc_hd__mux2_1
X_0950_ _1097_/B _0950_/B vssd1 vssd1 vccd1 vccd1 _0950_/Y sky130_fd_sc_hd__nor2_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0718__A3 _1003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0887__C1 _0866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0654__A2 _0595_/D vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_44 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_14_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput19 i_mode[1] vssd1 vssd1 vccd1 vccd1 _0595_/C sky130_fd_sc_hd__clkbuf_2
X_1080_ _1108_/A input7/X vssd1 vssd1 vccd1 vccd1 _1118_/A sky130_fd_sc_hd__and2_1
XFILLER_20_128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0830__B _0830_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0795_ _0811_/A _0831_/A vssd1 vssd1 vccd1 vccd1 _0805_/A sky130_fd_sc_hd__nor2_2
X_0864_ _0894_/A _0892_/A vssd1 vssd1 vccd1 vccd1 _0876_/A sky130_fd_sc_hd__nand2_1
XFILLER_9_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0933_ _0975_/A _0934_/B vssd1 vssd1 vccd1 vccd1 _0935_/A sky130_fd_sc_hd__nand2_2
XFILLER_3_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_231 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0650__B _0808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0580_ _0653_/A _0653_/B _0595_/C _0595_/D vssd1 vssd1 vccd1 vccd1 _0581_/A sky130_fd_sc_hd__and4b_1
X_1063_ _1064_/A _1064_/B _1152_/C vssd1 vssd1 vccd1 vccd1 _1091_/A sky130_fd_sc_hd__o21bai_1
X_1132_ _1132_/A _1132_/B _1132_/C _1131_/X vssd1 vssd1 vccd1 vccd1 _1133_/C sky130_fd_sc_hd__or4b_1
XFILLER_18_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0916_ _1173_/A _0957_/B _0957_/C vssd1 vssd1 vccd1 vccd1 _0916_/X sky130_fd_sc_hd__and3_1
X_0778_ _1006_/B _0778_/B _0778_/C vssd1 vssd1 vccd1 vccd1 _0784_/B sky130_fd_sc_hd__and3b_1
X_0847_ _0848_/A _0848_/B _0846_/X vssd1 vssd1 vccd1 vccd1 _0910_/A sky130_fd_sc_hd__o21bai_1
XFILLER_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input36_A i_r[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0661__A _1099_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_256 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0701_ _0693_/B _0661_/B _0700_/X vssd1 vssd1 vccd1 vccd1 _0725_/B sky130_fd_sc_hd__o21ai_2
X_0632_ _1155_/A input9/X _0711_/A _0781_/A vssd1 vssd1 vccd1 vccd1 _0632_/X sky130_fd_sc_hd__o211a_1
XFILLER_38_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1115_ _1115_/A _1115_/B _1151_/B vssd1 vssd1 vccd1 vccd1 _1115_/Y sky130_fd_sc_hd__nand3_1
X_1046_ _1152_/A _1152_/B vssd1 vssd1 vccd1 vccd1 _1064_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__0775__A1 _0779_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1016__A2 input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0615_ _0934_/B vssd1 vssd1 vccd1 vccd1 _0975_/B sky130_fd_sc_hd__clkbuf_4
X_1029_ _1124_/A _1029_/B vssd1 vssd1 vccd1 vccd1 _1029_/Y sky130_fd_sc_hd__nand2_1
XFILLER_30_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0987__A1 _1015_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1164__A1 _1173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0978__A1 _0975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_25_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_49_248 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_244 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_32_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0934__A _0975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0880_ _0878_/X _0879_/X _1073_/A vssd1 vssd1 vccd1 vccd1 _0880_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__0844__A _0894_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_26 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_11_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0887__B1 _0808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0932_ _0932_/A vssd1 vssd1 vccd1 vccd1 _1169_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_9_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0794_ _0815_/A _1131_/A vssd1 vssd1 vccd1 vccd1 _0831_/A sky130_fd_sc_hd__and2_1
X_0863_ _1097_/A _0734_/X _0738_/X _0884_/A vssd1 vssd1 vccd1 vccd1 _0863_/X sky130_fd_sc_hd__a22o_1
XFILLER_3_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1037__B1 _0808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1131_ _1131_/A _1131_/B _1131_/C _1131_/D vssd1 vssd1 vccd1 vccd1 _1131_/X sky130_fd_sc_hd__or4_1
X_1062_ _1062_/A _1061_/X vssd1 vssd1 vccd1 vccd1 _1152_/C sky130_fd_sc_hd__or2b_1
XFILLER_18_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0915_ _0914_/B _0914_/C _0914_/A vssd1 vssd1 vccd1 vccd1 _0957_/C sky130_fd_sc_hd__a21o_1
X_0777_ _0627_/X _0773_/X _0884_/B _1097_/A _1006_/A vssd1 vssd1 vccd1 vccd1 _0778_/C
+ sky130_fd_sc_hd__a221o_1
X_0846_ _0846_/A _0846_/B vssd1 vssd1 vccd1 vccd1 _0846_/X sky130_fd_sc_hd__or2_1
XFILLER_24_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1019__B1 _0824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input29_A i_r[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1103__A _1103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0700_ input1/X input2/X vssd1 vssd1 vccd1 vccd1 _0700_/X sky130_fd_sc_hd__or2b_1
XFILLER_30_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0631_ input2/X _0631_/B vssd1 vssd1 vccd1 vccd1 _0711_/A sky130_fd_sc_hd__or2_1
XFILLER_24_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1114_ _1114_/A _1114_/B vssd1 vssd1 vccd1 vccd1 _1151_/B sky130_fd_sc_hd__nand2_1
XFILLER_0_61 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1045_ _0957_/C _1042_/X _1043_/X _1044_/Y vssd1 vssd1 vccd1 vccd1 _1152_/B sky130_fd_sc_hd__o211a_1
XANTENNA__0775__A2 _0975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0829_ _0692_/X _0939_/B _0882_/A vssd1 vssd1 vccd1 vccd1 _0830_/B sky130_fd_sc_hd__mux2_2
XFILLER_9_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_268 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_5_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0656__B _0656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_7_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_290 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0614_ _0669_/A vssd1 vssd1 vccd1 vccd1 _0684_/A sky130_fd_sc_hd__buf_2
XANTENNA__0611__S _0738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0582__A _0695_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1028_ _0920_/X _1027_/X _1102_/S vssd1 vssd1 vccd1 vccd1 _1029_/B sky130_fd_sc_hd__mux2_1
XFILLER_39_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_44_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0987__A2 _0834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0667__A _1155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0969__A2 _0925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_256 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input11_A i_l[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0844__B _0892_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0887__A1 _0905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input3_A i_l[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_149 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_37_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0862_ _1097_/A _1097_/C _1006_/A vssd1 vssd1 vccd1 vccd1 _0862_/X sky130_fd_sc_hd__o21a_1
X_0931_ _1119_/A _0904_/Y _0916_/X _0930_/Y vssd1 vssd1 vccd1 vccd1 _0932_/A sky130_fd_sc_hd__a211o_1
XFILLER_9_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0793_ _0815_/A _1131_/A vssd1 vssd1 vccd1 vccd1 _0811_/A sky130_fd_sc_hd__nor2_1
XFILLER_9_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1037__A1 _1059_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_output42_A _1150_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1130_ _1130_/A _1155_/B vssd1 vssd1 vccd1 vccd1 _1132_/C sky130_fd_sc_hd__nor2_1
XFILLER_33_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1061_ _1061_/A input5/X _1061_/C vssd1 vssd1 vccd1 vccd1 _1061_/X sky130_fd_sc_hd__or3_1
XANTENNA__0675__A _1155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0845_ _0894_/A _0892_/A vssd1 vssd1 vccd1 vccd1 _0846_/B sky130_fd_sc_hd__and2_1
X_0914_ _0914_/A _0914_/B _0914_/C vssd1 vssd1 vccd1 vccd1 _0957_/B sky130_fd_sc_hd__nand3_1
X_0776_ _0781_/A _0684_/A _0774_/X _0775_/X vssd1 vssd1 vccd1 vccd1 _0884_/B sky130_fd_sc_hd__a31o_1
XFILLER_24_211 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0585__A _0954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0630_ _0693_/B vssd1 vssd1 vccd1 vccd1 _1155_/A sky130_fd_sc_hd__clkinv_2
X_1113_ _1113_/A input7/X _1173_/B vssd1 vssd1 vccd1 vccd1 _1114_/B sky130_fd_sc_hd__or3_1
X_1044_ _1014_/A _1018_/B _1018_/A vssd1 vssd1 vccd1 vccd1 _1044_/Y sky130_fd_sc_hd__a21boi_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_225 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0759_ _0759_/A _0796_/B vssd1 vssd1 vccd1 vccd1 _0759_/X sky130_fd_sc_hd__and2_1
X_0828_ _1007_/A _0828_/B vssd1 vssd1 vccd1 vccd1 _0882_/A sky130_fd_sc_hd__xnor2_2
XFILLER_9_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0613_ _0669_/A _0613_/B vssd1 vssd1 vccd1 vccd1 _0613_/Y sky130_fd_sc_hd__nand2_1
XFILLER_38_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1027_ _0979_/Y _1026_/Y _1101_/S vssd1 vssd1 vccd1 vccd1 _1027_/X sky130_fd_sc_hd__mux2_1
XFILLER_30_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_188 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1094__C1 _0866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1109__A _1110_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0948__A _0975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_128 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_6_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0593__A _0595_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_268 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_147 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0588__A input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0887__A2 _0834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0945__B _1003_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0792_ _0766_/S _0764_/B _0764_/A vssd1 vssd1 vccd1 vccd1 _0800_/A sky130_fd_sc_hd__a21o_1
X_0861_ _0744_/X _0860_/X _0882_/A vssd1 vssd1 vccd1 vccd1 _0861_/X sky130_fd_sc_hd__mux2_1
X_0930_ _0621_/X _1097_/B _1103_/A _0921_/X _0929_/X vssd1 vssd1 vccd1 vccd1 _0930_/Y
+ sky130_fd_sc_hd__o221ai_2
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_47_57 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0781__A _0781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1037__A2 _0834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1060_ _1061_/A input5/X _1061_/C vssd1 vssd1 vccd1 vccd1 _1062_/A sky130_fd_sc_hd__o21a_1
XANTENNA__0675__B input3/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_220 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_33_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0913_ _0913_/A _0913_/B _0913_/C _0800_/A vssd1 vssd1 vccd1 vccd1 _0914_/C sky130_fd_sc_hd__or4b_1
X_0775_ _0779_/S _0975_/B _0669_/A _0675_/X _0770_/A vssd1 vssd1 vccd1 vccd1 _0775_/X
+ sky130_fd_sc_hd__o2111a_1
X_0844_ _0894_/A _0892_/A vssd1 vssd1 vccd1 vccd1 _0846_/A sky130_fd_sc_hd__nor2_1
XANTENNA__0866__A _0866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0585__B _0975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_226 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_30_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1112_ _1113_/A input7/X _1173_/B vssd1 vssd1 vccd1 vccd1 _1114_/A sky130_fd_sc_hd__o21ai_1
XFILLER_0_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1043_ _1043_/A _1043_/B _1043_/C vssd1 vssd1 vccd1 vccd1 _1043_/X sky130_fd_sc_hd__or3_1
XFILLER_21_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0758_ _0764_/A _0758_/B vssd1 vssd1 vccd1 vccd1 _0758_/Y sky130_fd_sc_hd__xnor2_1
X_0827_ _0780_/Y _0826_/Y _0919_/A vssd1 vssd1 vccd1 vccd1 _0939_/B sky130_fd_sc_hd__mux2_1
X_0689_ _0733_/A _0781_/B vssd1 vssd1 vccd1 vccd1 _1155_/C sky130_fd_sc_hd__xnor2_2
XFILLER_29_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0999__A1 _1099_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input34_A i_r[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_90 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_7_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0612_ input3/X input4/X _0693_/B vssd1 vssd1 vccd1 vccd1 _0613_/B sky130_fd_sc_hd__mux2_1
XFILLER_38_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1026_ _0878_/X _1025_/X _1073_/A vssd1 vssd1 vccd1 vccd1 _1026_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__1024__B _1024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_16 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_39_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1094__B1 _0808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1109__B input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0948__B _0975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0832__B1 _0748_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__0874__A _0905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1009_ _1039_/A _0834_/X _0808_/X _1017_/C vssd1 vssd1 vccd1 vccd1 _1009_/X sky130_fd_sc_hd__a22o_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0587__C1 _0975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_151 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_262 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_48_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0694__A _0771_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_184 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1049__B1 _1119_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0791_ _0791_/A vssd1 vssd1 vccd1 vccd1 _1173_/A sky130_fd_sc_hd__buf_4
X_0860_ _0788_/Y _0859_/Y _0919_/A vssd1 vssd1 vccd1 vccd1 _0860_/X sky130_fd_sc_hd__mux2_1
XFILLER_13_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0689__A _0733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0989_ _1119_/A _0977_/Y _0988_/X vssd1 vssd1 vccd1 vccd1 _0989_/X sky130_fd_sc_hd__a21o_1
XFILLER_47_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_27_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_232 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0912_ _0912_/A _0912_/B vssd1 vssd1 vccd1 vccd1 _0913_/C sky130_fd_sc_hd__or2_1
XFILLER_33_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_0774_ _0874_/B _0952_/A _0779_/S vssd1 vssd1 vccd1 vccd1 _0774_/X sky130_fd_sc_hd__mux2_1
X_0843_ _0843_/A vssd1 vssd1 vccd1 vccd1 _0848_/A sky130_fd_sc_hd__inv_2
XFILLER_30_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1099__S _1099_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1042_ _1042_/A _1043_/A _1043_/C vssd1 vssd1 vccd1 vccd1 _1042_/X sky130_fd_sc_hd__or3_1
X_1111_ _1111_/A _1128_/A vssd1 vssd1 vccd1 vccd1 _1173_/B sky130_fd_sc_hd__and2_1
XFILLER_21_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0757_ _0757_/A _0757_/B vssd1 vssd1 vccd1 vccd1 _0758_/B sky130_fd_sc_hd__nand2_1
X_0688_ _0779_/S _0695_/A vssd1 vssd1 vccd1 vccd1 _0781_/B sky130_fd_sc_hd__nand2_2
X_0826_ _0878_/A _0825_/X _0787_/A vssd1 vssd1 vccd1 vccd1 _0826_/Y sky130_fd_sc_hd__o21ai_1
XANTENNA__1038__A input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0999__A2 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input27_A i_r[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0611_ _0733_/B _0608_/Y _0738_/S vssd1 vssd1 vccd1 vccd1 _0611_/X sky130_fd_sc_hd__mux2_1
XFILLER_7_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0773__S1 _0733_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1025_ input5/X input4/X _1099_/S vssd1 vssd1 vccd1 vccd1 _1025_/X sky130_fd_sc_hd__mux2_1
XFILLER_14_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_0809_ _0815_/A _0657_/X _0805_/A _0808_/X vssd1 vssd1 vccd1 vccd1 _0809_/Y sky130_fd_sc_hd__a22oi_1
XFILLER_39_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1094__A1 _1108_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_4_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0948__C _0948_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1141__A _1167_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_80 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_43_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__0874__B _0874_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1008_ _1097_/A _0769_/X _1007_/X vssd1 vssd1 vccd1 vccd1 _1008_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_25_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0587__B1 _0843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0814__A1 _1103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_163 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_40_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1136__A _1170_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_274 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_0_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0975__A _0975_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output58_A _1169_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_141 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_119 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_23_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1049__A1 input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0734__S _0781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0790_ _1007_/A _1007_/B _0600_/B _1003_/A _0789_/X vssd1 vssd1 vccd1 vccd1 _1024_/B
+ sky130_fd_sc_hd__o32a_2
XFILLER_9_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0988_ _0923_/A _0982_/Y _0983_/Y _0987_/X vssd1 vssd1 vccd1 vccd1 _0988_/X sky130_fd_sc_hd__a31o_1
XFILLER_22_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_15 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA_input1_A i_carry vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_255 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_10_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0842_ _0842_/A vssd1 vssd1 vccd1 vccd1 _1168_/B sky130_fd_sc_hd__clkbuf_1
XFILLER_33_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0911_ _0912_/A _0909_/Y _0912_/B _0910_/X _0895_/A vssd1 vssd1 vccd1 vccd1 _0914_/B
+ sky130_fd_sc_hd__o311a_1
X_0773_ _0796_/B _0815_/A _0848_/B _0892_/A _0858_/S _0733_/A vssd1 vssd1 vccd1 vccd1
+ _0773_/X sky130_fd_sc_hd__mux4_1
XFILLER_5_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0639__S _0738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0632__C1 _0781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0926__B1 _0808_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_output40_A _1176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1110_ _1110_/A input8/X vssd1 vssd1 vccd1 vccd1 _1128_/A sky130_fd_sc_hd__or2_1
X_1041_ _1039_/A _1038_/Y _1064_/A vssd1 vssd1 vccd1 vccd1 _1152_/A sky130_fd_sc_hd__a21o_1
X_0825_ _0848_/B _0815_/A _0858_/S vssd1 vssd1 vccd1 vccd1 _0825_/X sky130_fd_sc_hd__mux2_1
XFILLER_9_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0756_ _0711_/A _0711_/B _0711_/D _0724_/B _0745_/A vssd1 vssd1 vccd1 vccd1 _0757_/B
+ sky130_fd_sc_hd__a311o_1
X_0687_ _1006_/A _0950_/B _0686_/X _1006_/B vssd1 vssd1 vccd1 vccd1 _0719_/A sky130_fd_sc_hd__a211o_1
XANTENNA__0917__A0 _0952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1054__A _1086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0610_ _0781_/A vssd1 vssd1 vccd1 vccd1 _0738_/S sky130_fd_sc_hd__clkbuf_4
XFILLER_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0917__S _1099_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1024_ _1125_/A _1024_/B vssd1 vssd1 vccd1 vccd1 _1024_/Y sky130_fd_sc_hd__nand2_1
X_0808_ _0808_/A vssd1 vssd1 vccd1 vccd1 _0808_/X sky130_fd_sc_hd__clkbuf_4
XFILLER_30_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0888__A _0905_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0739_ _0736_/Y _0737_/X _0685_/Y _0738_/X vssd1 vssd1 vccd1 vccd1 _0739_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_29_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1094__A2 _0834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_279 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1141__B _1167_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1007_ _1007_/A _1007_/B _1131_/D vssd1 vssd1 vccd1 vccd1 _1007_/X sky130_fd_sc_hd__or3_1
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_19_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_227 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_1_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0587__A1 _1131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0814__A2 _1024_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_175 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_15_95 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1136__B _1176_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput50 _1167_/B vssd1 vssd1 vccd1 vccd1 o_out[1] sky130_fd_sc_hd__buf_2
XFILLER_48_286 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0975__B _0975_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0741__A1 _0824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1049__A2 _0656_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1147__A _1166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_21 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_259 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_36_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_0987_ _1015_/A _0834_/X _1132_/A _0984_/Y _0986_/X vssd1 vssd1 vccd1 vccd1 _0987_/X
+ sky130_fd_sc_hd__a2111o_1
XFILLER_47_27 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_267 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__0953__A1 _0954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0705__A1 _0738_/S vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0841_ _0841_/A _0841_/B _0841_/C _0841_/D vssd1 vssd1 vccd1 vccd1 _0842_/A sky130_fd_sc_hd__or4_1
XFILLER_41_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_0772_ _1006_/A _0772_/B vssd1 vssd1 vccd1 vccd1 _0778_/B sky130_fd_sc_hd__nand2_1
X_0910_ _0910_/A _0895_/B vssd1 vssd1 vccd1 vccd1 _0910_/X sky130_fd_sc_hd__or2b_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0623__B1 _1131_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0926__A1 _0954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1040_ _1039_/Y input4/X _1038_/B vssd1 vssd1 vccd1 vccd1 _1064_/A sky130_fd_sc_hd__o21a_1
X_0755_ _0755_/A vssd1 vssd1 vccd1 vccd1 _0764_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_0824_ _0824_/A _0824_/B vssd1 vssd1 vccd1 vccd1 _0841_/A sky130_fd_sc_hd__nor2_1
XANTENNA__0917__A1 _0925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0686_ _0884_/A _0681_/Y _0684_/Y _0685_/Y vssd1 vssd1 vccd1 vccd1 _0686_/X sky130_fd_sc_hd__a22o_1
XFILLER_28_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1054__B input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1169_ _1169_/A _1169_/B _1169_/C vssd1 vssd1 vccd1 vccd1 _1171_/C sky130_fd_sc_hd__or3_1
XFILLER_20_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1155__A _1155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0835__A0 _0729_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0994__A _1039_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1023_ _1023_/A vssd1 vssd1 vccd1 vccd1 _1166_/B sky130_fd_sc_hd__clkbuf_2
X_0807_ _0884_/A _0639_/X _0685_/Y _0618_/X vssd1 vssd1 vccd1 vccd1 _0807_/X sky130_fd_sc_hd__a22o_1
X_0738_ _0617_/Y _0635_/Y _0738_/S vssd1 vssd1 vccd1 vccd1 _0738_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0888__B _0925_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1065__A _1173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0669_ _0669_/A _0669_/B _0669_/C vssd1 vssd1 vccd1 vccd1 _0669_/Y sky130_fd_sc_hd__nand3_1
XFILLER_4_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_41 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_28_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input32_A i_r[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1006_ _1006_/A _1006_/B vssd1 vssd1 vccd1 vccd1 _1006_/Y sky130_fd_sc_hd__nor2_1
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__0899__A _0954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0602__A _0843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput51 _1167_/C vssd1 vssd1 vccd1 vccd1 o_out[2] sky130_fd_sc_hd__buf_2
Xoutput40 _1176_/A vssd1 vssd1 vccd1 vccd1 o_flags[2] sky130_fd_sc_hd__buf_2
XFILLER_48_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_121 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_42_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__0708__C1 _0866_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1147__B _1166_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_33 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_51_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_0986_ _0866_/X _0985_/X _0964_/A vssd1 vssd1 vccd1 vccd1 _0986_/X sky130_fd_sc_hd__o21ba_1
XANTENNA__0947__C1 _0866_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_39 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_27_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_3 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_2_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_0840_ _0848_/B _0657_/X _0855_/C _0836_/X _0839_/Y vssd1 vssd1 vccd1 vccd1 _0841_/D
+ sky130_fd_sc_hd__a221o_1
X_0771_ _0769_/X _0770_/X _0771_/S vssd1 vssd1 vccd1 vccd1 _0772_/B sky130_fd_sc_hd__mux2_1
XFILLER_5_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__0632__A1 _1155_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0969_ _0907_/A _0925_/A _0907_/C vssd1 vssd1 vccd1 vccd1 _0969_/X sky130_fd_sc_hd__o21a_1
XANTENNA__0700__A input1/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0871__A1 _1173_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0610__A _0781_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__0926__A2 _0834_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_0754_ _0754_/A _0754_/B vssd1 vssd1 vccd1 vccd1 _0755_/A sky130_fd_sc_hd__and2_1
X_0823_ _0913_/B _0823_/B vssd1 vssd1 vccd1 vccd1 _0824_/B sky130_fd_sc_hd__xnor2_1
X_0685_ _1006_/A _1007_/A vssd1 vssd1 vccd1 vccd1 _0685_/Y sky130_fd_sc_hd__nor2_1
XFILLER_28_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1168_ _1168_/A _1168_/B _1168_/C vssd1 vssd1 vccd1 vccd1 _1169_/C sky130_fd_sc_hd__or3_1
XFILLER_44_29 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
X_1099_ input7/X input6/X _1099_/S vssd1 vssd1 vccd1 vccd1 _1099_/X sky130_fd_sc_hd__mux2_1
XANTENNA__0605__A1 input8/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0994__B input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__0835__A1 _0808_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1088__A1 _1086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1022_ _0997_/Y _0998_/X _1013_/X _1021_/X vssd1 vssd1 vccd1 vccd1 _1023_/A sky130_fd_sc_hd__a211o_1
X_0806_ _1097_/A _0611_/X _1006_/A vssd1 vssd1 vccd1 vccd1 _0806_/X sky130_fd_sc_hd__o21a_1
X_0737_ _0738_/S _0684_/A _0629_/X _0771_/S _0759_/A vssd1 vssd1 vccd1 vccd1 _0737_/X
+ sky130_fd_sc_hd__a311o_1
XANTENNA__0888__C _0948_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_0668_ _0693_/B input6/X vssd1 vssd1 vccd1 vccd1 _0669_/C sky130_fd_sc_hd__or2_1
X_0599_ _0878_/A _1161_/A _1126_/A vssd1 vssd1 vccd1 vccd1 _0923_/A sky130_fd_sc_hd__o21a_2
XFILLER_37_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_53 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XFILLER_35_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input25_A i_r[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_281 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__1166__A _1166_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1005_ _1124_/A _1002_/Y _1003_/Y _1004_/Y _0945_/Y vssd1 vssd1 vccd1 vccd1 _1005_/X
+ sky130_fd_sc_hd__a32o_1
XFILLER_41_19 vssd1 vccd1 vccd1 vssd1 sky130_ef_sc_hd__decap_12
XANTENNA__0899__B _0952_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1076__A _1103_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput52 _1167_/D vssd1 vssd1 vccd1 vccd1 o_out[3] sky130_fd_sc_hd__buf_2
XFILLER_31_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput41 _1175_/X vssd1 vssd1 vccd1 vccd1 o_flags[3] sky130_fd_sc_hd__buf_2
XANTENNA__0602__B _0954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1160__B1 _0848_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

