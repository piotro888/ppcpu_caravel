VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO int_ram
  CLASS BLOCK ;
  FOREIGN int_ram ;
  ORIGIN 0.000 0.000 ;
  SIZE 800.000 BY 350.000 ;
  PIN i_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 36.960 800.000 37.520 ;
    END
  END i_addr[0]
  PIN i_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 60.480 800.000 61.040 ;
    END
  END i_addr[1]
  PIN i_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 84.000 800.000 84.560 ;
    END
  END i_addr[2]
  PIN i_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 107.520 800.000 108.080 ;
    END
  END i_addr[3]
  PIN i_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 131.040 800.000 131.600 ;
    END
  END i_addr[4]
  PIN i_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 154.560 800.000 155.120 ;
    END
  END i_addr[5]
  PIN i_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 21.280 800.000 21.840 ;
    END
  END i_clk
  PIN i_data[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 44.800 800.000 45.360 ;
    END
  END i_data[0]
  PIN i_data[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 240.800 800.000 241.360 ;
    END
  END i_data[10]
  PIN i_data[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 256.480 800.000 257.040 ;
    END
  END i_data[11]
  PIN i_data[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 272.160 800.000 272.720 ;
    END
  END i_data[12]
  PIN i_data[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 287.840 800.000 288.400 ;
    END
  END i_data[13]
  PIN i_data[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 303.520 800.000 304.080 ;
    END
  END i_data[14]
  PIN i_data[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 319.200 800.000 319.760 ;
    END
  END i_data[15]
  PIN i_data[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 68.320 800.000 68.880 ;
    END
  END i_data[1]
  PIN i_data[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 91.840 800.000 92.400 ;
    END
  END i_data[2]
  PIN i_data[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 115.360 800.000 115.920 ;
    END
  END i_data[3]
  PIN i_data[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 138.880 800.000 139.440 ;
    END
  END i_data[4]
  PIN i_data[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 162.400 800.000 162.960 ;
    END
  END i_data[5]
  PIN i_data[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 178.080 800.000 178.640 ;
    END
  END i_data[6]
  PIN i_data[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 193.760 800.000 194.320 ;
    END
  END i_data[7]
  PIN i_data[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 209.440 800.000 210.000 ;
    END
  END i_data[8]
  PIN i_data[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 225.120 800.000 225.680 ;
    END
  END i_data[9]
  PIN i_we
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 29.120 800.000 29.680 ;
    END
  END i_we
  PIN o_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 52.640 800.000 53.200 ;
    END
  END o_data[0]
  PIN o_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 248.640 800.000 249.200 ;
    END
  END o_data[10]
  PIN o_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 264.320 800.000 264.880 ;
    END
  END o_data[11]
  PIN o_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 280.000 800.000 280.560 ;
    END
  END o_data[12]
  PIN o_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 295.680 800.000 296.240 ;
    END
  END o_data[13]
  PIN o_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 311.360 800.000 311.920 ;
    END
  END o_data[14]
  PIN o_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 327.040 800.000 327.600 ;
    END
  END o_data[15]
  PIN o_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 76.160 800.000 76.720 ;
    END
  END o_data[1]
  PIN o_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 99.680 800.000 100.240 ;
    END
  END o_data[2]
  PIN o_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 123.200 800.000 123.760 ;
    END
  END o_data[3]
  PIN o_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 146.720 800.000 147.280 ;
    END
  END o_data[4]
  PIN o_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 170.240 800.000 170.800 ;
    END
  END o_data[5]
  PIN o_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 185.920 800.000 186.480 ;
    END
  END o_data[6]
  PIN o_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 201.600 800.000 202.160 ;
    END
  END o_data[7]
  PIN o_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 217.280 800.000 217.840 ;
    END
  END o_data[8]
  PIN o_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.080400 ;
    PORT
      LAYER Metal3 ;
        RECT 796.000 232.960 800.000 233.520 ;
    END
  END o_data[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 333.500 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 333.500 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 333.500 ;
    END
  END vssd1
  OBS
      LAYER Nwell ;
        RECT 6.290 331.165 793.390 333.630 ;
        RECT 6.290 331.040 151.240 331.165 ;
      LAYER Pwell ;
        RECT 6.290 327.520 793.390 331.040 ;
      LAYER Nwell ;
        RECT 6.290 327.395 73.745 327.520 ;
        RECT 6.290 323.325 793.390 327.395 ;
        RECT 6.290 323.200 73.185 323.325 ;
      LAYER Pwell ;
        RECT 6.290 319.680 793.390 323.200 ;
      LAYER Nwell ;
        RECT 6.290 319.555 95.025 319.680 ;
        RECT 6.290 315.485 793.390 319.555 ;
        RECT 6.290 315.360 51.905 315.485 ;
      LAYER Pwell ;
        RECT 6.290 311.840 793.390 315.360 ;
      LAYER Nwell ;
        RECT 6.290 311.715 71.505 311.840 ;
        RECT 6.290 307.645 793.390 311.715 ;
        RECT 6.290 307.520 124.145 307.645 ;
      LAYER Pwell ;
        RECT 6.290 304.000 793.390 307.520 ;
      LAYER Nwell ;
        RECT 6.290 303.875 51.905 304.000 ;
        RECT 6.290 299.805 793.390 303.875 ;
        RECT 6.290 299.680 49.105 299.805 ;
      LAYER Pwell ;
        RECT 6.290 296.160 793.390 299.680 ;
      LAYER Nwell ;
        RECT 6.290 296.035 68.145 296.160 ;
        RECT 6.290 291.965 793.390 296.035 ;
        RECT 6.290 291.840 127.160 291.965 ;
      LAYER Pwell ;
        RECT 6.290 288.320 793.390 291.840 ;
      LAYER Nwell ;
        RECT 6.290 288.195 51.905 288.320 ;
        RECT 6.290 284.125 793.390 288.195 ;
        RECT 6.290 284.000 47.985 284.125 ;
      LAYER Pwell ;
        RECT 6.290 280.480 793.390 284.000 ;
      LAYER Nwell ;
        RECT 6.290 280.355 149.905 280.480 ;
        RECT 6.290 276.285 793.390 280.355 ;
        RECT 6.290 276.160 52.465 276.285 ;
      LAYER Pwell ;
        RECT 6.290 272.640 793.390 276.160 ;
      LAYER Nwell ;
        RECT 6.290 272.515 93.345 272.640 ;
        RECT 6.290 268.445 793.390 272.515 ;
        RECT 6.290 268.320 35.105 268.445 ;
      LAYER Pwell ;
        RECT 6.290 264.800 793.390 268.320 ;
      LAYER Nwell ;
        RECT 6.290 264.675 34.545 264.800 ;
        RECT 6.290 260.605 793.390 264.675 ;
        RECT 6.290 260.480 39.025 260.605 ;
      LAYER Pwell ;
        RECT 6.290 256.960 793.390 260.480 ;
      LAYER Nwell ;
        RECT 6.290 256.835 65.905 256.960 ;
        RECT 6.290 252.765 793.390 256.835 ;
        RECT 6.290 252.640 32.305 252.765 ;
      LAYER Pwell ;
        RECT 6.290 249.120 793.390 252.640 ;
      LAYER Nwell ;
        RECT 6.290 248.995 93.345 249.120 ;
        RECT 6.290 244.925 793.390 248.995 ;
        RECT 6.290 244.800 41.825 244.925 ;
      LAYER Pwell ;
        RECT 6.290 241.280 793.390 244.800 ;
      LAYER Nwell ;
        RECT 6.290 241.155 31.745 241.280 ;
        RECT 6.290 237.085 793.390 241.155 ;
        RECT 6.290 236.960 46.305 237.085 ;
      LAYER Pwell ;
        RECT 6.290 233.440 793.390 236.960 ;
      LAYER Nwell ;
        RECT 6.290 233.315 98.385 233.440 ;
        RECT 6.290 229.245 793.390 233.315 ;
        RECT 6.290 229.120 14.945 229.245 ;
      LAYER Pwell ;
        RECT 6.290 225.600 793.390 229.120 ;
      LAYER Nwell ;
        RECT 6.290 225.475 51.905 225.600 ;
        RECT 6.290 221.405 793.390 225.475 ;
        RECT 6.290 221.280 47.425 221.405 ;
      LAYER Pwell ;
        RECT 6.290 217.760 793.390 221.280 ;
      LAYER Nwell ;
        RECT 6.290 217.635 17.745 217.760 ;
        RECT 6.290 213.565 793.390 217.635 ;
        RECT 6.290 213.440 14.945 213.565 ;
      LAYER Pwell ;
        RECT 6.290 209.920 793.390 213.440 ;
      LAYER Nwell ;
        RECT 6.290 209.795 110.145 209.920 ;
        RECT 6.290 205.725 793.390 209.795 ;
        RECT 6.290 205.600 71.505 205.725 ;
      LAYER Pwell ;
        RECT 6.290 202.080 793.390 205.600 ;
      LAYER Nwell ;
        RECT 6.290 201.955 16.065 202.080 ;
        RECT 6.290 197.885 793.390 201.955 ;
        RECT 6.290 197.760 14.945 197.885 ;
      LAYER Pwell ;
        RECT 6.290 194.240 793.390 197.760 ;
      LAYER Nwell ;
        RECT 6.290 194.115 70.600 194.240 ;
        RECT 6.290 190.045 793.390 194.115 ;
        RECT 6.290 189.920 14.945 190.045 ;
      LAYER Pwell ;
        RECT 6.290 186.400 793.390 189.920 ;
      LAYER Nwell ;
        RECT 6.290 186.275 97.825 186.400 ;
        RECT 6.290 182.205 793.390 186.275 ;
        RECT 6.290 182.080 43.505 182.205 ;
      LAYER Pwell ;
        RECT 6.290 178.560 793.390 182.080 ;
      LAYER Nwell ;
        RECT 6.290 178.435 23.345 178.560 ;
        RECT 6.290 174.365 793.390 178.435 ;
        RECT 6.290 174.240 14.945 174.365 ;
      LAYER Pwell ;
        RECT 6.290 170.720 793.390 174.240 ;
      LAYER Nwell ;
        RECT 6.290 170.595 22.225 170.720 ;
        RECT 6.290 166.525 793.390 170.595 ;
        RECT 6.290 166.400 32.305 166.525 ;
      LAYER Pwell ;
        RECT 6.290 162.880 793.390 166.400 ;
      LAYER Nwell ;
        RECT 6.290 162.755 102.865 162.880 ;
        RECT 6.290 158.685 793.390 162.755 ;
        RECT 6.290 158.560 163.345 158.685 ;
      LAYER Pwell ;
        RECT 6.290 155.040 793.390 158.560 ;
      LAYER Nwell ;
        RECT 6.290 154.915 20.545 155.040 ;
        RECT 6.290 150.845 793.390 154.915 ;
        RECT 6.290 150.720 37.905 150.845 ;
      LAYER Pwell ;
        RECT 6.290 147.200 793.390 150.720 ;
      LAYER Nwell ;
        RECT 6.290 147.075 29.505 147.200 ;
        RECT 6.290 143.005 793.390 147.075 ;
        RECT 6.290 142.880 40.705 143.005 ;
      LAYER Pwell ;
        RECT 6.290 139.360 793.390 142.880 ;
      LAYER Nwell ;
        RECT 6.290 139.235 63.665 139.360 ;
        RECT 6.290 135.165 793.390 139.235 ;
        RECT 6.290 135.040 132.545 135.165 ;
      LAYER Pwell ;
        RECT 6.290 131.520 793.390 135.040 ;
      LAYER Nwell ;
        RECT 6.290 131.395 69.825 131.520 ;
        RECT 6.290 127.325 793.390 131.395 ;
        RECT 6.290 127.200 42.945 127.325 ;
      LAYER Pwell ;
        RECT 6.290 123.680 793.390 127.200 ;
      LAYER Nwell ;
        RECT 6.290 123.555 56.385 123.680 ;
        RECT 6.290 119.485 793.390 123.555 ;
        RECT 6.290 119.360 33.985 119.485 ;
      LAYER Pwell ;
        RECT 6.290 115.840 793.390 119.360 ;
      LAYER Nwell ;
        RECT 6.290 115.715 96.705 115.840 ;
        RECT 6.290 111.645 793.390 115.715 ;
        RECT 6.290 111.520 51.905 111.645 ;
      LAYER Pwell ;
        RECT 6.290 108.000 793.390 111.520 ;
      LAYER Nwell ;
        RECT 6.290 107.875 34.545 108.000 ;
        RECT 6.290 103.805 793.390 107.875 ;
        RECT 6.290 103.680 91.665 103.805 ;
      LAYER Pwell ;
        RECT 6.290 100.160 793.390 103.680 ;
      LAYER Nwell ;
        RECT 6.290 100.035 34.545 100.160 ;
        RECT 6.290 95.965 793.390 100.035 ;
        RECT 6.290 95.840 71.505 95.965 ;
      LAYER Pwell ;
        RECT 6.290 92.320 793.390 95.840 ;
      LAYER Nwell ;
        RECT 6.290 92.195 139.265 92.320 ;
        RECT 6.290 88.125 793.390 92.195 ;
        RECT 6.290 88.000 44.065 88.125 ;
      LAYER Pwell ;
        RECT 6.290 84.480 793.390 88.000 ;
      LAYER Nwell ;
        RECT 6.290 84.355 38.680 84.480 ;
        RECT 6.290 80.285 793.390 84.355 ;
        RECT 6.290 80.160 71.505 80.285 ;
      LAYER Pwell ;
        RECT 6.290 76.640 793.390 80.160 ;
      LAYER Nwell ;
        RECT 6.290 76.515 93.345 76.640 ;
        RECT 6.290 72.445 793.390 76.515 ;
        RECT 6.290 72.320 128.625 72.445 ;
      LAYER Pwell ;
        RECT 6.290 68.800 793.390 72.320 ;
      LAYER Nwell ;
        RECT 6.290 68.675 108.680 68.800 ;
        RECT 6.290 64.605 793.390 68.675 ;
        RECT 6.290 64.480 49.105 64.605 ;
      LAYER Pwell ;
        RECT 6.290 60.960 793.390 64.480 ;
      LAYER Nwell ;
        RECT 6.290 60.835 51.905 60.960 ;
        RECT 6.290 56.765 793.390 60.835 ;
        RECT 6.290 56.640 171.745 56.765 ;
      LAYER Pwell ;
        RECT 6.290 53.120 793.390 56.640 ;
      LAYER Nwell ;
        RECT 6.290 52.995 103.425 53.120 ;
        RECT 6.290 48.925 793.390 52.995 ;
        RECT 6.290 48.800 54.145 48.925 ;
      LAYER Pwell ;
        RECT 6.290 45.280 793.390 48.800 ;
      LAYER Nwell ;
        RECT 6.290 45.155 56.385 45.280 ;
        RECT 6.290 41.085 793.390 45.155 ;
        RECT 6.290 40.960 79.905 41.085 ;
      LAYER Pwell ;
        RECT 6.290 37.440 793.390 40.960 ;
      LAYER Nwell ;
        RECT 6.290 37.315 181.825 37.440 ;
        RECT 6.290 33.245 793.390 37.315 ;
        RECT 6.290 33.120 71.505 33.245 ;
      LAYER Pwell ;
        RECT 6.290 29.600 793.390 33.120 ;
      LAYER Nwell ;
        RECT 6.290 29.475 98.945 29.600 ;
        RECT 6.290 25.405 793.390 29.475 ;
        RECT 6.290 25.280 86.065 25.405 ;
      LAYER Pwell ;
        RECT 6.290 21.760 793.390 25.280 ;
      LAYER Nwell ;
        RECT 6.290 21.635 70.945 21.760 ;
        RECT 6.290 17.565 793.390 21.635 ;
        RECT 6.290 17.440 165.025 17.565 ;
      LAYER Pwell ;
        RECT 6.290 15.250 793.390 17.440 ;
      LAYER Metal1 ;
        RECT 6.720 15.380 792.960 334.170 ;
      LAYER Metal2 ;
        RECT 9.660 2.890 792.820 339.830 ;
      LAYER Metal3 ;
        RECT 9.610 327.900 796.000 339.780 ;
        RECT 9.610 326.740 795.700 327.900 ;
        RECT 9.610 320.060 796.000 326.740 ;
        RECT 9.610 318.900 795.700 320.060 ;
        RECT 9.610 312.220 796.000 318.900 ;
        RECT 9.610 311.060 795.700 312.220 ;
        RECT 9.610 304.380 796.000 311.060 ;
        RECT 9.610 303.220 795.700 304.380 ;
        RECT 9.610 296.540 796.000 303.220 ;
        RECT 9.610 295.380 795.700 296.540 ;
        RECT 9.610 288.700 796.000 295.380 ;
        RECT 9.610 287.540 795.700 288.700 ;
        RECT 9.610 280.860 796.000 287.540 ;
        RECT 9.610 279.700 795.700 280.860 ;
        RECT 9.610 273.020 796.000 279.700 ;
        RECT 9.610 271.860 795.700 273.020 ;
        RECT 9.610 265.180 796.000 271.860 ;
        RECT 9.610 264.020 795.700 265.180 ;
        RECT 9.610 257.340 796.000 264.020 ;
        RECT 9.610 256.180 795.700 257.340 ;
        RECT 9.610 249.500 796.000 256.180 ;
        RECT 9.610 248.340 795.700 249.500 ;
        RECT 9.610 241.660 796.000 248.340 ;
        RECT 9.610 240.500 795.700 241.660 ;
        RECT 9.610 233.820 796.000 240.500 ;
        RECT 9.610 232.660 795.700 233.820 ;
        RECT 9.610 225.980 796.000 232.660 ;
        RECT 9.610 224.820 795.700 225.980 ;
        RECT 9.610 218.140 796.000 224.820 ;
        RECT 9.610 216.980 795.700 218.140 ;
        RECT 9.610 210.300 796.000 216.980 ;
        RECT 9.610 209.140 795.700 210.300 ;
        RECT 9.610 202.460 796.000 209.140 ;
        RECT 9.610 201.300 795.700 202.460 ;
        RECT 9.610 194.620 796.000 201.300 ;
        RECT 9.610 193.460 795.700 194.620 ;
        RECT 9.610 186.780 796.000 193.460 ;
        RECT 9.610 185.620 795.700 186.780 ;
        RECT 9.610 178.940 796.000 185.620 ;
        RECT 9.610 177.780 795.700 178.940 ;
        RECT 9.610 171.100 796.000 177.780 ;
        RECT 9.610 169.940 795.700 171.100 ;
        RECT 9.610 163.260 796.000 169.940 ;
        RECT 9.610 162.100 795.700 163.260 ;
        RECT 9.610 155.420 796.000 162.100 ;
        RECT 9.610 154.260 795.700 155.420 ;
        RECT 9.610 147.580 796.000 154.260 ;
        RECT 9.610 146.420 795.700 147.580 ;
        RECT 9.610 139.740 796.000 146.420 ;
        RECT 9.610 138.580 795.700 139.740 ;
        RECT 9.610 131.900 796.000 138.580 ;
        RECT 9.610 130.740 795.700 131.900 ;
        RECT 9.610 124.060 796.000 130.740 ;
        RECT 9.610 122.900 795.700 124.060 ;
        RECT 9.610 116.220 796.000 122.900 ;
        RECT 9.610 115.060 795.700 116.220 ;
        RECT 9.610 108.380 796.000 115.060 ;
        RECT 9.610 107.220 795.700 108.380 ;
        RECT 9.610 100.540 796.000 107.220 ;
        RECT 9.610 99.380 795.700 100.540 ;
        RECT 9.610 92.700 796.000 99.380 ;
        RECT 9.610 91.540 795.700 92.700 ;
        RECT 9.610 84.860 796.000 91.540 ;
        RECT 9.610 83.700 795.700 84.860 ;
        RECT 9.610 77.020 796.000 83.700 ;
        RECT 9.610 75.860 795.700 77.020 ;
        RECT 9.610 69.180 796.000 75.860 ;
        RECT 9.610 68.020 795.700 69.180 ;
        RECT 9.610 61.340 796.000 68.020 ;
        RECT 9.610 60.180 795.700 61.340 ;
        RECT 9.610 53.500 796.000 60.180 ;
        RECT 9.610 52.340 795.700 53.500 ;
        RECT 9.610 45.660 796.000 52.340 ;
        RECT 9.610 44.500 795.700 45.660 ;
        RECT 9.610 37.820 796.000 44.500 ;
        RECT 9.610 36.660 795.700 37.820 ;
        RECT 9.610 29.980 796.000 36.660 ;
        RECT 9.610 28.820 795.700 29.980 ;
        RECT 9.610 22.140 796.000 28.820 ;
        RECT 9.610 20.980 795.700 22.140 ;
        RECT 9.610 2.940 796.000 20.980 ;
      LAYER Metal4 ;
        RECT 48.300 333.800 778.820 337.590 ;
        RECT 48.300 15.080 98.740 333.800 ;
        RECT 100.940 15.080 175.540 333.800 ;
        RECT 177.740 15.080 252.340 333.800 ;
        RECT 254.540 15.080 329.140 333.800 ;
        RECT 331.340 15.080 405.940 333.800 ;
        RECT 408.140 15.080 482.740 333.800 ;
        RECT 484.940 15.080 559.540 333.800 ;
        RECT 561.740 15.080 636.340 333.800 ;
        RECT 638.540 15.080 713.140 333.800 ;
        RECT 715.340 15.080 778.820 333.800 ;
        RECT 48.300 3.450 778.820 15.080 ;
  END
END int_ram
END LIBRARY

