VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO uprj_w_const
  CLASS BLOCK ;
  FOREIGN uprj_w_const ;
  ORIGIN 0.000 0.000 ;
  SIZE 150.000 BY 150.000 ;
  PIN b0_drv[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 146.000 35.790 150.000 ;
    END
  END b0_drv[0]
  PIN b0_drv[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.040 4.000 85.640 ;
    END
  END b0_drv[10]
  PIN b0_drv[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 146.000 148.490 150.000 ;
    END
  END b0_drv[11]
  PIN b0_drv[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END b0_drv[12]
  PIN b0_drv[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END b0_drv[13]
  PIN b0_drv[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 47.640 150.000 48.240 ;
    END
  END b0_drv[14]
  PIN b0_drv[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 125.840 150.000 126.440 ;
    END
  END b0_drv[15]
  PIN b0_drv[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 85.040 150.000 85.640 ;
    END
  END b0_drv[16]
  PIN b0_drv[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 146.000 96.970 150.000 ;
    END
  END b0_drv[17]
  PIN b0_drv[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 20.440 150.000 21.040 ;
    END
  END b0_drv[18]
  PIN b0_drv[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 95.240 150.000 95.840 ;
    END
  END b0_drv[19]
  PIN b0_drv[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END b0_drv[1]
  PIN b0_drv[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 146.000 119.510 150.000 ;
    END
  END b0_drv[20]
  PIN b0_drv[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END b0_drv[21]
  PIN b0_drv[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END b0_drv[22]
  PIN b0_drv[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 146.000 142.050 150.000 ;
    END
  END b0_drv[23]
  PIN b0_drv[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END b0_drv[24]
  PIN b0_drv[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 146.000 29.350 150.000 ;
    END
  END b0_drv[25]
  PIN b0_drv[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 146.000 3.590 150.000 ;
    END
  END b0_drv[26]
  PIN b0_drv[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 146.000 67.990 150.000 ;
    END
  END b0_drv[27]
  PIN b0_drv[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 54.440 150.000 55.040 ;
    END
  END b0_drv[28]
  PIN b0_drv[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 13.640 150.000 14.240 ;
    END
  END b0_drv[29]
  PIN b0_drv[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END b0_drv[2]
  PIN b0_drv[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 136.040 150.000 136.640 ;
    END
  END b0_drv[30]
  PIN b0_drv[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 146.000 80.870 150.000 ;
    END
  END b0_drv[31]
  PIN b0_drv[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 146.000 58.330 150.000 ;
    END
  END b0_drv[32]
  PIN b0_drv[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END b0_drv[33]
  PIN b0_drv[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 146.000 90.530 150.000 ;
    END
  END b0_drv[34]
  PIN b0_drv[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END b0_drv[35]
  PIN b0_drv[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END b0_drv[36]
  PIN b0_drv[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END b0_drv[37]
  PIN b0_drv[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 119.040 150.000 119.640 ;
    END
  END b0_drv[38]
  PIN b0_drv[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 146.000 129.170 150.000 ;
    END
  END b0_drv[39]
  PIN b0_drv[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END b0_drv[3]
  PIN b0_drv[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 146.000 84.090 150.000 ;
    END
  END b0_drv[40]
  PIN b0_drv[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END b0_drv[41]
  PIN b0_drv[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 34.040 150.000 34.640 ;
    END
  END b0_drv[42]
  PIN b0_drv[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 146.000 39.010 150.000 ;
    END
  END b0_drv[43]
  PIN b0_drv[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 6.840 150.000 7.440 ;
    END
  END b0_drv[44]
  PIN b0_drv[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END b0_drv[45]
  PIN b0_drv[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END b0_drv[46]
  PIN b0_drv[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END b0_drv[47]
  PIN b0_drv[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 146.000 135.610 150.000 ;
    END
  END b0_drv[48]
  PIN b0_drv[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 146.000 71.210 150.000 ;
    END
  END b0_drv[49]
  PIN b0_drv[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 139.440 4.000 140.040 ;
    END
  END b0_drv[4]
  PIN b0_drv[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 0.040 150.000 0.640 ;
    END
  END b0_drv[50]
  PIN b0_drv[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END b0_drv[51]
  PIN b0_drv[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END b0_drv[52]
  PIN b0_drv[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END b0_drv[53]
  PIN b0_drv[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END b0_drv[54]
  PIN b0_drv[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 146.000 61.550 150.000 ;
    END
  END b0_drv[55]
  PIN b0_drv[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 146.000 87.310 150.000 ;
    END
  END b0_drv[56]
  PIN b0_drv[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END b0_drv[57]
  PIN b0_drv[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END b0_drv[58]
  PIN b0_drv[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 122.440 150.000 123.040 ;
    END
  END b0_drv[59]
  PIN b0_drv[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 146.000 13.250 150.000 ;
    END
  END b0_drv[5]
  PIN b0_drv[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END b0_drv[60]
  PIN b0_drv[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END b0_drv[61]
  PIN b0_drv[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END b0_drv[62]
  PIN b0_drv[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 78.240 150.000 78.840 ;
    END
  END b0_drv[63]
  PIN b0_drv[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 146.000 64.770 150.000 ;
    END
  END b0_drv[64]
  PIN b0_drv[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 108.840 150.000 109.440 ;
    END
  END b0_drv[65]
  PIN b0_drv[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 146.000 132.390 150.000 ;
    END
  END b0_drv[66]
  PIN b0_drv[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END b0_drv[67]
  PIN b0_drv[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 146.000 122.730 150.000 ;
    END
  END b0_drv[68]
  PIN b0_drv[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END b0_drv[69]
  PIN b0_drv[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 146.000 48.670 150.000 ;
    END
  END b0_drv[6]
  PIN b0_drv[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END b0_drv[70]
  PIN b0_drv[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 57.840 150.000 58.440 ;
    END
  END b0_drv[71]
  PIN b0_drv[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 10.240 150.000 10.840 ;
    END
  END b0_drv[72]
  PIN b0_drv[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END b0_drv[73]
  PIN b0_drv[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 139.440 150.000 140.040 ;
    END
  END b0_drv[74]
  PIN b0_drv[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 105.440 150.000 106.040 ;
    END
  END b0_drv[75]
  PIN b0_drv[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END b0_drv[76]
  PIN b0_drv[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END b0_drv[77]
  PIN b0_drv[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END b0_drv[78]
  PIN b0_drv[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END b0_drv[79]
  PIN b0_drv[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 64.640 150.000 65.240 ;
    END
  END b0_drv[7]
  PIN b0_drv[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END b0_drv[80]
  PIN b0_drv[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 0.000 6.810 4.000 ;
    END
  END b0_drv[81]
  PIN b0_drv[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END b0_drv[82]
  PIN b0_drv[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END b0_drv[8]
  PIN b0_drv[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END b0_drv[9]
  PIN cw_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END cw_clk_i
  PIN cw_clk_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 146.000 116.290 150.000 ;
    END
  END cw_clk_o
  PIN cw_dir
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END cw_dir
  PIN cw_dir_b_o
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END cw_dir_b_o
  PIN cw_dir_b_oo
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 68.040 150.000 68.640 ;
    END
  END cw_dir_b_oo
  PIN cw_dir_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 37.440 150.000 38.040 ;
    END
  END cw_dir_o
  PIN cw_req_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 146.000 138.830 150.000 ;
    END
  END cw_req_i
  PIN cw_req_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END cw_req_o
  PIN cw_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END cw_rst_i
  PIN cw_rst_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 129.240 150.000 129.840 ;
    END
  END cw_rst_o
  PIN io_oeb_15_0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END io_oeb_15_0[0]
  PIN io_oeb_15_0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END io_oeb_15_0[10]
  PIN io_oeb_15_0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 146.000 26.130 150.000 ;
    END
  END io_oeb_15_0[11]
  PIN io_oeb_15_0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 146.000 32.570 150.000 ;
    END
  END io_oeb_15_0[12]
  PIN io_oeb_15_0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 146.000 6.810 150.000 ;
    END
  END io_oeb_15_0[13]
  PIN io_oeb_15_0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END io_oeb_15_0[14]
  PIN io_oeb_15_0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 74.840 150.000 75.440 ;
    END
  END io_oeb_15_0[15]
  PIN io_oeb_15_0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END io_oeb_15_0[1]
  PIN io_oeb_15_0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 146.000 55.110 150.000 ;
    END
  END io_oeb_15_0[2]
  PIN io_oeb_15_0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 81.640 150.000 82.240 ;
    END
  END io_oeb_15_0[3]
  PIN io_oeb_15_0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END io_oeb_15_0[4]
  PIN io_oeb_15_0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END io_oeb_15_0[5]
  PIN io_oeb_15_0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END io_oeb_15_0[6]
  PIN io_oeb_15_0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END io_oeb_15_0[7]
  PIN io_oeb_15_0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 132.640 4.000 133.240 ;
    END
  END io_oeb_15_0[8]
  PIN io_oeb_15_0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 142.840 150.000 143.440 ;
    END
  END io_oeb_15_0[9]
  PIN io_oeb_18_16[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END io_oeb_18_16[0]
  PIN io_oeb_18_16[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END io_oeb_18_16[1]
  PIN io_oeb_18_16[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 146.000 100.190 150.000 ;
    END
  END io_oeb_18_16[2]
  PIN io_oeb_20_19[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 146.000 93.750 150.000 ;
    END
  END io_oeb_20_19[0]
  PIN io_oeb_20_19[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END io_oeb_20_19[1]
  PIN io_oeb_21
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END io_oeb_21
  PIN io_oeb_22
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 17.040 150.000 17.640 ;
    END
  END io_oeb_22
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 115.640 150.000 116.240 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 146.000 42.230 150.000 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 30.640 150.000 31.240 ;
    END
  END io_out[14]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 88.440 150.000 89.040 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 146.000 45.450 150.000 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 61.240 150.000 61.840 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 146.000 10.030 150.000 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 0.000 80.870 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 112.240 150.000 112.840 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 146.000 113.070 150.000 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 40.840 150.000 41.440 ;
    END
  END io_out[9]
  PIN io_out_20_19[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END io_out_20_19[0]
  PIN io_out_20_19[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 3.440 150.000 4.040 ;
    END
  END io_out_20_19[1]
  PIN io_out_22
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 146.000 16.470 150.000 ;
    END
  END io_out_22
  PIN la_data_out_16_17[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 0.000 125.950 4.000 ;
    END
  END la_data_out_16_17[0]
  PIN la_data_out_16_17[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END la_data_out_16_17[1]
  PIN la_data_out_21
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END la_data_out_21
  PIN la_data_out_37_36[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 27.240 150.000 27.840 ;
    END
  END la_data_out_37_36[0]
  PIN la_data_out_37_36[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 132.640 150.000 133.240 ;
    END
  END la_data_out_37_36[1]
  PIN la_data_out_77_62[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 91.840 150.000 92.440 ;
    END
  END la_data_out_77_62[0]
  PIN la_data_out_77_62[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END la_data_out_77_62[10]
  PIN la_data_out_77_62[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END la_data_out_77_62[11]
  PIN la_data_out_77_62[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 51.040 150.000 51.640 ;
    END
  END la_data_out_77_62[12]
  PIN la_data_out_77_62[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END la_data_out_77_62[13]
  PIN la_data_out_77_62[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END la_data_out_77_62[14]
  PIN la_data_out_77_62[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 146.240 150.000 146.840 ;
    END
  END la_data_out_77_62[15]
  PIN la_data_out_77_62[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END la_data_out_77_62[1]
  PIN la_data_out_77_62[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 146.000 145.270 150.000 ;
    END
  END la_data_out_77_62[2]
  PIN la_data_out_77_62[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END la_data_out_77_62[3]
  PIN la_data_out_77_62[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END la_data_out_77_62[4]
  PIN la_data_out_77_62[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END la_data_out_77_62[5]
  PIN la_data_out_77_62[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END la_data_out_77_62[6]
  PIN la_data_out_77_62[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 13.640 4.000 14.240 ;
    END
  END la_data_out_77_62[7]
  PIN la_data_out_77_62[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END la_data_out_77_62[8]
  PIN la_data_out_77_62[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 146.000 19.690 150.000 ;
    END
  END la_data_out_77_62[9]
  PIN la_data_out_97_95[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 146.000 77.650 150.000 ;
    END
  END la_data_out_97_95[0]
  PIN la_data_out_97_95[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END la_data_out_97_95[1]
  PIN la_data_out_97_95[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END la_data_out_97_95[2]
  PIN la_datb_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END la_datb_i[0]
  PIN la_datb_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 146.000 103.410 150.000 ;
    END
  END la_datb_i[1]
  PIN la_datb_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 146.000 74.430 150.000 ;
    END
  END la_datb_i[2]
  PIN la_datb_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END la_datb_o[0]
  PIN la_datb_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 146.000 125.950 150.000 ;
    END
  END la_datb_o[1]
  PIN la_datb_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 23.840 150.000 24.440 ;
    END
  END la_datb_o[2]
  PIN oeb_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END oeb_out[0]
  PIN oeb_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 102.040 150.000 102.640 ;
    END
  END oeb_out[10]
  PIN oeb_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 29.070 0.000 29.350 4.000 ;
    END
  END oeb_out[11]
  PIN oeb_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END oeb_out[12]
  PIN oeb_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 30.640 4.000 31.240 ;
    END
  END oeb_out[13]
  PIN oeb_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 98.640 150.000 99.240 ;
    END
  END oeb_out[14]
  PIN oeb_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END oeb_out[1]
  PIN oeb_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 146.000 109.850 150.000 ;
    END
  END oeb_out[2]
  PIN oeb_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 146.000 106.630 150.000 ;
    END
  END oeb_out[3]
  PIN oeb_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 146.000 0.370 150.000 ;
    END
  END oeb_out[4]
  PIN oeb_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 146.000 22.910 150.000 ;
    END
  END oeb_out[5]
  PIN oeb_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 0.000 103.410 4.000 ;
    END
  END oeb_out[6]
  PIN oeb_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END oeb_out[7]
  PIN oeb_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END oeb_out[8]
  PIN oeb_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 146.000 71.440 150.000 72.040 ;
    END
  END oeb_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 22.090 10.640 23.690 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.830 10.640 58.430 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 91.570 10.640 93.170 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 126.310 10.640 127.910 138.960 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 39.460 10.640 41.060 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 74.200 10.640 75.800 138.960 ;
    END
    PORT
      LAYER met4 ;
        RECT 108.940 10.640 110.540 138.960 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 144.440 138.805 ;
      LAYER met1 ;
        RECT 0.070 10.640 148.510 138.960 ;
      LAYER met2 ;
        RECT 0.650 145.720 3.030 146.725 ;
        RECT 3.870 145.720 6.250 146.725 ;
        RECT 7.090 145.720 9.470 146.725 ;
        RECT 10.310 145.720 12.690 146.725 ;
        RECT 13.530 145.720 15.910 146.725 ;
        RECT 16.750 145.720 19.130 146.725 ;
        RECT 19.970 145.720 22.350 146.725 ;
        RECT 23.190 145.720 25.570 146.725 ;
        RECT 26.410 145.720 28.790 146.725 ;
        RECT 29.630 145.720 32.010 146.725 ;
        RECT 32.850 145.720 35.230 146.725 ;
        RECT 36.070 145.720 38.450 146.725 ;
        RECT 39.290 145.720 41.670 146.725 ;
        RECT 42.510 145.720 44.890 146.725 ;
        RECT 45.730 145.720 48.110 146.725 ;
        RECT 48.950 145.720 54.550 146.725 ;
        RECT 55.390 145.720 57.770 146.725 ;
        RECT 58.610 145.720 60.990 146.725 ;
        RECT 61.830 145.720 64.210 146.725 ;
        RECT 65.050 145.720 67.430 146.725 ;
        RECT 68.270 145.720 70.650 146.725 ;
        RECT 71.490 145.720 73.870 146.725 ;
        RECT 74.710 145.720 77.090 146.725 ;
        RECT 77.930 145.720 80.310 146.725 ;
        RECT 81.150 145.720 83.530 146.725 ;
        RECT 84.370 145.720 86.750 146.725 ;
        RECT 87.590 145.720 89.970 146.725 ;
        RECT 90.810 145.720 93.190 146.725 ;
        RECT 94.030 145.720 96.410 146.725 ;
        RECT 97.250 145.720 99.630 146.725 ;
        RECT 100.470 145.720 102.850 146.725 ;
        RECT 103.690 145.720 106.070 146.725 ;
        RECT 106.910 145.720 109.290 146.725 ;
        RECT 110.130 145.720 112.510 146.725 ;
        RECT 113.350 145.720 115.730 146.725 ;
        RECT 116.570 145.720 118.950 146.725 ;
        RECT 119.790 145.720 122.170 146.725 ;
        RECT 123.010 145.720 125.390 146.725 ;
        RECT 126.230 145.720 128.610 146.725 ;
        RECT 129.450 145.720 131.830 146.725 ;
        RECT 132.670 145.720 135.050 146.725 ;
        RECT 135.890 145.720 138.270 146.725 ;
        RECT 139.110 145.720 141.490 146.725 ;
        RECT 142.330 145.720 144.710 146.725 ;
        RECT 145.550 145.720 147.930 146.725 ;
        RECT 0.100 4.280 148.480 145.720 ;
        RECT 0.650 0.155 3.030 4.280 ;
        RECT 3.870 0.155 6.250 4.280 ;
        RECT 7.090 0.155 9.470 4.280 ;
        RECT 10.310 0.155 12.690 4.280 ;
        RECT 13.530 0.155 15.910 4.280 ;
        RECT 16.750 0.155 19.130 4.280 ;
        RECT 19.970 0.155 22.350 4.280 ;
        RECT 23.190 0.155 25.570 4.280 ;
        RECT 26.410 0.155 28.790 4.280 ;
        RECT 29.630 0.155 32.010 4.280 ;
        RECT 32.850 0.155 35.230 4.280 ;
        RECT 36.070 0.155 38.450 4.280 ;
        RECT 39.290 0.155 41.670 4.280 ;
        RECT 42.510 0.155 44.890 4.280 ;
        RECT 45.730 0.155 48.110 4.280 ;
        RECT 48.950 0.155 51.330 4.280 ;
        RECT 52.170 0.155 54.550 4.280 ;
        RECT 55.390 0.155 57.770 4.280 ;
        RECT 58.610 0.155 60.990 4.280 ;
        RECT 61.830 0.155 64.210 4.280 ;
        RECT 65.050 0.155 67.430 4.280 ;
        RECT 68.270 0.155 70.650 4.280 ;
        RECT 71.490 0.155 73.870 4.280 ;
        RECT 74.710 0.155 77.090 4.280 ;
        RECT 77.930 0.155 80.310 4.280 ;
        RECT 81.150 0.155 83.530 4.280 ;
        RECT 84.370 0.155 86.750 4.280 ;
        RECT 87.590 0.155 89.970 4.280 ;
        RECT 90.810 0.155 93.190 4.280 ;
        RECT 94.030 0.155 96.410 4.280 ;
        RECT 97.250 0.155 99.630 4.280 ;
        RECT 100.470 0.155 102.850 4.280 ;
        RECT 103.690 0.155 106.070 4.280 ;
        RECT 106.910 0.155 109.290 4.280 ;
        RECT 110.130 0.155 112.510 4.280 ;
        RECT 113.350 0.155 115.730 4.280 ;
        RECT 116.570 0.155 118.950 4.280 ;
        RECT 119.790 0.155 122.170 4.280 ;
        RECT 123.010 0.155 125.390 4.280 ;
        RECT 126.230 0.155 128.610 4.280 ;
        RECT 129.450 0.155 131.830 4.280 ;
        RECT 132.670 0.155 135.050 4.280 ;
        RECT 135.890 0.155 138.270 4.280 ;
        RECT 139.110 0.155 141.490 4.280 ;
        RECT 142.330 0.155 144.710 4.280 ;
        RECT 145.550 0.155 147.930 4.280 ;
      LAYER met3 ;
        RECT 4.400 145.840 145.600 146.705 ;
        RECT 4.000 143.840 146.000 145.840 ;
        RECT 4.400 142.440 145.600 143.840 ;
        RECT 4.000 140.440 146.000 142.440 ;
        RECT 4.400 139.040 145.600 140.440 ;
        RECT 4.000 137.040 146.000 139.040 ;
        RECT 4.400 135.640 145.600 137.040 ;
        RECT 4.000 133.640 146.000 135.640 ;
        RECT 4.400 132.240 145.600 133.640 ;
        RECT 4.000 130.240 146.000 132.240 ;
        RECT 4.400 128.840 145.600 130.240 ;
        RECT 4.000 126.840 146.000 128.840 ;
        RECT 4.400 125.440 145.600 126.840 ;
        RECT 4.000 123.440 146.000 125.440 ;
        RECT 4.400 122.040 145.600 123.440 ;
        RECT 4.000 120.040 146.000 122.040 ;
        RECT 4.400 118.640 145.600 120.040 ;
        RECT 4.000 116.640 146.000 118.640 ;
        RECT 4.400 115.240 145.600 116.640 ;
        RECT 4.000 113.240 146.000 115.240 ;
        RECT 4.400 111.840 145.600 113.240 ;
        RECT 4.000 109.840 146.000 111.840 ;
        RECT 4.400 108.440 145.600 109.840 ;
        RECT 4.000 106.440 146.000 108.440 ;
        RECT 4.400 105.040 145.600 106.440 ;
        RECT 4.000 103.040 146.000 105.040 ;
        RECT 4.400 101.640 145.600 103.040 ;
        RECT 4.000 99.640 146.000 101.640 ;
        RECT 4.400 98.240 145.600 99.640 ;
        RECT 4.000 96.240 146.000 98.240 ;
        RECT 4.400 94.840 145.600 96.240 ;
        RECT 4.000 92.840 146.000 94.840 ;
        RECT 4.400 91.440 145.600 92.840 ;
        RECT 4.000 89.440 146.000 91.440 ;
        RECT 4.400 88.040 145.600 89.440 ;
        RECT 4.000 86.040 146.000 88.040 ;
        RECT 4.400 84.640 145.600 86.040 ;
        RECT 4.000 82.640 146.000 84.640 ;
        RECT 4.400 81.240 145.600 82.640 ;
        RECT 4.000 79.240 146.000 81.240 ;
        RECT 4.400 77.840 145.600 79.240 ;
        RECT 4.000 75.840 146.000 77.840 ;
        RECT 4.400 74.440 145.600 75.840 ;
        RECT 4.000 72.440 146.000 74.440 ;
        RECT 4.400 71.040 145.600 72.440 ;
        RECT 4.000 69.040 146.000 71.040 ;
        RECT 4.400 67.640 145.600 69.040 ;
        RECT 4.000 65.640 146.000 67.640 ;
        RECT 4.400 64.240 145.600 65.640 ;
        RECT 4.000 62.240 146.000 64.240 ;
        RECT 4.400 60.840 145.600 62.240 ;
        RECT 4.000 58.840 146.000 60.840 ;
        RECT 4.400 57.440 145.600 58.840 ;
        RECT 4.000 55.440 146.000 57.440 ;
        RECT 4.400 54.040 145.600 55.440 ;
        RECT 4.000 52.040 146.000 54.040 ;
        RECT 4.400 50.640 145.600 52.040 ;
        RECT 4.000 48.640 146.000 50.640 ;
        RECT 4.400 47.240 145.600 48.640 ;
        RECT 4.000 45.240 146.000 47.240 ;
        RECT 4.400 43.840 146.000 45.240 ;
        RECT 4.000 41.840 146.000 43.840 ;
        RECT 4.400 40.440 145.600 41.840 ;
        RECT 4.000 38.440 146.000 40.440 ;
        RECT 4.400 37.040 145.600 38.440 ;
        RECT 4.000 35.040 146.000 37.040 ;
        RECT 4.400 33.640 145.600 35.040 ;
        RECT 4.000 31.640 146.000 33.640 ;
        RECT 4.400 30.240 145.600 31.640 ;
        RECT 4.000 28.240 146.000 30.240 ;
        RECT 4.400 26.840 145.600 28.240 ;
        RECT 4.000 24.840 146.000 26.840 ;
        RECT 4.400 23.440 145.600 24.840 ;
        RECT 4.000 21.440 146.000 23.440 ;
        RECT 4.400 20.040 145.600 21.440 ;
        RECT 4.000 18.040 146.000 20.040 ;
        RECT 4.400 16.640 145.600 18.040 ;
        RECT 4.000 14.640 146.000 16.640 ;
        RECT 4.400 13.240 145.600 14.640 ;
        RECT 4.000 11.240 146.000 13.240 ;
        RECT 4.400 9.840 145.600 11.240 ;
        RECT 4.000 7.840 146.000 9.840 ;
        RECT 4.400 6.440 145.600 7.840 ;
        RECT 4.000 4.440 146.000 6.440 ;
        RECT 4.400 3.040 145.600 4.440 ;
        RECT 4.000 1.040 146.000 3.040 ;
        RECT 4.000 0.175 145.600 1.040 ;
  END
END uprj_w_const
END LIBRARY

