magic
tech gf180mcuD
magscale 1 5
timestamp 1700070097
<< obsm1 >>
rect 672 463 119280 35310
<< metal2 >>
rect 3024 36600 3080 37000
rect 3920 36600 3976 37000
rect 4816 36600 4872 37000
rect 5712 36600 5768 37000
rect 6608 36600 6664 37000
rect 7504 36600 7560 37000
rect 8400 36600 8456 37000
rect 9296 36600 9352 37000
rect 10192 36600 10248 37000
rect 11088 36600 11144 37000
rect 11984 36600 12040 37000
rect 12880 36600 12936 37000
rect 13776 36600 13832 37000
rect 14672 36600 14728 37000
rect 15568 36600 15624 37000
rect 16464 36600 16520 37000
rect 17360 36600 17416 37000
rect 18256 36600 18312 37000
rect 19152 36600 19208 37000
rect 20048 36600 20104 37000
rect 20944 36600 21000 37000
rect 21840 36600 21896 37000
rect 22736 36600 22792 37000
rect 23632 36600 23688 37000
rect 24528 36600 24584 37000
rect 25424 36600 25480 37000
rect 26320 36600 26376 37000
rect 27216 36600 27272 37000
rect 28112 36600 28168 37000
rect 29008 36600 29064 37000
rect 29904 36600 29960 37000
rect 30800 36600 30856 37000
rect 31696 36600 31752 37000
rect 32592 36600 32648 37000
rect 33488 36600 33544 37000
rect 34384 36600 34440 37000
rect 35280 36600 35336 37000
rect 36176 36600 36232 37000
rect 37072 36600 37128 37000
rect 37968 36600 38024 37000
rect 38864 36600 38920 37000
rect 39760 36600 39816 37000
rect 40656 36600 40712 37000
rect 41552 36600 41608 37000
rect 42448 36600 42504 37000
rect 43344 36600 43400 37000
rect 44240 36600 44296 37000
rect 45136 36600 45192 37000
rect 46032 36600 46088 37000
rect 46928 36600 46984 37000
rect 47824 36600 47880 37000
rect 48720 36600 48776 37000
rect 49616 36600 49672 37000
rect 50512 36600 50568 37000
rect 51408 36600 51464 37000
rect 52304 36600 52360 37000
rect 53200 36600 53256 37000
rect 54096 36600 54152 37000
rect 54992 36600 55048 37000
rect 55888 36600 55944 37000
rect 56784 36600 56840 37000
rect 57680 36600 57736 37000
rect 58576 36600 58632 37000
rect 59472 36600 59528 37000
rect 60368 36600 60424 37000
rect 61264 36600 61320 37000
rect 62160 36600 62216 37000
rect 63056 36600 63112 37000
rect 63952 36600 64008 37000
rect 64848 36600 64904 37000
rect 65744 36600 65800 37000
rect 66640 36600 66696 37000
rect 67536 36600 67592 37000
rect 68432 36600 68488 37000
rect 69328 36600 69384 37000
rect 70224 36600 70280 37000
rect 71120 36600 71176 37000
rect 72016 36600 72072 37000
rect 72912 36600 72968 37000
rect 73808 36600 73864 37000
rect 74704 36600 74760 37000
rect 75600 36600 75656 37000
rect 76496 36600 76552 37000
rect 77392 36600 77448 37000
rect 78288 36600 78344 37000
rect 79184 36600 79240 37000
rect 80080 36600 80136 37000
rect 80976 36600 81032 37000
rect 81872 36600 81928 37000
rect 82768 36600 82824 37000
rect 83664 36600 83720 37000
rect 84560 36600 84616 37000
rect 85456 36600 85512 37000
rect 86352 36600 86408 37000
rect 87248 36600 87304 37000
rect 88144 36600 88200 37000
rect 89040 36600 89096 37000
rect 89936 36600 89992 37000
rect 90832 36600 90888 37000
rect 91728 36600 91784 37000
rect 92624 36600 92680 37000
rect 93520 36600 93576 37000
rect 94416 36600 94472 37000
rect 95312 36600 95368 37000
rect 96208 36600 96264 37000
rect 97104 36600 97160 37000
rect 98000 36600 98056 37000
rect 98896 36600 98952 37000
rect 99792 36600 99848 37000
rect 100688 36600 100744 37000
rect 101584 36600 101640 37000
rect 102480 36600 102536 37000
rect 103376 36600 103432 37000
rect 104272 36600 104328 37000
rect 105168 36600 105224 37000
rect 106064 36600 106120 37000
rect 106960 36600 107016 37000
rect 107856 36600 107912 37000
rect 108752 36600 108808 37000
rect 109648 36600 109704 37000
rect 110544 36600 110600 37000
rect 111440 36600 111496 37000
rect 112336 36600 112392 37000
rect 113232 36600 113288 37000
rect 114128 36600 114184 37000
rect 115024 36600 115080 37000
rect 115920 36600 115976 37000
rect 116816 36600 116872 37000
rect 8512 0 8568 400
rect 8736 0 8792 400
rect 8960 0 9016 400
rect 9184 0 9240 400
rect 9408 0 9464 400
rect 9632 0 9688 400
rect 9856 0 9912 400
rect 10080 0 10136 400
rect 10304 0 10360 400
rect 10528 0 10584 400
rect 10752 0 10808 400
rect 10976 0 11032 400
rect 11200 0 11256 400
rect 11424 0 11480 400
rect 11648 0 11704 400
rect 11872 0 11928 400
rect 12096 0 12152 400
rect 12320 0 12376 400
rect 12544 0 12600 400
rect 12768 0 12824 400
rect 12992 0 13048 400
rect 13216 0 13272 400
rect 13440 0 13496 400
rect 13664 0 13720 400
rect 13888 0 13944 400
rect 14112 0 14168 400
rect 14336 0 14392 400
rect 14560 0 14616 400
rect 14784 0 14840 400
rect 15008 0 15064 400
rect 15232 0 15288 400
rect 15456 0 15512 400
rect 15680 0 15736 400
rect 15904 0 15960 400
rect 16128 0 16184 400
rect 16352 0 16408 400
rect 16576 0 16632 400
rect 16800 0 16856 400
rect 17024 0 17080 400
rect 17248 0 17304 400
rect 17472 0 17528 400
rect 17696 0 17752 400
rect 17920 0 17976 400
rect 18144 0 18200 400
rect 18368 0 18424 400
rect 18592 0 18648 400
rect 18816 0 18872 400
rect 19040 0 19096 400
rect 19264 0 19320 400
rect 19488 0 19544 400
rect 19712 0 19768 400
rect 19936 0 19992 400
rect 20160 0 20216 400
rect 20384 0 20440 400
rect 20608 0 20664 400
rect 20832 0 20888 400
rect 21056 0 21112 400
rect 21280 0 21336 400
rect 21504 0 21560 400
rect 21728 0 21784 400
rect 21952 0 22008 400
rect 22176 0 22232 400
rect 22400 0 22456 400
rect 22624 0 22680 400
rect 22848 0 22904 400
rect 23072 0 23128 400
rect 23296 0 23352 400
rect 23520 0 23576 400
rect 23744 0 23800 400
rect 23968 0 24024 400
rect 24192 0 24248 400
rect 24416 0 24472 400
rect 24640 0 24696 400
rect 24864 0 24920 400
rect 25088 0 25144 400
rect 25312 0 25368 400
rect 25536 0 25592 400
rect 25760 0 25816 400
rect 25984 0 26040 400
rect 26208 0 26264 400
rect 26432 0 26488 400
rect 26656 0 26712 400
rect 26880 0 26936 400
rect 27104 0 27160 400
rect 27328 0 27384 400
rect 27552 0 27608 400
rect 27776 0 27832 400
rect 28000 0 28056 400
rect 28224 0 28280 400
rect 28448 0 28504 400
rect 28672 0 28728 400
rect 28896 0 28952 400
rect 29120 0 29176 400
rect 29344 0 29400 400
rect 29568 0 29624 400
rect 29792 0 29848 400
rect 30016 0 30072 400
rect 30240 0 30296 400
rect 30464 0 30520 400
rect 30688 0 30744 400
rect 30912 0 30968 400
rect 31136 0 31192 400
rect 31360 0 31416 400
rect 31584 0 31640 400
rect 31808 0 31864 400
rect 32032 0 32088 400
rect 32256 0 32312 400
rect 32480 0 32536 400
rect 32704 0 32760 400
rect 32928 0 32984 400
rect 33152 0 33208 400
rect 33376 0 33432 400
rect 33600 0 33656 400
rect 33824 0 33880 400
rect 34048 0 34104 400
rect 34272 0 34328 400
rect 34496 0 34552 400
rect 34720 0 34776 400
rect 34944 0 35000 400
rect 35168 0 35224 400
rect 35392 0 35448 400
rect 35616 0 35672 400
rect 35840 0 35896 400
rect 36064 0 36120 400
rect 36288 0 36344 400
rect 36512 0 36568 400
rect 36736 0 36792 400
rect 36960 0 37016 400
rect 37184 0 37240 400
rect 37408 0 37464 400
rect 37632 0 37688 400
rect 37856 0 37912 400
rect 38080 0 38136 400
rect 38304 0 38360 400
rect 38528 0 38584 400
rect 38752 0 38808 400
rect 38976 0 39032 400
rect 39200 0 39256 400
rect 39424 0 39480 400
rect 39648 0 39704 400
rect 39872 0 39928 400
rect 40096 0 40152 400
rect 40320 0 40376 400
rect 40544 0 40600 400
rect 40768 0 40824 400
rect 40992 0 41048 400
rect 41216 0 41272 400
rect 41440 0 41496 400
rect 41664 0 41720 400
rect 41888 0 41944 400
rect 42112 0 42168 400
rect 42336 0 42392 400
rect 42560 0 42616 400
rect 42784 0 42840 400
rect 43008 0 43064 400
rect 43232 0 43288 400
rect 43456 0 43512 400
rect 43680 0 43736 400
rect 43904 0 43960 400
rect 44128 0 44184 400
rect 44352 0 44408 400
rect 44576 0 44632 400
rect 44800 0 44856 400
rect 45024 0 45080 400
rect 45248 0 45304 400
rect 45472 0 45528 400
rect 45696 0 45752 400
rect 45920 0 45976 400
rect 46144 0 46200 400
rect 46368 0 46424 400
rect 46592 0 46648 400
rect 46816 0 46872 400
rect 47040 0 47096 400
rect 47264 0 47320 400
rect 47488 0 47544 400
rect 47712 0 47768 400
rect 47936 0 47992 400
rect 48160 0 48216 400
rect 48384 0 48440 400
rect 48608 0 48664 400
rect 48832 0 48888 400
rect 49056 0 49112 400
rect 49280 0 49336 400
rect 49504 0 49560 400
rect 49728 0 49784 400
rect 49952 0 50008 400
rect 50176 0 50232 400
rect 50400 0 50456 400
rect 50624 0 50680 400
rect 50848 0 50904 400
rect 51072 0 51128 400
rect 51296 0 51352 400
rect 51520 0 51576 400
rect 51744 0 51800 400
rect 51968 0 52024 400
rect 52192 0 52248 400
rect 52416 0 52472 400
rect 52640 0 52696 400
rect 52864 0 52920 400
rect 53088 0 53144 400
rect 53312 0 53368 400
rect 53536 0 53592 400
rect 53760 0 53816 400
rect 53984 0 54040 400
rect 54208 0 54264 400
rect 54432 0 54488 400
rect 54656 0 54712 400
rect 54880 0 54936 400
rect 55104 0 55160 400
rect 55328 0 55384 400
rect 55552 0 55608 400
rect 55776 0 55832 400
rect 56000 0 56056 400
rect 56224 0 56280 400
rect 56448 0 56504 400
rect 56672 0 56728 400
rect 56896 0 56952 400
rect 57120 0 57176 400
rect 57344 0 57400 400
rect 57568 0 57624 400
rect 57792 0 57848 400
rect 58016 0 58072 400
rect 58240 0 58296 400
rect 58464 0 58520 400
rect 58688 0 58744 400
rect 58912 0 58968 400
rect 59136 0 59192 400
rect 59360 0 59416 400
rect 59584 0 59640 400
rect 59808 0 59864 400
rect 60032 0 60088 400
rect 60256 0 60312 400
rect 60480 0 60536 400
rect 60704 0 60760 400
rect 60928 0 60984 400
rect 61152 0 61208 400
rect 61376 0 61432 400
rect 61600 0 61656 400
rect 61824 0 61880 400
rect 62048 0 62104 400
rect 62272 0 62328 400
rect 62496 0 62552 400
rect 62720 0 62776 400
rect 62944 0 63000 400
rect 63168 0 63224 400
rect 63392 0 63448 400
rect 63616 0 63672 400
rect 63840 0 63896 400
rect 64064 0 64120 400
rect 64288 0 64344 400
rect 64512 0 64568 400
rect 64736 0 64792 400
rect 64960 0 65016 400
rect 65184 0 65240 400
rect 65408 0 65464 400
rect 65632 0 65688 400
rect 65856 0 65912 400
rect 66080 0 66136 400
rect 66304 0 66360 400
rect 66528 0 66584 400
rect 66752 0 66808 400
rect 66976 0 67032 400
rect 67200 0 67256 400
rect 67424 0 67480 400
rect 67648 0 67704 400
rect 67872 0 67928 400
rect 68096 0 68152 400
rect 68320 0 68376 400
rect 68544 0 68600 400
rect 68768 0 68824 400
rect 68992 0 69048 400
rect 69216 0 69272 400
rect 69440 0 69496 400
rect 69664 0 69720 400
rect 69888 0 69944 400
rect 70112 0 70168 400
rect 70336 0 70392 400
rect 70560 0 70616 400
rect 70784 0 70840 400
rect 71008 0 71064 400
rect 71232 0 71288 400
rect 71456 0 71512 400
rect 71680 0 71736 400
rect 71904 0 71960 400
rect 72128 0 72184 400
rect 72352 0 72408 400
rect 72576 0 72632 400
rect 72800 0 72856 400
rect 73024 0 73080 400
rect 73248 0 73304 400
rect 73472 0 73528 400
rect 73696 0 73752 400
rect 73920 0 73976 400
rect 74144 0 74200 400
rect 74368 0 74424 400
rect 74592 0 74648 400
rect 74816 0 74872 400
rect 75040 0 75096 400
rect 75264 0 75320 400
rect 75488 0 75544 400
rect 75712 0 75768 400
rect 75936 0 75992 400
rect 76160 0 76216 400
rect 76384 0 76440 400
rect 76608 0 76664 400
rect 76832 0 76888 400
rect 77056 0 77112 400
rect 77280 0 77336 400
rect 77504 0 77560 400
rect 77728 0 77784 400
rect 77952 0 78008 400
rect 78176 0 78232 400
rect 78400 0 78456 400
rect 78624 0 78680 400
rect 78848 0 78904 400
rect 79072 0 79128 400
rect 79296 0 79352 400
rect 79520 0 79576 400
rect 79744 0 79800 400
rect 79968 0 80024 400
rect 80192 0 80248 400
rect 80416 0 80472 400
rect 80640 0 80696 400
rect 80864 0 80920 400
rect 81088 0 81144 400
rect 81312 0 81368 400
rect 81536 0 81592 400
rect 81760 0 81816 400
rect 81984 0 82040 400
rect 82208 0 82264 400
rect 82432 0 82488 400
rect 82656 0 82712 400
rect 82880 0 82936 400
rect 83104 0 83160 400
rect 83328 0 83384 400
rect 83552 0 83608 400
rect 83776 0 83832 400
rect 84000 0 84056 400
rect 84224 0 84280 400
rect 84448 0 84504 400
rect 84672 0 84728 400
rect 84896 0 84952 400
rect 85120 0 85176 400
rect 85344 0 85400 400
rect 85568 0 85624 400
rect 85792 0 85848 400
rect 86016 0 86072 400
rect 86240 0 86296 400
rect 86464 0 86520 400
rect 86688 0 86744 400
rect 86912 0 86968 400
rect 87136 0 87192 400
rect 87360 0 87416 400
rect 87584 0 87640 400
rect 87808 0 87864 400
rect 88032 0 88088 400
rect 88256 0 88312 400
rect 88480 0 88536 400
rect 88704 0 88760 400
rect 88928 0 88984 400
rect 89152 0 89208 400
rect 89376 0 89432 400
rect 89600 0 89656 400
rect 89824 0 89880 400
rect 90048 0 90104 400
rect 90272 0 90328 400
rect 90496 0 90552 400
rect 90720 0 90776 400
rect 90944 0 91000 400
rect 91168 0 91224 400
rect 91392 0 91448 400
rect 91616 0 91672 400
rect 91840 0 91896 400
rect 92064 0 92120 400
rect 92288 0 92344 400
rect 92512 0 92568 400
rect 92736 0 92792 400
rect 92960 0 93016 400
rect 93184 0 93240 400
rect 93408 0 93464 400
rect 93632 0 93688 400
rect 93856 0 93912 400
rect 94080 0 94136 400
rect 94304 0 94360 400
rect 94528 0 94584 400
rect 94752 0 94808 400
rect 94976 0 95032 400
rect 95200 0 95256 400
rect 95424 0 95480 400
rect 95648 0 95704 400
rect 95872 0 95928 400
rect 96096 0 96152 400
rect 96320 0 96376 400
rect 96544 0 96600 400
rect 96768 0 96824 400
rect 96992 0 97048 400
rect 97216 0 97272 400
rect 97440 0 97496 400
rect 97664 0 97720 400
rect 97888 0 97944 400
rect 98112 0 98168 400
rect 98336 0 98392 400
rect 98560 0 98616 400
rect 98784 0 98840 400
rect 99008 0 99064 400
rect 99232 0 99288 400
rect 99456 0 99512 400
rect 99680 0 99736 400
rect 99904 0 99960 400
rect 100128 0 100184 400
rect 100352 0 100408 400
rect 100576 0 100632 400
rect 100800 0 100856 400
rect 101024 0 101080 400
rect 101248 0 101304 400
rect 101472 0 101528 400
rect 101696 0 101752 400
rect 101920 0 101976 400
rect 102144 0 102200 400
rect 102368 0 102424 400
rect 102592 0 102648 400
rect 102816 0 102872 400
rect 103040 0 103096 400
rect 103264 0 103320 400
rect 103488 0 103544 400
rect 103712 0 103768 400
rect 103936 0 103992 400
rect 104160 0 104216 400
rect 104384 0 104440 400
rect 104608 0 104664 400
rect 104832 0 104888 400
rect 105056 0 105112 400
rect 105280 0 105336 400
rect 105504 0 105560 400
rect 105728 0 105784 400
rect 105952 0 106008 400
rect 106176 0 106232 400
rect 106400 0 106456 400
rect 106624 0 106680 400
rect 106848 0 106904 400
rect 107072 0 107128 400
rect 107296 0 107352 400
rect 107520 0 107576 400
rect 107744 0 107800 400
rect 107968 0 108024 400
rect 108192 0 108248 400
rect 108416 0 108472 400
rect 108640 0 108696 400
rect 108864 0 108920 400
rect 109088 0 109144 400
rect 109312 0 109368 400
rect 109536 0 109592 400
rect 109760 0 109816 400
rect 109984 0 110040 400
rect 110208 0 110264 400
rect 110432 0 110488 400
rect 110656 0 110712 400
rect 110880 0 110936 400
rect 111104 0 111160 400
rect 111328 0 111384 400
<< obsm2 >>
rect 630 36570 2994 36666
rect 3110 36570 3890 36666
rect 4006 36570 4786 36666
rect 4902 36570 5682 36666
rect 5798 36570 6578 36666
rect 6694 36570 7474 36666
rect 7590 36570 8370 36666
rect 8486 36570 9266 36666
rect 9382 36570 10162 36666
rect 10278 36570 11058 36666
rect 11174 36570 11954 36666
rect 12070 36570 12850 36666
rect 12966 36570 13746 36666
rect 13862 36570 14642 36666
rect 14758 36570 15538 36666
rect 15654 36570 16434 36666
rect 16550 36570 17330 36666
rect 17446 36570 18226 36666
rect 18342 36570 19122 36666
rect 19238 36570 20018 36666
rect 20134 36570 20914 36666
rect 21030 36570 21810 36666
rect 21926 36570 22706 36666
rect 22822 36570 23602 36666
rect 23718 36570 24498 36666
rect 24614 36570 25394 36666
rect 25510 36570 26290 36666
rect 26406 36570 27186 36666
rect 27302 36570 28082 36666
rect 28198 36570 28978 36666
rect 29094 36570 29874 36666
rect 29990 36570 30770 36666
rect 30886 36570 31666 36666
rect 31782 36570 32562 36666
rect 32678 36570 33458 36666
rect 33574 36570 34354 36666
rect 34470 36570 35250 36666
rect 35366 36570 36146 36666
rect 36262 36570 37042 36666
rect 37158 36570 37938 36666
rect 38054 36570 38834 36666
rect 38950 36570 39730 36666
rect 39846 36570 40626 36666
rect 40742 36570 41522 36666
rect 41638 36570 42418 36666
rect 42534 36570 43314 36666
rect 43430 36570 44210 36666
rect 44326 36570 45106 36666
rect 45222 36570 46002 36666
rect 46118 36570 46898 36666
rect 47014 36570 47794 36666
rect 47910 36570 48690 36666
rect 48806 36570 49586 36666
rect 49702 36570 50482 36666
rect 50598 36570 51378 36666
rect 51494 36570 52274 36666
rect 52390 36570 53170 36666
rect 53286 36570 54066 36666
rect 54182 36570 54962 36666
rect 55078 36570 55858 36666
rect 55974 36570 56754 36666
rect 56870 36570 57650 36666
rect 57766 36570 58546 36666
rect 58662 36570 59442 36666
rect 59558 36570 60338 36666
rect 60454 36570 61234 36666
rect 61350 36570 62130 36666
rect 62246 36570 63026 36666
rect 63142 36570 63922 36666
rect 64038 36570 64818 36666
rect 64934 36570 65714 36666
rect 65830 36570 66610 36666
rect 66726 36570 67506 36666
rect 67622 36570 68402 36666
rect 68518 36570 69298 36666
rect 69414 36570 70194 36666
rect 70310 36570 71090 36666
rect 71206 36570 71986 36666
rect 72102 36570 72882 36666
rect 72998 36570 73778 36666
rect 73894 36570 74674 36666
rect 74790 36570 75570 36666
rect 75686 36570 76466 36666
rect 76582 36570 77362 36666
rect 77478 36570 78258 36666
rect 78374 36570 79154 36666
rect 79270 36570 80050 36666
rect 80166 36570 80946 36666
rect 81062 36570 81842 36666
rect 81958 36570 82738 36666
rect 82854 36570 83634 36666
rect 83750 36570 84530 36666
rect 84646 36570 85426 36666
rect 85542 36570 86322 36666
rect 86438 36570 87218 36666
rect 87334 36570 88114 36666
rect 88230 36570 89010 36666
rect 89126 36570 89906 36666
rect 90022 36570 90802 36666
rect 90918 36570 91698 36666
rect 91814 36570 92594 36666
rect 92710 36570 93490 36666
rect 93606 36570 94386 36666
rect 94502 36570 95282 36666
rect 95398 36570 96178 36666
rect 96294 36570 97074 36666
rect 97190 36570 97970 36666
rect 98086 36570 98866 36666
rect 98982 36570 99762 36666
rect 99878 36570 100658 36666
rect 100774 36570 101554 36666
rect 101670 36570 102450 36666
rect 102566 36570 103346 36666
rect 103462 36570 104242 36666
rect 104358 36570 105138 36666
rect 105254 36570 106034 36666
rect 106150 36570 106930 36666
rect 107046 36570 107826 36666
rect 107942 36570 108722 36666
rect 108838 36570 109618 36666
rect 109734 36570 110514 36666
rect 110630 36570 111410 36666
rect 111526 36570 112306 36666
rect 112422 36570 113202 36666
rect 113318 36570 114098 36666
rect 114214 36570 114994 36666
rect 115110 36570 115890 36666
rect 116006 36570 116786 36666
rect 116902 36570 119266 36666
rect 630 430 119266 36570
rect 630 289 8482 430
rect 8598 289 8706 430
rect 8822 289 8930 430
rect 9046 289 9154 430
rect 9270 289 9378 430
rect 9494 289 9602 430
rect 9718 289 9826 430
rect 9942 289 10050 430
rect 10166 289 10274 430
rect 10390 289 10498 430
rect 10614 289 10722 430
rect 10838 289 10946 430
rect 11062 289 11170 430
rect 11286 289 11394 430
rect 11510 289 11618 430
rect 11734 289 11842 430
rect 11958 289 12066 430
rect 12182 289 12290 430
rect 12406 289 12514 430
rect 12630 289 12738 430
rect 12854 289 12962 430
rect 13078 289 13186 430
rect 13302 289 13410 430
rect 13526 289 13634 430
rect 13750 289 13858 430
rect 13974 289 14082 430
rect 14198 289 14306 430
rect 14422 289 14530 430
rect 14646 289 14754 430
rect 14870 289 14978 430
rect 15094 289 15202 430
rect 15318 289 15426 430
rect 15542 289 15650 430
rect 15766 289 15874 430
rect 15990 289 16098 430
rect 16214 289 16322 430
rect 16438 289 16546 430
rect 16662 289 16770 430
rect 16886 289 16994 430
rect 17110 289 17218 430
rect 17334 289 17442 430
rect 17558 289 17666 430
rect 17782 289 17890 430
rect 18006 289 18114 430
rect 18230 289 18338 430
rect 18454 289 18562 430
rect 18678 289 18786 430
rect 18902 289 19010 430
rect 19126 289 19234 430
rect 19350 289 19458 430
rect 19574 289 19682 430
rect 19798 289 19906 430
rect 20022 289 20130 430
rect 20246 289 20354 430
rect 20470 289 20578 430
rect 20694 289 20802 430
rect 20918 289 21026 430
rect 21142 289 21250 430
rect 21366 289 21474 430
rect 21590 289 21698 430
rect 21814 289 21922 430
rect 22038 289 22146 430
rect 22262 289 22370 430
rect 22486 289 22594 430
rect 22710 289 22818 430
rect 22934 289 23042 430
rect 23158 289 23266 430
rect 23382 289 23490 430
rect 23606 289 23714 430
rect 23830 289 23938 430
rect 24054 289 24162 430
rect 24278 289 24386 430
rect 24502 289 24610 430
rect 24726 289 24834 430
rect 24950 289 25058 430
rect 25174 289 25282 430
rect 25398 289 25506 430
rect 25622 289 25730 430
rect 25846 289 25954 430
rect 26070 289 26178 430
rect 26294 289 26402 430
rect 26518 289 26626 430
rect 26742 289 26850 430
rect 26966 289 27074 430
rect 27190 289 27298 430
rect 27414 289 27522 430
rect 27638 289 27746 430
rect 27862 289 27970 430
rect 28086 289 28194 430
rect 28310 289 28418 430
rect 28534 289 28642 430
rect 28758 289 28866 430
rect 28982 289 29090 430
rect 29206 289 29314 430
rect 29430 289 29538 430
rect 29654 289 29762 430
rect 29878 289 29986 430
rect 30102 289 30210 430
rect 30326 289 30434 430
rect 30550 289 30658 430
rect 30774 289 30882 430
rect 30998 289 31106 430
rect 31222 289 31330 430
rect 31446 289 31554 430
rect 31670 289 31778 430
rect 31894 289 32002 430
rect 32118 289 32226 430
rect 32342 289 32450 430
rect 32566 289 32674 430
rect 32790 289 32898 430
rect 33014 289 33122 430
rect 33238 289 33346 430
rect 33462 289 33570 430
rect 33686 289 33794 430
rect 33910 289 34018 430
rect 34134 289 34242 430
rect 34358 289 34466 430
rect 34582 289 34690 430
rect 34806 289 34914 430
rect 35030 289 35138 430
rect 35254 289 35362 430
rect 35478 289 35586 430
rect 35702 289 35810 430
rect 35926 289 36034 430
rect 36150 289 36258 430
rect 36374 289 36482 430
rect 36598 289 36706 430
rect 36822 289 36930 430
rect 37046 289 37154 430
rect 37270 289 37378 430
rect 37494 289 37602 430
rect 37718 289 37826 430
rect 37942 289 38050 430
rect 38166 289 38274 430
rect 38390 289 38498 430
rect 38614 289 38722 430
rect 38838 289 38946 430
rect 39062 289 39170 430
rect 39286 289 39394 430
rect 39510 289 39618 430
rect 39734 289 39842 430
rect 39958 289 40066 430
rect 40182 289 40290 430
rect 40406 289 40514 430
rect 40630 289 40738 430
rect 40854 289 40962 430
rect 41078 289 41186 430
rect 41302 289 41410 430
rect 41526 289 41634 430
rect 41750 289 41858 430
rect 41974 289 42082 430
rect 42198 289 42306 430
rect 42422 289 42530 430
rect 42646 289 42754 430
rect 42870 289 42978 430
rect 43094 289 43202 430
rect 43318 289 43426 430
rect 43542 289 43650 430
rect 43766 289 43874 430
rect 43990 289 44098 430
rect 44214 289 44322 430
rect 44438 289 44546 430
rect 44662 289 44770 430
rect 44886 289 44994 430
rect 45110 289 45218 430
rect 45334 289 45442 430
rect 45558 289 45666 430
rect 45782 289 45890 430
rect 46006 289 46114 430
rect 46230 289 46338 430
rect 46454 289 46562 430
rect 46678 289 46786 430
rect 46902 289 47010 430
rect 47126 289 47234 430
rect 47350 289 47458 430
rect 47574 289 47682 430
rect 47798 289 47906 430
rect 48022 289 48130 430
rect 48246 289 48354 430
rect 48470 289 48578 430
rect 48694 289 48802 430
rect 48918 289 49026 430
rect 49142 289 49250 430
rect 49366 289 49474 430
rect 49590 289 49698 430
rect 49814 289 49922 430
rect 50038 289 50146 430
rect 50262 289 50370 430
rect 50486 289 50594 430
rect 50710 289 50818 430
rect 50934 289 51042 430
rect 51158 289 51266 430
rect 51382 289 51490 430
rect 51606 289 51714 430
rect 51830 289 51938 430
rect 52054 289 52162 430
rect 52278 289 52386 430
rect 52502 289 52610 430
rect 52726 289 52834 430
rect 52950 289 53058 430
rect 53174 289 53282 430
rect 53398 289 53506 430
rect 53622 289 53730 430
rect 53846 289 53954 430
rect 54070 289 54178 430
rect 54294 289 54402 430
rect 54518 289 54626 430
rect 54742 289 54850 430
rect 54966 289 55074 430
rect 55190 289 55298 430
rect 55414 289 55522 430
rect 55638 289 55746 430
rect 55862 289 55970 430
rect 56086 289 56194 430
rect 56310 289 56418 430
rect 56534 289 56642 430
rect 56758 289 56866 430
rect 56982 289 57090 430
rect 57206 289 57314 430
rect 57430 289 57538 430
rect 57654 289 57762 430
rect 57878 289 57986 430
rect 58102 289 58210 430
rect 58326 289 58434 430
rect 58550 289 58658 430
rect 58774 289 58882 430
rect 58998 289 59106 430
rect 59222 289 59330 430
rect 59446 289 59554 430
rect 59670 289 59778 430
rect 59894 289 60002 430
rect 60118 289 60226 430
rect 60342 289 60450 430
rect 60566 289 60674 430
rect 60790 289 60898 430
rect 61014 289 61122 430
rect 61238 289 61346 430
rect 61462 289 61570 430
rect 61686 289 61794 430
rect 61910 289 62018 430
rect 62134 289 62242 430
rect 62358 289 62466 430
rect 62582 289 62690 430
rect 62806 289 62914 430
rect 63030 289 63138 430
rect 63254 289 63362 430
rect 63478 289 63586 430
rect 63702 289 63810 430
rect 63926 289 64034 430
rect 64150 289 64258 430
rect 64374 289 64482 430
rect 64598 289 64706 430
rect 64822 289 64930 430
rect 65046 289 65154 430
rect 65270 289 65378 430
rect 65494 289 65602 430
rect 65718 289 65826 430
rect 65942 289 66050 430
rect 66166 289 66274 430
rect 66390 289 66498 430
rect 66614 289 66722 430
rect 66838 289 66946 430
rect 67062 289 67170 430
rect 67286 289 67394 430
rect 67510 289 67618 430
rect 67734 289 67842 430
rect 67958 289 68066 430
rect 68182 289 68290 430
rect 68406 289 68514 430
rect 68630 289 68738 430
rect 68854 289 68962 430
rect 69078 289 69186 430
rect 69302 289 69410 430
rect 69526 289 69634 430
rect 69750 289 69858 430
rect 69974 289 70082 430
rect 70198 289 70306 430
rect 70422 289 70530 430
rect 70646 289 70754 430
rect 70870 289 70978 430
rect 71094 289 71202 430
rect 71318 289 71426 430
rect 71542 289 71650 430
rect 71766 289 71874 430
rect 71990 289 72098 430
rect 72214 289 72322 430
rect 72438 289 72546 430
rect 72662 289 72770 430
rect 72886 289 72994 430
rect 73110 289 73218 430
rect 73334 289 73442 430
rect 73558 289 73666 430
rect 73782 289 73890 430
rect 74006 289 74114 430
rect 74230 289 74338 430
rect 74454 289 74562 430
rect 74678 289 74786 430
rect 74902 289 75010 430
rect 75126 289 75234 430
rect 75350 289 75458 430
rect 75574 289 75682 430
rect 75798 289 75906 430
rect 76022 289 76130 430
rect 76246 289 76354 430
rect 76470 289 76578 430
rect 76694 289 76802 430
rect 76918 289 77026 430
rect 77142 289 77250 430
rect 77366 289 77474 430
rect 77590 289 77698 430
rect 77814 289 77922 430
rect 78038 289 78146 430
rect 78262 289 78370 430
rect 78486 289 78594 430
rect 78710 289 78818 430
rect 78934 289 79042 430
rect 79158 289 79266 430
rect 79382 289 79490 430
rect 79606 289 79714 430
rect 79830 289 79938 430
rect 80054 289 80162 430
rect 80278 289 80386 430
rect 80502 289 80610 430
rect 80726 289 80834 430
rect 80950 289 81058 430
rect 81174 289 81282 430
rect 81398 289 81506 430
rect 81622 289 81730 430
rect 81846 289 81954 430
rect 82070 289 82178 430
rect 82294 289 82402 430
rect 82518 289 82626 430
rect 82742 289 82850 430
rect 82966 289 83074 430
rect 83190 289 83298 430
rect 83414 289 83522 430
rect 83638 289 83746 430
rect 83862 289 83970 430
rect 84086 289 84194 430
rect 84310 289 84418 430
rect 84534 289 84642 430
rect 84758 289 84866 430
rect 84982 289 85090 430
rect 85206 289 85314 430
rect 85430 289 85538 430
rect 85654 289 85762 430
rect 85878 289 85986 430
rect 86102 289 86210 430
rect 86326 289 86434 430
rect 86550 289 86658 430
rect 86774 289 86882 430
rect 86998 289 87106 430
rect 87222 289 87330 430
rect 87446 289 87554 430
rect 87670 289 87778 430
rect 87894 289 88002 430
rect 88118 289 88226 430
rect 88342 289 88450 430
rect 88566 289 88674 430
rect 88790 289 88898 430
rect 89014 289 89122 430
rect 89238 289 89346 430
rect 89462 289 89570 430
rect 89686 289 89794 430
rect 89910 289 90018 430
rect 90134 289 90242 430
rect 90358 289 90466 430
rect 90582 289 90690 430
rect 90806 289 90914 430
rect 91030 289 91138 430
rect 91254 289 91362 430
rect 91478 289 91586 430
rect 91702 289 91810 430
rect 91926 289 92034 430
rect 92150 289 92258 430
rect 92374 289 92482 430
rect 92598 289 92706 430
rect 92822 289 92930 430
rect 93046 289 93154 430
rect 93270 289 93378 430
rect 93494 289 93602 430
rect 93718 289 93826 430
rect 93942 289 94050 430
rect 94166 289 94274 430
rect 94390 289 94498 430
rect 94614 289 94722 430
rect 94838 289 94946 430
rect 95062 289 95170 430
rect 95286 289 95394 430
rect 95510 289 95618 430
rect 95734 289 95842 430
rect 95958 289 96066 430
rect 96182 289 96290 430
rect 96406 289 96514 430
rect 96630 289 96738 430
rect 96854 289 96962 430
rect 97078 289 97186 430
rect 97302 289 97410 430
rect 97526 289 97634 430
rect 97750 289 97858 430
rect 97974 289 98082 430
rect 98198 289 98306 430
rect 98422 289 98530 430
rect 98646 289 98754 430
rect 98870 289 98978 430
rect 99094 289 99202 430
rect 99318 289 99426 430
rect 99542 289 99650 430
rect 99766 289 99874 430
rect 99990 289 100098 430
rect 100214 289 100322 430
rect 100438 289 100546 430
rect 100662 289 100770 430
rect 100886 289 100994 430
rect 101110 289 101218 430
rect 101334 289 101442 430
rect 101558 289 101666 430
rect 101782 289 101890 430
rect 102006 289 102114 430
rect 102230 289 102338 430
rect 102454 289 102562 430
rect 102678 289 102786 430
rect 102902 289 103010 430
rect 103126 289 103234 430
rect 103350 289 103458 430
rect 103574 289 103682 430
rect 103798 289 103906 430
rect 104022 289 104130 430
rect 104246 289 104354 430
rect 104470 289 104578 430
rect 104694 289 104802 430
rect 104918 289 105026 430
rect 105142 289 105250 430
rect 105366 289 105474 430
rect 105590 289 105698 430
rect 105814 289 105922 430
rect 106038 289 106146 430
rect 106262 289 106370 430
rect 106486 289 106594 430
rect 106710 289 106818 430
rect 106934 289 107042 430
rect 107158 289 107266 430
rect 107382 289 107490 430
rect 107606 289 107714 430
rect 107830 289 107938 430
rect 108054 289 108162 430
rect 108278 289 108386 430
rect 108502 289 108610 430
rect 108726 289 108834 430
rect 108950 289 109058 430
rect 109174 289 109282 430
rect 109398 289 109506 430
rect 109622 289 109730 430
rect 109846 289 109954 430
rect 110070 289 110178 430
rect 110294 289 110402 430
rect 110518 289 110626 430
rect 110742 289 110850 430
rect 110966 289 111074 430
rect 111190 289 111298 430
rect 111414 289 119266 430
<< metal3 >>
rect 0 33712 400 33768
rect 119600 33712 120000 33768
rect 0 33376 400 33432
rect 119600 33376 120000 33432
rect 0 33040 400 33096
rect 119600 33040 120000 33096
rect 0 32704 400 32760
rect 119600 32704 120000 32760
rect 0 32368 400 32424
rect 119600 32368 120000 32424
rect 0 32032 400 32088
rect 119600 32032 120000 32088
rect 0 31696 400 31752
rect 119600 31696 120000 31752
rect 0 31360 400 31416
rect 119600 31360 120000 31416
rect 0 31024 400 31080
rect 119600 31024 120000 31080
rect 0 30688 400 30744
rect 119600 30688 120000 30744
rect 0 30352 400 30408
rect 119600 30352 120000 30408
rect 0 30016 400 30072
rect 119600 30016 120000 30072
rect 0 29680 400 29736
rect 119600 29680 120000 29736
rect 0 29344 400 29400
rect 119600 29344 120000 29400
rect 0 29008 400 29064
rect 119600 29008 120000 29064
rect 0 28672 400 28728
rect 119600 28672 120000 28728
rect 0 28336 400 28392
rect 119600 28336 120000 28392
rect 0 28000 400 28056
rect 119600 28000 120000 28056
rect 0 27664 400 27720
rect 119600 27664 120000 27720
rect 0 27328 400 27384
rect 119600 27328 120000 27384
rect 0 26992 400 27048
rect 119600 26992 120000 27048
rect 0 26656 400 26712
rect 119600 26656 120000 26712
rect 0 26320 400 26376
rect 119600 26320 120000 26376
rect 0 25984 400 26040
rect 119600 25984 120000 26040
rect 0 25648 400 25704
rect 119600 25648 120000 25704
rect 0 25312 400 25368
rect 119600 25312 120000 25368
rect 0 24976 400 25032
rect 119600 24976 120000 25032
rect 0 24640 400 24696
rect 119600 24640 120000 24696
rect 0 24304 400 24360
rect 119600 24304 120000 24360
rect 0 23968 400 24024
rect 119600 23968 120000 24024
rect 0 23632 400 23688
rect 119600 23632 120000 23688
rect 0 23296 400 23352
rect 119600 23296 120000 23352
rect 0 22960 400 23016
rect 119600 22960 120000 23016
rect 0 22624 400 22680
rect 119600 22624 120000 22680
rect 0 22288 400 22344
rect 119600 22288 120000 22344
rect 0 21952 400 22008
rect 119600 21952 120000 22008
rect 0 21616 400 21672
rect 119600 21616 120000 21672
rect 0 21280 400 21336
rect 119600 21280 120000 21336
rect 0 20944 400 21000
rect 119600 20944 120000 21000
rect 0 20608 400 20664
rect 119600 20608 120000 20664
rect 0 20272 400 20328
rect 119600 20272 120000 20328
rect 0 19936 400 19992
rect 119600 19936 120000 19992
rect 0 19600 400 19656
rect 119600 19600 120000 19656
rect 0 19264 400 19320
rect 119600 19264 120000 19320
rect 0 18928 400 18984
rect 119600 18928 120000 18984
rect 0 18592 400 18648
rect 119600 18592 120000 18648
rect 0 18256 400 18312
rect 119600 18256 120000 18312
rect 0 17920 400 17976
rect 119600 17920 120000 17976
rect 0 17584 400 17640
rect 119600 17584 120000 17640
rect 0 17248 400 17304
rect 119600 17248 120000 17304
rect 0 16912 400 16968
rect 119600 16912 120000 16968
rect 0 16576 400 16632
rect 119600 16576 120000 16632
rect 0 16240 400 16296
rect 119600 16240 120000 16296
rect 0 15904 400 15960
rect 119600 15904 120000 15960
rect 0 15568 400 15624
rect 119600 15568 120000 15624
rect 0 15232 400 15288
rect 119600 15232 120000 15288
rect 0 14896 400 14952
rect 119600 14896 120000 14952
rect 0 14560 400 14616
rect 119600 14560 120000 14616
rect 0 14224 400 14280
rect 119600 14224 120000 14280
rect 0 13888 400 13944
rect 119600 13888 120000 13944
rect 0 13552 400 13608
rect 119600 13552 120000 13608
rect 0 13216 400 13272
rect 119600 13216 120000 13272
rect 0 12880 400 12936
rect 119600 12880 120000 12936
rect 0 12544 400 12600
rect 119600 12544 120000 12600
rect 0 12208 400 12264
rect 119600 12208 120000 12264
rect 0 11872 400 11928
rect 119600 11872 120000 11928
rect 0 11536 400 11592
rect 119600 11536 120000 11592
rect 0 11200 400 11256
rect 119600 11200 120000 11256
rect 0 10864 400 10920
rect 119600 10864 120000 10920
rect 0 10528 400 10584
rect 119600 10528 120000 10584
rect 0 10192 400 10248
rect 119600 10192 120000 10248
rect 0 9856 400 9912
rect 119600 9856 120000 9912
rect 0 9520 400 9576
rect 119600 9520 120000 9576
rect 0 9184 400 9240
rect 119600 9184 120000 9240
rect 0 8848 400 8904
rect 119600 8848 120000 8904
rect 0 8512 400 8568
rect 119600 8512 120000 8568
rect 0 8176 400 8232
rect 119600 8176 120000 8232
rect 0 7840 400 7896
rect 119600 7840 120000 7896
rect 0 7504 400 7560
rect 119600 7504 120000 7560
rect 0 7168 400 7224
rect 119600 7168 120000 7224
rect 0 6832 400 6888
rect 119600 6832 120000 6888
rect 0 6496 400 6552
rect 119600 6496 120000 6552
rect 0 6160 400 6216
rect 119600 6160 120000 6216
rect 0 5824 400 5880
rect 119600 5824 120000 5880
rect 0 5488 400 5544
rect 119600 5488 120000 5544
rect 0 5152 400 5208
rect 119600 5152 120000 5208
rect 0 4816 400 4872
rect 119600 4816 120000 4872
rect 0 4480 400 4536
rect 119600 4480 120000 4536
rect 0 4144 400 4200
rect 119600 4144 120000 4200
rect 0 3808 400 3864
rect 119600 3808 120000 3864
rect 0 3472 400 3528
rect 119600 3472 120000 3528
rect 0 3136 400 3192
rect 119600 3136 120000 3192
<< obsm3 >>
rect 400 33798 119600 36498
rect 430 33682 119570 33798
rect 400 33462 119600 33682
rect 430 33346 119570 33462
rect 400 33126 119600 33346
rect 430 33010 119570 33126
rect 400 32790 119600 33010
rect 430 32674 119570 32790
rect 400 32454 119600 32674
rect 430 32338 119570 32454
rect 400 32118 119600 32338
rect 430 32002 119570 32118
rect 400 31782 119600 32002
rect 430 31666 119570 31782
rect 400 31446 119600 31666
rect 430 31330 119570 31446
rect 400 31110 119600 31330
rect 430 30994 119570 31110
rect 400 30774 119600 30994
rect 430 30658 119570 30774
rect 400 30438 119600 30658
rect 430 30322 119570 30438
rect 400 30102 119600 30322
rect 430 29986 119570 30102
rect 400 29766 119600 29986
rect 430 29650 119570 29766
rect 400 29430 119600 29650
rect 430 29314 119570 29430
rect 400 29094 119600 29314
rect 430 28978 119570 29094
rect 400 28758 119600 28978
rect 430 28642 119570 28758
rect 400 28422 119600 28642
rect 430 28306 119570 28422
rect 400 28086 119600 28306
rect 430 27970 119570 28086
rect 400 27750 119600 27970
rect 430 27634 119570 27750
rect 400 27414 119600 27634
rect 430 27298 119570 27414
rect 400 27078 119600 27298
rect 430 26962 119570 27078
rect 400 26742 119600 26962
rect 430 26626 119570 26742
rect 400 26406 119600 26626
rect 430 26290 119570 26406
rect 400 26070 119600 26290
rect 430 25954 119570 26070
rect 400 25734 119600 25954
rect 430 25618 119570 25734
rect 400 25398 119600 25618
rect 430 25282 119570 25398
rect 400 25062 119600 25282
rect 430 24946 119570 25062
rect 400 24726 119600 24946
rect 430 24610 119570 24726
rect 400 24390 119600 24610
rect 430 24274 119570 24390
rect 400 24054 119600 24274
rect 430 23938 119570 24054
rect 400 23718 119600 23938
rect 430 23602 119570 23718
rect 400 23382 119600 23602
rect 430 23266 119570 23382
rect 400 23046 119600 23266
rect 430 22930 119570 23046
rect 400 22710 119600 22930
rect 430 22594 119570 22710
rect 400 22374 119600 22594
rect 430 22258 119570 22374
rect 400 22038 119600 22258
rect 430 21922 119570 22038
rect 400 21702 119600 21922
rect 430 21586 119570 21702
rect 400 21366 119600 21586
rect 430 21250 119570 21366
rect 400 21030 119600 21250
rect 430 20914 119570 21030
rect 400 20694 119600 20914
rect 430 20578 119570 20694
rect 400 20358 119600 20578
rect 430 20242 119570 20358
rect 400 20022 119600 20242
rect 430 19906 119570 20022
rect 400 19686 119600 19906
rect 430 19570 119570 19686
rect 400 19350 119600 19570
rect 430 19234 119570 19350
rect 400 19014 119600 19234
rect 430 18898 119570 19014
rect 400 18678 119600 18898
rect 430 18562 119570 18678
rect 400 18342 119600 18562
rect 430 18226 119570 18342
rect 400 18006 119600 18226
rect 430 17890 119570 18006
rect 400 17670 119600 17890
rect 430 17554 119570 17670
rect 400 17334 119600 17554
rect 430 17218 119570 17334
rect 400 16998 119600 17218
rect 430 16882 119570 16998
rect 400 16662 119600 16882
rect 430 16546 119570 16662
rect 400 16326 119600 16546
rect 430 16210 119570 16326
rect 400 15990 119600 16210
rect 430 15874 119570 15990
rect 400 15654 119600 15874
rect 430 15538 119570 15654
rect 400 15318 119600 15538
rect 430 15202 119570 15318
rect 400 14982 119600 15202
rect 430 14866 119570 14982
rect 400 14646 119600 14866
rect 430 14530 119570 14646
rect 400 14310 119600 14530
rect 430 14194 119570 14310
rect 400 13974 119600 14194
rect 430 13858 119570 13974
rect 400 13638 119600 13858
rect 430 13522 119570 13638
rect 400 13302 119600 13522
rect 430 13186 119570 13302
rect 400 12966 119600 13186
rect 430 12850 119570 12966
rect 400 12630 119600 12850
rect 430 12514 119570 12630
rect 400 12294 119600 12514
rect 430 12178 119570 12294
rect 400 11958 119600 12178
rect 430 11842 119570 11958
rect 400 11622 119600 11842
rect 430 11506 119570 11622
rect 400 11286 119600 11506
rect 430 11170 119570 11286
rect 400 10950 119600 11170
rect 430 10834 119570 10950
rect 400 10614 119600 10834
rect 430 10498 119570 10614
rect 400 10278 119600 10498
rect 430 10162 119570 10278
rect 400 9942 119600 10162
rect 430 9826 119570 9942
rect 400 9606 119600 9826
rect 430 9490 119570 9606
rect 400 9270 119600 9490
rect 430 9154 119570 9270
rect 400 8934 119600 9154
rect 430 8818 119570 8934
rect 400 8598 119600 8818
rect 430 8482 119570 8598
rect 400 8262 119600 8482
rect 430 8146 119570 8262
rect 400 7926 119600 8146
rect 430 7810 119570 7926
rect 400 7590 119600 7810
rect 430 7474 119570 7590
rect 400 7254 119600 7474
rect 430 7138 119570 7254
rect 400 6918 119600 7138
rect 430 6802 119570 6918
rect 400 6582 119600 6802
rect 430 6466 119570 6582
rect 400 6246 119600 6466
rect 430 6130 119570 6246
rect 400 5910 119600 6130
rect 430 5794 119570 5910
rect 400 5574 119600 5794
rect 430 5458 119570 5574
rect 400 5238 119600 5458
rect 430 5122 119570 5238
rect 400 4902 119600 5122
rect 430 4786 119570 4902
rect 400 4566 119600 4786
rect 430 4450 119570 4566
rect 400 4230 119600 4450
rect 430 4114 119570 4230
rect 400 3894 119600 4114
rect 430 3778 119570 3894
rect 400 3558 119600 3778
rect 430 3442 119570 3558
rect 400 3222 119600 3442
rect 430 3106 119570 3222
rect 400 294 119600 3106
<< metal4 >>
rect 2224 1538 2384 35310
rect 9904 1538 10064 35310
rect 17584 1538 17744 35310
rect 25264 1538 25424 35310
rect 32944 1538 33104 35310
rect 40624 1538 40784 35310
rect 48304 1538 48464 35310
rect 55984 1538 56144 35310
rect 63664 1538 63824 35310
rect 71344 1538 71504 35310
rect 79024 1538 79184 35310
rect 86704 1538 86864 35310
rect 94384 1538 94544 35310
rect 102064 1538 102224 35310
rect 109744 1538 109904 35310
rect 117424 1538 117584 35310
<< obsm4 >>
rect 1022 35340 118930 36447
rect 1022 1508 2194 35340
rect 2414 1508 9874 35340
rect 10094 1508 17554 35340
rect 17774 1508 25234 35340
rect 25454 1508 32914 35340
rect 33134 1508 40594 35340
rect 40814 1508 48274 35340
rect 48494 1508 55954 35340
rect 56174 1508 63634 35340
rect 63854 1508 71314 35340
rect 71534 1508 78994 35340
rect 79214 1508 86674 35340
rect 86894 1508 94354 35340
rect 94574 1508 102034 35340
rect 102254 1508 109714 35340
rect 109934 1508 117394 35340
rect 117614 1508 118930 35340
rect 1022 289 118930 1508
<< labels >>
rlabel metal2 s 8512 0 8568 400 6 c0_disable
port 1 nsew signal output
rlabel metal2 s 12320 0 12376 400 6 c0_i_core_int_sreg[0]
port 2 nsew signal output
rlabel metal2 s 34272 0 34328 400 6 c0_i_core_int_sreg[10]
port 3 nsew signal output
rlabel metal2 s 36064 0 36120 400 6 c0_i_core_int_sreg[11]
port 4 nsew signal output
rlabel metal2 s 37856 0 37912 400 6 c0_i_core_int_sreg[12]
port 5 nsew signal output
rlabel metal2 s 39648 0 39704 400 6 c0_i_core_int_sreg[13]
port 6 nsew signal output
rlabel metal2 s 41440 0 41496 400 6 c0_i_core_int_sreg[14]
port 7 nsew signal output
rlabel metal2 s 43232 0 43288 400 6 c0_i_core_int_sreg[15]
port 8 nsew signal output
rlabel metal2 s 14784 0 14840 400 6 c0_i_core_int_sreg[1]
port 9 nsew signal output
rlabel metal2 s 17248 0 17304 400 6 c0_i_core_int_sreg[2]
port 10 nsew signal output
rlabel metal2 s 19488 0 19544 400 6 c0_i_core_int_sreg[3]
port 11 nsew signal output
rlabel metal2 s 21728 0 21784 400 6 c0_i_core_int_sreg[4]
port 12 nsew signal output
rlabel metal2 s 23968 0 24024 400 6 c0_i_core_int_sreg[5]
port 13 nsew signal output
rlabel metal2 s 26208 0 26264 400 6 c0_i_core_int_sreg[6]
port 14 nsew signal output
rlabel metal2 s 28448 0 28504 400 6 c0_i_core_int_sreg[7]
port 15 nsew signal output
rlabel metal2 s 30688 0 30744 400 6 c0_i_core_int_sreg[8]
port 16 nsew signal output
rlabel metal2 s 32480 0 32536 400 6 c0_i_core_int_sreg[9]
port 17 nsew signal output
rlabel metal2 s 8736 0 8792 400 6 c0_i_irq
port 18 nsew signal output
rlabel metal2 s 8960 0 9016 400 6 c0_i_mc_core_int
port 19 nsew signal output
rlabel metal2 s 9184 0 9240 400 6 c0_i_mem_ack
port 20 nsew signal output
rlabel metal2 s 12544 0 12600 400 6 c0_i_mem_data[0]
port 21 nsew signal output
rlabel metal2 s 34496 0 34552 400 6 c0_i_mem_data[10]
port 22 nsew signal output
rlabel metal2 s 36288 0 36344 400 6 c0_i_mem_data[11]
port 23 nsew signal output
rlabel metal2 s 38080 0 38136 400 6 c0_i_mem_data[12]
port 24 nsew signal output
rlabel metal2 s 39872 0 39928 400 6 c0_i_mem_data[13]
port 25 nsew signal output
rlabel metal2 s 41664 0 41720 400 6 c0_i_mem_data[14]
port 26 nsew signal output
rlabel metal2 s 43456 0 43512 400 6 c0_i_mem_data[15]
port 27 nsew signal output
rlabel metal2 s 15008 0 15064 400 6 c0_i_mem_data[1]
port 28 nsew signal output
rlabel metal2 s 17472 0 17528 400 6 c0_i_mem_data[2]
port 29 nsew signal output
rlabel metal2 s 19712 0 19768 400 6 c0_i_mem_data[3]
port 30 nsew signal output
rlabel metal2 s 21952 0 22008 400 6 c0_i_mem_data[4]
port 31 nsew signal output
rlabel metal2 s 24192 0 24248 400 6 c0_i_mem_data[5]
port 32 nsew signal output
rlabel metal2 s 26432 0 26488 400 6 c0_i_mem_data[6]
port 33 nsew signal output
rlabel metal2 s 28672 0 28728 400 6 c0_i_mem_data[7]
port 34 nsew signal output
rlabel metal2 s 30912 0 30968 400 6 c0_i_mem_data[8]
port 35 nsew signal output
rlabel metal2 s 32704 0 32760 400 6 c0_i_mem_data[9]
port 36 nsew signal output
rlabel metal2 s 9408 0 9464 400 6 c0_i_mem_exception
port 37 nsew signal output
rlabel metal2 s 12768 0 12824 400 6 c0_i_req_data[0]
port 38 nsew signal output
rlabel metal2 s 34720 0 34776 400 6 c0_i_req_data[10]
port 39 nsew signal output
rlabel metal2 s 36512 0 36568 400 6 c0_i_req_data[11]
port 40 nsew signal output
rlabel metal2 s 38304 0 38360 400 6 c0_i_req_data[12]
port 41 nsew signal output
rlabel metal2 s 40096 0 40152 400 6 c0_i_req_data[13]
port 42 nsew signal output
rlabel metal2 s 41888 0 41944 400 6 c0_i_req_data[14]
port 43 nsew signal output
rlabel metal2 s 43680 0 43736 400 6 c0_i_req_data[15]
port 44 nsew signal output
rlabel metal2 s 45024 0 45080 400 6 c0_i_req_data[16]
port 45 nsew signal output
rlabel metal2 s 45248 0 45304 400 6 c0_i_req_data[17]
port 46 nsew signal output
rlabel metal2 s 45472 0 45528 400 6 c0_i_req_data[18]
port 47 nsew signal output
rlabel metal2 s 45696 0 45752 400 6 c0_i_req_data[19]
port 48 nsew signal output
rlabel metal2 s 15232 0 15288 400 6 c0_i_req_data[1]
port 49 nsew signal output
rlabel metal2 s 45920 0 45976 400 6 c0_i_req_data[20]
port 50 nsew signal output
rlabel metal2 s 46144 0 46200 400 6 c0_i_req_data[21]
port 51 nsew signal output
rlabel metal2 s 46368 0 46424 400 6 c0_i_req_data[22]
port 52 nsew signal output
rlabel metal2 s 46592 0 46648 400 6 c0_i_req_data[23]
port 53 nsew signal output
rlabel metal2 s 46816 0 46872 400 6 c0_i_req_data[24]
port 54 nsew signal output
rlabel metal2 s 47040 0 47096 400 6 c0_i_req_data[25]
port 55 nsew signal output
rlabel metal2 s 47264 0 47320 400 6 c0_i_req_data[26]
port 56 nsew signal output
rlabel metal2 s 47488 0 47544 400 6 c0_i_req_data[27]
port 57 nsew signal output
rlabel metal2 s 47712 0 47768 400 6 c0_i_req_data[28]
port 58 nsew signal output
rlabel metal2 s 47936 0 47992 400 6 c0_i_req_data[29]
port 59 nsew signal output
rlabel metal2 s 17696 0 17752 400 6 c0_i_req_data[2]
port 60 nsew signal output
rlabel metal2 s 48160 0 48216 400 6 c0_i_req_data[30]
port 61 nsew signal output
rlabel metal2 s 48384 0 48440 400 6 c0_i_req_data[31]
port 62 nsew signal output
rlabel metal2 s 19936 0 19992 400 6 c0_i_req_data[3]
port 63 nsew signal output
rlabel metal2 s 22176 0 22232 400 6 c0_i_req_data[4]
port 64 nsew signal output
rlabel metal2 s 24416 0 24472 400 6 c0_i_req_data[5]
port 65 nsew signal output
rlabel metal2 s 26656 0 26712 400 6 c0_i_req_data[6]
port 66 nsew signal output
rlabel metal2 s 28896 0 28952 400 6 c0_i_req_data[7]
port 67 nsew signal output
rlabel metal2 s 31136 0 31192 400 6 c0_i_req_data[8]
port 68 nsew signal output
rlabel metal2 s 32928 0 32984 400 6 c0_i_req_data[9]
port 69 nsew signal output
rlabel metal2 s 9632 0 9688 400 6 c0_i_req_data_valid
port 70 nsew signal output
rlabel metal2 s 9856 0 9912 400 6 c0_o_c_data_page
port 71 nsew signal input
rlabel metal2 s 10080 0 10136 400 6 c0_o_c_instr_long
port 72 nsew signal input
rlabel metal2 s 10304 0 10360 400 6 c0_o_c_instr_page
port 73 nsew signal input
rlabel metal2 s 10528 0 10584 400 6 c0_o_icache_flush
port 74 nsew signal input
rlabel metal2 s 12992 0 13048 400 6 c0_o_instr_long_addr[0]
port 75 nsew signal input
rlabel metal2 s 15456 0 15512 400 6 c0_o_instr_long_addr[1]
port 76 nsew signal input
rlabel metal2 s 17920 0 17976 400 6 c0_o_instr_long_addr[2]
port 77 nsew signal input
rlabel metal2 s 20160 0 20216 400 6 c0_o_instr_long_addr[3]
port 78 nsew signal input
rlabel metal2 s 22400 0 22456 400 6 c0_o_instr_long_addr[4]
port 79 nsew signal input
rlabel metal2 s 24640 0 24696 400 6 c0_o_instr_long_addr[5]
port 80 nsew signal input
rlabel metal2 s 26880 0 26936 400 6 c0_o_instr_long_addr[6]
port 81 nsew signal input
rlabel metal2 s 29120 0 29176 400 6 c0_o_instr_long_addr[7]
port 82 nsew signal input
rlabel metal2 s 13216 0 13272 400 6 c0_o_mem_addr[0]
port 83 nsew signal input
rlabel metal2 s 34944 0 35000 400 6 c0_o_mem_addr[10]
port 84 nsew signal input
rlabel metal2 s 36736 0 36792 400 6 c0_o_mem_addr[11]
port 85 nsew signal input
rlabel metal2 s 38528 0 38584 400 6 c0_o_mem_addr[12]
port 86 nsew signal input
rlabel metal2 s 40320 0 40376 400 6 c0_o_mem_addr[13]
port 87 nsew signal input
rlabel metal2 s 42112 0 42168 400 6 c0_o_mem_addr[14]
port 88 nsew signal input
rlabel metal2 s 43904 0 43960 400 6 c0_o_mem_addr[15]
port 89 nsew signal input
rlabel metal2 s 15680 0 15736 400 6 c0_o_mem_addr[1]
port 90 nsew signal input
rlabel metal2 s 18144 0 18200 400 6 c0_o_mem_addr[2]
port 91 nsew signal input
rlabel metal2 s 20384 0 20440 400 6 c0_o_mem_addr[3]
port 92 nsew signal input
rlabel metal2 s 22624 0 22680 400 6 c0_o_mem_addr[4]
port 93 nsew signal input
rlabel metal2 s 24864 0 24920 400 6 c0_o_mem_addr[5]
port 94 nsew signal input
rlabel metal2 s 27104 0 27160 400 6 c0_o_mem_addr[6]
port 95 nsew signal input
rlabel metal2 s 29344 0 29400 400 6 c0_o_mem_addr[7]
port 96 nsew signal input
rlabel metal2 s 31360 0 31416 400 6 c0_o_mem_addr[8]
port 97 nsew signal input
rlabel metal2 s 33152 0 33208 400 6 c0_o_mem_addr[9]
port 98 nsew signal input
rlabel metal2 s 13440 0 13496 400 6 c0_o_mem_data[0]
port 99 nsew signal input
rlabel metal2 s 35168 0 35224 400 6 c0_o_mem_data[10]
port 100 nsew signal input
rlabel metal2 s 36960 0 37016 400 6 c0_o_mem_data[11]
port 101 nsew signal input
rlabel metal2 s 38752 0 38808 400 6 c0_o_mem_data[12]
port 102 nsew signal input
rlabel metal2 s 40544 0 40600 400 6 c0_o_mem_data[13]
port 103 nsew signal input
rlabel metal2 s 42336 0 42392 400 6 c0_o_mem_data[14]
port 104 nsew signal input
rlabel metal2 s 44128 0 44184 400 6 c0_o_mem_data[15]
port 105 nsew signal input
rlabel metal2 s 15904 0 15960 400 6 c0_o_mem_data[1]
port 106 nsew signal input
rlabel metal2 s 18368 0 18424 400 6 c0_o_mem_data[2]
port 107 nsew signal input
rlabel metal2 s 20608 0 20664 400 6 c0_o_mem_data[3]
port 108 nsew signal input
rlabel metal2 s 22848 0 22904 400 6 c0_o_mem_data[4]
port 109 nsew signal input
rlabel metal2 s 25088 0 25144 400 6 c0_o_mem_data[5]
port 110 nsew signal input
rlabel metal2 s 27328 0 27384 400 6 c0_o_mem_data[6]
port 111 nsew signal input
rlabel metal2 s 29568 0 29624 400 6 c0_o_mem_data[7]
port 112 nsew signal input
rlabel metal2 s 31584 0 31640 400 6 c0_o_mem_data[8]
port 113 nsew signal input
rlabel metal2 s 33376 0 33432 400 6 c0_o_mem_data[9]
port 114 nsew signal input
rlabel metal2 s 13664 0 13720 400 6 c0_o_mem_high_addr[0]
port 115 nsew signal input
rlabel metal2 s 16128 0 16184 400 6 c0_o_mem_high_addr[1]
port 116 nsew signal input
rlabel metal2 s 18592 0 18648 400 6 c0_o_mem_high_addr[2]
port 117 nsew signal input
rlabel metal2 s 20832 0 20888 400 6 c0_o_mem_high_addr[3]
port 118 nsew signal input
rlabel metal2 s 23072 0 23128 400 6 c0_o_mem_high_addr[4]
port 119 nsew signal input
rlabel metal2 s 25312 0 25368 400 6 c0_o_mem_high_addr[5]
port 120 nsew signal input
rlabel metal2 s 27552 0 27608 400 6 c0_o_mem_high_addr[6]
port 121 nsew signal input
rlabel metal2 s 29792 0 29848 400 6 c0_o_mem_high_addr[7]
port 122 nsew signal input
rlabel metal2 s 10752 0 10808 400 6 c0_o_mem_long_mode
port 123 nsew signal input
rlabel metal2 s 10976 0 11032 400 6 c0_o_mem_req
port 124 nsew signal input
rlabel metal2 s 13888 0 13944 400 6 c0_o_mem_sel[0]
port 125 nsew signal input
rlabel metal2 s 16352 0 16408 400 6 c0_o_mem_sel[1]
port 126 nsew signal input
rlabel metal2 s 11200 0 11256 400 6 c0_o_mem_we
port 127 nsew signal input
rlabel metal2 s 11424 0 11480 400 6 c0_o_req_active
port 128 nsew signal input
rlabel metal2 s 14112 0 14168 400 6 c0_o_req_addr[0]
port 129 nsew signal input
rlabel metal2 s 35392 0 35448 400 6 c0_o_req_addr[10]
port 130 nsew signal input
rlabel metal2 s 37184 0 37240 400 6 c0_o_req_addr[11]
port 131 nsew signal input
rlabel metal2 s 38976 0 39032 400 6 c0_o_req_addr[12]
port 132 nsew signal input
rlabel metal2 s 40768 0 40824 400 6 c0_o_req_addr[13]
port 133 nsew signal input
rlabel metal2 s 42560 0 42616 400 6 c0_o_req_addr[14]
port 134 nsew signal input
rlabel metal2 s 44352 0 44408 400 6 c0_o_req_addr[15]
port 135 nsew signal input
rlabel metal2 s 16576 0 16632 400 6 c0_o_req_addr[1]
port 136 nsew signal input
rlabel metal2 s 18816 0 18872 400 6 c0_o_req_addr[2]
port 137 nsew signal input
rlabel metal2 s 21056 0 21112 400 6 c0_o_req_addr[3]
port 138 nsew signal input
rlabel metal2 s 23296 0 23352 400 6 c0_o_req_addr[4]
port 139 nsew signal input
rlabel metal2 s 25536 0 25592 400 6 c0_o_req_addr[5]
port 140 nsew signal input
rlabel metal2 s 27776 0 27832 400 6 c0_o_req_addr[6]
port 141 nsew signal input
rlabel metal2 s 30016 0 30072 400 6 c0_o_req_addr[7]
port 142 nsew signal input
rlabel metal2 s 31808 0 31864 400 6 c0_o_req_addr[8]
port 143 nsew signal input
rlabel metal2 s 33600 0 33656 400 6 c0_o_req_addr[9]
port 144 nsew signal input
rlabel metal2 s 11648 0 11704 400 6 c0_o_req_ppl_submit
port 145 nsew signal input
rlabel metal2 s 11872 0 11928 400 6 c0_rst
port 146 nsew signal output
rlabel metal2 s 14336 0 14392 400 6 c0_sr_bus_addr[0]
port 147 nsew signal input
rlabel metal2 s 35616 0 35672 400 6 c0_sr_bus_addr[10]
port 148 nsew signal input
rlabel metal2 s 37408 0 37464 400 6 c0_sr_bus_addr[11]
port 149 nsew signal input
rlabel metal2 s 39200 0 39256 400 6 c0_sr_bus_addr[12]
port 150 nsew signal input
rlabel metal2 s 40992 0 41048 400 6 c0_sr_bus_addr[13]
port 151 nsew signal input
rlabel metal2 s 42784 0 42840 400 6 c0_sr_bus_addr[14]
port 152 nsew signal input
rlabel metal2 s 44576 0 44632 400 6 c0_sr_bus_addr[15]
port 153 nsew signal input
rlabel metal2 s 16800 0 16856 400 6 c0_sr_bus_addr[1]
port 154 nsew signal input
rlabel metal2 s 19040 0 19096 400 6 c0_sr_bus_addr[2]
port 155 nsew signal input
rlabel metal2 s 21280 0 21336 400 6 c0_sr_bus_addr[3]
port 156 nsew signal input
rlabel metal2 s 23520 0 23576 400 6 c0_sr_bus_addr[4]
port 157 nsew signal input
rlabel metal2 s 25760 0 25816 400 6 c0_sr_bus_addr[5]
port 158 nsew signal input
rlabel metal2 s 28000 0 28056 400 6 c0_sr_bus_addr[6]
port 159 nsew signal input
rlabel metal2 s 30240 0 30296 400 6 c0_sr_bus_addr[7]
port 160 nsew signal input
rlabel metal2 s 32032 0 32088 400 6 c0_sr_bus_addr[8]
port 161 nsew signal input
rlabel metal2 s 33824 0 33880 400 6 c0_sr_bus_addr[9]
port 162 nsew signal input
rlabel metal2 s 14560 0 14616 400 6 c0_sr_bus_data_o[0]
port 163 nsew signal input
rlabel metal2 s 35840 0 35896 400 6 c0_sr_bus_data_o[10]
port 164 nsew signal input
rlabel metal2 s 37632 0 37688 400 6 c0_sr_bus_data_o[11]
port 165 nsew signal input
rlabel metal2 s 39424 0 39480 400 6 c0_sr_bus_data_o[12]
port 166 nsew signal input
rlabel metal2 s 41216 0 41272 400 6 c0_sr_bus_data_o[13]
port 167 nsew signal input
rlabel metal2 s 43008 0 43064 400 6 c0_sr_bus_data_o[14]
port 168 nsew signal input
rlabel metal2 s 44800 0 44856 400 6 c0_sr_bus_data_o[15]
port 169 nsew signal input
rlabel metal2 s 17024 0 17080 400 6 c0_sr_bus_data_o[1]
port 170 nsew signal input
rlabel metal2 s 19264 0 19320 400 6 c0_sr_bus_data_o[2]
port 171 nsew signal input
rlabel metal2 s 21504 0 21560 400 6 c0_sr_bus_data_o[3]
port 172 nsew signal input
rlabel metal2 s 23744 0 23800 400 6 c0_sr_bus_data_o[4]
port 173 nsew signal input
rlabel metal2 s 25984 0 26040 400 6 c0_sr_bus_data_o[5]
port 174 nsew signal input
rlabel metal2 s 28224 0 28280 400 6 c0_sr_bus_data_o[6]
port 175 nsew signal input
rlabel metal2 s 30464 0 30520 400 6 c0_sr_bus_data_o[7]
port 176 nsew signal input
rlabel metal2 s 32256 0 32312 400 6 c0_sr_bus_data_o[8]
port 177 nsew signal input
rlabel metal2 s 34048 0 34104 400 6 c0_sr_bus_data_o[9]
port 178 nsew signal input
rlabel metal2 s 12096 0 12152 400 6 c0_sr_bus_we
port 179 nsew signal input
rlabel metal2 s 68096 0 68152 400 6 c1_dbg_pc[0]
port 180 nsew signal input
rlabel metal2 s 94528 0 94584 400 6 c1_dbg_pc[10]
port 181 nsew signal input
rlabel metal2 s 96768 0 96824 400 6 c1_dbg_pc[11]
port 182 nsew signal input
rlabel metal2 s 99008 0 99064 400 6 c1_dbg_pc[12]
port 183 nsew signal input
rlabel metal2 s 101248 0 101304 400 6 c1_dbg_pc[13]
port 184 nsew signal input
rlabel metal2 s 103488 0 103544 400 6 c1_dbg_pc[14]
port 185 nsew signal input
rlabel metal2 s 105728 0 105784 400 6 c1_dbg_pc[15]
port 186 nsew signal input
rlabel metal2 s 71008 0 71064 400 6 c1_dbg_pc[1]
port 187 nsew signal input
rlabel metal2 s 73920 0 73976 400 6 c1_dbg_pc[2]
port 188 nsew signal input
rlabel metal2 s 76608 0 76664 400 6 c1_dbg_pc[3]
port 189 nsew signal input
rlabel metal2 s 79296 0 79352 400 6 c1_dbg_pc[4]
port 190 nsew signal input
rlabel metal2 s 81984 0 82040 400 6 c1_dbg_pc[5]
port 191 nsew signal input
rlabel metal2 s 84672 0 84728 400 6 c1_dbg_pc[6]
port 192 nsew signal input
rlabel metal2 s 87360 0 87416 400 6 c1_dbg_pc[7]
port 193 nsew signal input
rlabel metal2 s 90048 0 90104 400 6 c1_dbg_pc[8]
port 194 nsew signal input
rlabel metal2 s 92288 0 92344 400 6 c1_dbg_pc[9]
port 195 nsew signal input
rlabel metal2 s 68320 0 68376 400 6 c1_dbg_r0[0]
port 196 nsew signal input
rlabel metal2 s 94752 0 94808 400 6 c1_dbg_r0[10]
port 197 nsew signal input
rlabel metal2 s 96992 0 97048 400 6 c1_dbg_r0[11]
port 198 nsew signal input
rlabel metal2 s 99232 0 99288 400 6 c1_dbg_r0[12]
port 199 nsew signal input
rlabel metal2 s 101472 0 101528 400 6 c1_dbg_r0[13]
port 200 nsew signal input
rlabel metal2 s 103712 0 103768 400 6 c1_dbg_r0[14]
port 201 nsew signal input
rlabel metal2 s 105952 0 106008 400 6 c1_dbg_r0[15]
port 202 nsew signal input
rlabel metal2 s 71232 0 71288 400 6 c1_dbg_r0[1]
port 203 nsew signal input
rlabel metal2 s 74144 0 74200 400 6 c1_dbg_r0[2]
port 204 nsew signal input
rlabel metal2 s 76832 0 76888 400 6 c1_dbg_r0[3]
port 205 nsew signal input
rlabel metal2 s 79520 0 79576 400 6 c1_dbg_r0[4]
port 206 nsew signal input
rlabel metal2 s 82208 0 82264 400 6 c1_dbg_r0[5]
port 207 nsew signal input
rlabel metal2 s 84896 0 84952 400 6 c1_dbg_r0[6]
port 208 nsew signal input
rlabel metal2 s 87584 0 87640 400 6 c1_dbg_r0[7]
port 209 nsew signal input
rlabel metal2 s 90272 0 90328 400 6 c1_dbg_r0[8]
port 210 nsew signal input
rlabel metal2 s 92512 0 92568 400 6 c1_dbg_r0[9]
port 211 nsew signal input
rlabel metal2 s 64288 0 64344 400 6 c1_disable
port 212 nsew signal output
rlabel metal2 s 68544 0 68600 400 6 c1_i_core_int_sreg[0]
port 213 nsew signal output
rlabel metal2 s 94976 0 95032 400 6 c1_i_core_int_sreg[10]
port 214 nsew signal output
rlabel metal2 s 97216 0 97272 400 6 c1_i_core_int_sreg[11]
port 215 nsew signal output
rlabel metal2 s 99456 0 99512 400 6 c1_i_core_int_sreg[12]
port 216 nsew signal output
rlabel metal2 s 101696 0 101752 400 6 c1_i_core_int_sreg[13]
port 217 nsew signal output
rlabel metal2 s 103936 0 103992 400 6 c1_i_core_int_sreg[14]
port 218 nsew signal output
rlabel metal2 s 106176 0 106232 400 6 c1_i_core_int_sreg[15]
port 219 nsew signal output
rlabel metal2 s 71456 0 71512 400 6 c1_i_core_int_sreg[1]
port 220 nsew signal output
rlabel metal2 s 74368 0 74424 400 6 c1_i_core_int_sreg[2]
port 221 nsew signal output
rlabel metal2 s 77056 0 77112 400 6 c1_i_core_int_sreg[3]
port 222 nsew signal output
rlabel metal2 s 79744 0 79800 400 6 c1_i_core_int_sreg[4]
port 223 nsew signal output
rlabel metal2 s 82432 0 82488 400 6 c1_i_core_int_sreg[5]
port 224 nsew signal output
rlabel metal2 s 85120 0 85176 400 6 c1_i_core_int_sreg[6]
port 225 nsew signal output
rlabel metal2 s 87808 0 87864 400 6 c1_i_core_int_sreg[7]
port 226 nsew signal output
rlabel metal2 s 90496 0 90552 400 6 c1_i_core_int_sreg[8]
port 227 nsew signal output
rlabel metal2 s 92736 0 92792 400 6 c1_i_core_int_sreg[9]
port 228 nsew signal output
rlabel metal2 s 64512 0 64568 400 6 c1_i_irq
port 229 nsew signal output
rlabel metal2 s 64736 0 64792 400 6 c1_i_mc_core_int
port 230 nsew signal output
rlabel metal2 s 64960 0 65016 400 6 c1_i_mem_ack
port 231 nsew signal output
rlabel metal2 s 68768 0 68824 400 6 c1_i_mem_data[0]
port 232 nsew signal output
rlabel metal2 s 95200 0 95256 400 6 c1_i_mem_data[10]
port 233 nsew signal output
rlabel metal2 s 97440 0 97496 400 6 c1_i_mem_data[11]
port 234 nsew signal output
rlabel metal2 s 99680 0 99736 400 6 c1_i_mem_data[12]
port 235 nsew signal output
rlabel metal2 s 101920 0 101976 400 6 c1_i_mem_data[13]
port 236 nsew signal output
rlabel metal2 s 104160 0 104216 400 6 c1_i_mem_data[14]
port 237 nsew signal output
rlabel metal2 s 106400 0 106456 400 6 c1_i_mem_data[15]
port 238 nsew signal output
rlabel metal2 s 71680 0 71736 400 6 c1_i_mem_data[1]
port 239 nsew signal output
rlabel metal2 s 74592 0 74648 400 6 c1_i_mem_data[2]
port 240 nsew signal output
rlabel metal2 s 77280 0 77336 400 6 c1_i_mem_data[3]
port 241 nsew signal output
rlabel metal2 s 79968 0 80024 400 6 c1_i_mem_data[4]
port 242 nsew signal output
rlabel metal2 s 82656 0 82712 400 6 c1_i_mem_data[5]
port 243 nsew signal output
rlabel metal2 s 85344 0 85400 400 6 c1_i_mem_data[6]
port 244 nsew signal output
rlabel metal2 s 88032 0 88088 400 6 c1_i_mem_data[7]
port 245 nsew signal output
rlabel metal2 s 90720 0 90776 400 6 c1_i_mem_data[8]
port 246 nsew signal output
rlabel metal2 s 92960 0 93016 400 6 c1_i_mem_data[9]
port 247 nsew signal output
rlabel metal2 s 65184 0 65240 400 6 c1_i_mem_exception
port 248 nsew signal output
rlabel metal2 s 68992 0 69048 400 6 c1_i_req_data[0]
port 249 nsew signal output
rlabel metal2 s 95424 0 95480 400 6 c1_i_req_data[10]
port 250 nsew signal output
rlabel metal2 s 97664 0 97720 400 6 c1_i_req_data[11]
port 251 nsew signal output
rlabel metal2 s 99904 0 99960 400 6 c1_i_req_data[12]
port 252 nsew signal output
rlabel metal2 s 102144 0 102200 400 6 c1_i_req_data[13]
port 253 nsew signal output
rlabel metal2 s 104384 0 104440 400 6 c1_i_req_data[14]
port 254 nsew signal output
rlabel metal2 s 106624 0 106680 400 6 c1_i_req_data[15]
port 255 nsew signal output
rlabel metal2 s 107968 0 108024 400 6 c1_i_req_data[16]
port 256 nsew signal output
rlabel metal2 s 108192 0 108248 400 6 c1_i_req_data[17]
port 257 nsew signal output
rlabel metal2 s 108416 0 108472 400 6 c1_i_req_data[18]
port 258 nsew signal output
rlabel metal2 s 108640 0 108696 400 6 c1_i_req_data[19]
port 259 nsew signal output
rlabel metal2 s 71904 0 71960 400 6 c1_i_req_data[1]
port 260 nsew signal output
rlabel metal2 s 108864 0 108920 400 6 c1_i_req_data[20]
port 261 nsew signal output
rlabel metal2 s 109088 0 109144 400 6 c1_i_req_data[21]
port 262 nsew signal output
rlabel metal2 s 109312 0 109368 400 6 c1_i_req_data[22]
port 263 nsew signal output
rlabel metal2 s 109536 0 109592 400 6 c1_i_req_data[23]
port 264 nsew signal output
rlabel metal2 s 109760 0 109816 400 6 c1_i_req_data[24]
port 265 nsew signal output
rlabel metal2 s 109984 0 110040 400 6 c1_i_req_data[25]
port 266 nsew signal output
rlabel metal2 s 110208 0 110264 400 6 c1_i_req_data[26]
port 267 nsew signal output
rlabel metal2 s 110432 0 110488 400 6 c1_i_req_data[27]
port 268 nsew signal output
rlabel metal2 s 110656 0 110712 400 6 c1_i_req_data[28]
port 269 nsew signal output
rlabel metal2 s 110880 0 110936 400 6 c1_i_req_data[29]
port 270 nsew signal output
rlabel metal2 s 74816 0 74872 400 6 c1_i_req_data[2]
port 271 nsew signal output
rlabel metal2 s 111104 0 111160 400 6 c1_i_req_data[30]
port 272 nsew signal output
rlabel metal2 s 111328 0 111384 400 6 c1_i_req_data[31]
port 273 nsew signal output
rlabel metal2 s 77504 0 77560 400 6 c1_i_req_data[3]
port 274 nsew signal output
rlabel metal2 s 80192 0 80248 400 6 c1_i_req_data[4]
port 275 nsew signal output
rlabel metal2 s 82880 0 82936 400 6 c1_i_req_data[5]
port 276 nsew signal output
rlabel metal2 s 85568 0 85624 400 6 c1_i_req_data[6]
port 277 nsew signal output
rlabel metal2 s 88256 0 88312 400 6 c1_i_req_data[7]
port 278 nsew signal output
rlabel metal2 s 90944 0 91000 400 6 c1_i_req_data[8]
port 279 nsew signal output
rlabel metal2 s 93184 0 93240 400 6 c1_i_req_data[9]
port 280 nsew signal output
rlabel metal2 s 65408 0 65464 400 6 c1_i_req_data_valid
port 281 nsew signal output
rlabel metal2 s 65632 0 65688 400 6 c1_o_c_data_page
port 282 nsew signal input
rlabel metal2 s 65856 0 65912 400 6 c1_o_c_instr_long
port 283 nsew signal input
rlabel metal2 s 66080 0 66136 400 6 c1_o_c_instr_page
port 284 nsew signal input
rlabel metal2 s 66304 0 66360 400 6 c1_o_icache_flush
port 285 nsew signal input
rlabel metal2 s 69216 0 69272 400 6 c1_o_instr_long_addr[0]
port 286 nsew signal input
rlabel metal2 s 72128 0 72184 400 6 c1_o_instr_long_addr[1]
port 287 nsew signal input
rlabel metal2 s 75040 0 75096 400 6 c1_o_instr_long_addr[2]
port 288 nsew signal input
rlabel metal2 s 77728 0 77784 400 6 c1_o_instr_long_addr[3]
port 289 nsew signal input
rlabel metal2 s 80416 0 80472 400 6 c1_o_instr_long_addr[4]
port 290 nsew signal input
rlabel metal2 s 83104 0 83160 400 6 c1_o_instr_long_addr[5]
port 291 nsew signal input
rlabel metal2 s 85792 0 85848 400 6 c1_o_instr_long_addr[6]
port 292 nsew signal input
rlabel metal2 s 88480 0 88536 400 6 c1_o_instr_long_addr[7]
port 293 nsew signal input
rlabel metal2 s 69440 0 69496 400 6 c1_o_mem_addr[0]
port 294 nsew signal input
rlabel metal2 s 95648 0 95704 400 6 c1_o_mem_addr[10]
port 295 nsew signal input
rlabel metal2 s 97888 0 97944 400 6 c1_o_mem_addr[11]
port 296 nsew signal input
rlabel metal2 s 100128 0 100184 400 6 c1_o_mem_addr[12]
port 297 nsew signal input
rlabel metal2 s 102368 0 102424 400 6 c1_o_mem_addr[13]
port 298 nsew signal input
rlabel metal2 s 104608 0 104664 400 6 c1_o_mem_addr[14]
port 299 nsew signal input
rlabel metal2 s 106848 0 106904 400 6 c1_o_mem_addr[15]
port 300 nsew signal input
rlabel metal2 s 72352 0 72408 400 6 c1_o_mem_addr[1]
port 301 nsew signal input
rlabel metal2 s 75264 0 75320 400 6 c1_o_mem_addr[2]
port 302 nsew signal input
rlabel metal2 s 77952 0 78008 400 6 c1_o_mem_addr[3]
port 303 nsew signal input
rlabel metal2 s 80640 0 80696 400 6 c1_o_mem_addr[4]
port 304 nsew signal input
rlabel metal2 s 83328 0 83384 400 6 c1_o_mem_addr[5]
port 305 nsew signal input
rlabel metal2 s 86016 0 86072 400 6 c1_o_mem_addr[6]
port 306 nsew signal input
rlabel metal2 s 88704 0 88760 400 6 c1_o_mem_addr[7]
port 307 nsew signal input
rlabel metal2 s 91168 0 91224 400 6 c1_o_mem_addr[8]
port 308 nsew signal input
rlabel metal2 s 93408 0 93464 400 6 c1_o_mem_addr[9]
port 309 nsew signal input
rlabel metal2 s 69664 0 69720 400 6 c1_o_mem_data[0]
port 310 nsew signal input
rlabel metal2 s 95872 0 95928 400 6 c1_o_mem_data[10]
port 311 nsew signal input
rlabel metal2 s 98112 0 98168 400 6 c1_o_mem_data[11]
port 312 nsew signal input
rlabel metal2 s 100352 0 100408 400 6 c1_o_mem_data[12]
port 313 nsew signal input
rlabel metal2 s 102592 0 102648 400 6 c1_o_mem_data[13]
port 314 nsew signal input
rlabel metal2 s 104832 0 104888 400 6 c1_o_mem_data[14]
port 315 nsew signal input
rlabel metal2 s 107072 0 107128 400 6 c1_o_mem_data[15]
port 316 nsew signal input
rlabel metal2 s 72576 0 72632 400 6 c1_o_mem_data[1]
port 317 nsew signal input
rlabel metal2 s 75488 0 75544 400 6 c1_o_mem_data[2]
port 318 nsew signal input
rlabel metal2 s 78176 0 78232 400 6 c1_o_mem_data[3]
port 319 nsew signal input
rlabel metal2 s 80864 0 80920 400 6 c1_o_mem_data[4]
port 320 nsew signal input
rlabel metal2 s 83552 0 83608 400 6 c1_o_mem_data[5]
port 321 nsew signal input
rlabel metal2 s 86240 0 86296 400 6 c1_o_mem_data[6]
port 322 nsew signal input
rlabel metal2 s 88928 0 88984 400 6 c1_o_mem_data[7]
port 323 nsew signal input
rlabel metal2 s 91392 0 91448 400 6 c1_o_mem_data[8]
port 324 nsew signal input
rlabel metal2 s 93632 0 93688 400 6 c1_o_mem_data[9]
port 325 nsew signal input
rlabel metal2 s 69888 0 69944 400 6 c1_o_mem_high_addr[0]
port 326 nsew signal input
rlabel metal2 s 72800 0 72856 400 6 c1_o_mem_high_addr[1]
port 327 nsew signal input
rlabel metal2 s 75712 0 75768 400 6 c1_o_mem_high_addr[2]
port 328 nsew signal input
rlabel metal2 s 78400 0 78456 400 6 c1_o_mem_high_addr[3]
port 329 nsew signal input
rlabel metal2 s 81088 0 81144 400 6 c1_o_mem_high_addr[4]
port 330 nsew signal input
rlabel metal2 s 83776 0 83832 400 6 c1_o_mem_high_addr[5]
port 331 nsew signal input
rlabel metal2 s 86464 0 86520 400 6 c1_o_mem_high_addr[6]
port 332 nsew signal input
rlabel metal2 s 89152 0 89208 400 6 c1_o_mem_high_addr[7]
port 333 nsew signal input
rlabel metal2 s 66528 0 66584 400 6 c1_o_mem_long_mode
port 334 nsew signal input
rlabel metal2 s 66752 0 66808 400 6 c1_o_mem_req
port 335 nsew signal input
rlabel metal2 s 70112 0 70168 400 6 c1_o_mem_sel[0]
port 336 nsew signal input
rlabel metal2 s 73024 0 73080 400 6 c1_o_mem_sel[1]
port 337 nsew signal input
rlabel metal2 s 66976 0 67032 400 6 c1_o_mem_we
port 338 nsew signal input
rlabel metal2 s 67200 0 67256 400 6 c1_o_req_active
port 339 nsew signal input
rlabel metal2 s 70336 0 70392 400 6 c1_o_req_addr[0]
port 340 nsew signal input
rlabel metal2 s 96096 0 96152 400 6 c1_o_req_addr[10]
port 341 nsew signal input
rlabel metal2 s 98336 0 98392 400 6 c1_o_req_addr[11]
port 342 nsew signal input
rlabel metal2 s 100576 0 100632 400 6 c1_o_req_addr[12]
port 343 nsew signal input
rlabel metal2 s 102816 0 102872 400 6 c1_o_req_addr[13]
port 344 nsew signal input
rlabel metal2 s 105056 0 105112 400 6 c1_o_req_addr[14]
port 345 nsew signal input
rlabel metal2 s 107296 0 107352 400 6 c1_o_req_addr[15]
port 346 nsew signal input
rlabel metal2 s 73248 0 73304 400 6 c1_o_req_addr[1]
port 347 nsew signal input
rlabel metal2 s 75936 0 75992 400 6 c1_o_req_addr[2]
port 348 nsew signal input
rlabel metal2 s 78624 0 78680 400 6 c1_o_req_addr[3]
port 349 nsew signal input
rlabel metal2 s 81312 0 81368 400 6 c1_o_req_addr[4]
port 350 nsew signal input
rlabel metal2 s 84000 0 84056 400 6 c1_o_req_addr[5]
port 351 nsew signal input
rlabel metal2 s 86688 0 86744 400 6 c1_o_req_addr[6]
port 352 nsew signal input
rlabel metal2 s 89376 0 89432 400 6 c1_o_req_addr[7]
port 353 nsew signal input
rlabel metal2 s 91616 0 91672 400 6 c1_o_req_addr[8]
port 354 nsew signal input
rlabel metal2 s 93856 0 93912 400 6 c1_o_req_addr[9]
port 355 nsew signal input
rlabel metal2 s 67424 0 67480 400 6 c1_o_req_ppl_submit
port 356 nsew signal input
rlabel metal2 s 67648 0 67704 400 6 c1_rst
port 357 nsew signal output
rlabel metal2 s 70560 0 70616 400 6 c1_sr_bus_addr[0]
port 358 nsew signal input
rlabel metal2 s 96320 0 96376 400 6 c1_sr_bus_addr[10]
port 359 nsew signal input
rlabel metal2 s 98560 0 98616 400 6 c1_sr_bus_addr[11]
port 360 nsew signal input
rlabel metal2 s 100800 0 100856 400 6 c1_sr_bus_addr[12]
port 361 nsew signal input
rlabel metal2 s 103040 0 103096 400 6 c1_sr_bus_addr[13]
port 362 nsew signal input
rlabel metal2 s 105280 0 105336 400 6 c1_sr_bus_addr[14]
port 363 nsew signal input
rlabel metal2 s 107520 0 107576 400 6 c1_sr_bus_addr[15]
port 364 nsew signal input
rlabel metal2 s 73472 0 73528 400 6 c1_sr_bus_addr[1]
port 365 nsew signal input
rlabel metal2 s 76160 0 76216 400 6 c1_sr_bus_addr[2]
port 366 nsew signal input
rlabel metal2 s 78848 0 78904 400 6 c1_sr_bus_addr[3]
port 367 nsew signal input
rlabel metal2 s 81536 0 81592 400 6 c1_sr_bus_addr[4]
port 368 nsew signal input
rlabel metal2 s 84224 0 84280 400 6 c1_sr_bus_addr[5]
port 369 nsew signal input
rlabel metal2 s 86912 0 86968 400 6 c1_sr_bus_addr[6]
port 370 nsew signal input
rlabel metal2 s 89600 0 89656 400 6 c1_sr_bus_addr[7]
port 371 nsew signal input
rlabel metal2 s 91840 0 91896 400 6 c1_sr_bus_addr[8]
port 372 nsew signal input
rlabel metal2 s 94080 0 94136 400 6 c1_sr_bus_addr[9]
port 373 nsew signal input
rlabel metal2 s 70784 0 70840 400 6 c1_sr_bus_data_o[0]
port 374 nsew signal input
rlabel metal2 s 96544 0 96600 400 6 c1_sr_bus_data_o[10]
port 375 nsew signal input
rlabel metal2 s 98784 0 98840 400 6 c1_sr_bus_data_o[11]
port 376 nsew signal input
rlabel metal2 s 101024 0 101080 400 6 c1_sr_bus_data_o[12]
port 377 nsew signal input
rlabel metal2 s 103264 0 103320 400 6 c1_sr_bus_data_o[13]
port 378 nsew signal input
rlabel metal2 s 105504 0 105560 400 6 c1_sr_bus_data_o[14]
port 379 nsew signal input
rlabel metal2 s 107744 0 107800 400 6 c1_sr_bus_data_o[15]
port 380 nsew signal input
rlabel metal2 s 73696 0 73752 400 6 c1_sr_bus_data_o[1]
port 381 nsew signal input
rlabel metal2 s 76384 0 76440 400 6 c1_sr_bus_data_o[2]
port 382 nsew signal input
rlabel metal2 s 79072 0 79128 400 6 c1_sr_bus_data_o[3]
port 383 nsew signal input
rlabel metal2 s 81760 0 81816 400 6 c1_sr_bus_data_o[4]
port 384 nsew signal input
rlabel metal2 s 84448 0 84504 400 6 c1_sr_bus_data_o[5]
port 385 nsew signal input
rlabel metal2 s 87136 0 87192 400 6 c1_sr_bus_data_o[6]
port 386 nsew signal input
rlabel metal2 s 89824 0 89880 400 6 c1_sr_bus_data_o[7]
port 387 nsew signal input
rlabel metal2 s 92064 0 92120 400 6 c1_sr_bus_data_o[8]
port 388 nsew signal input
rlabel metal2 s 94304 0 94360 400 6 c1_sr_bus_data_o[9]
port 389 nsew signal input
rlabel metal2 s 67872 0 67928 400 6 c1_sr_bus_we
port 390 nsew signal input
rlabel metal2 s 48608 0 48664 400 6 core_clock
port 391 nsew signal input
rlabel metal2 s 48832 0 48888 400 6 core_reset
port 392 nsew signal input
rlabel metal2 s 3024 36600 3080 37000 6 dcache_mem_ack
port 393 nsew signal input
rlabel metal2 s 13776 36600 13832 37000 6 dcache_mem_addr[0]
port 394 nsew signal output
rlabel metal2 s 71120 36600 71176 37000 6 dcache_mem_addr[10]
port 395 nsew signal output
rlabel metal2 s 76496 36600 76552 37000 6 dcache_mem_addr[11]
port 396 nsew signal output
rlabel metal2 s 81872 36600 81928 37000 6 dcache_mem_addr[12]
port 397 nsew signal output
rlabel metal2 s 87248 36600 87304 37000 6 dcache_mem_addr[13]
port 398 nsew signal output
rlabel metal2 s 92624 36600 92680 37000 6 dcache_mem_addr[14]
port 399 nsew signal output
rlabel metal2 s 98000 36600 98056 37000 6 dcache_mem_addr[15]
port 400 nsew signal output
rlabel metal2 s 103376 36600 103432 37000 6 dcache_mem_addr[16]
port 401 nsew signal output
rlabel metal2 s 105168 36600 105224 37000 6 dcache_mem_addr[17]
port 402 nsew signal output
rlabel metal2 s 106960 36600 107016 37000 6 dcache_mem_addr[18]
port 403 nsew signal output
rlabel metal2 s 108752 36600 108808 37000 6 dcache_mem_addr[19]
port 404 nsew signal output
rlabel metal2 s 20944 36600 21000 37000 6 dcache_mem_addr[1]
port 405 nsew signal output
rlabel metal2 s 110544 36600 110600 37000 6 dcache_mem_addr[20]
port 406 nsew signal output
rlabel metal2 s 112336 36600 112392 37000 6 dcache_mem_addr[21]
port 407 nsew signal output
rlabel metal2 s 114128 36600 114184 37000 6 dcache_mem_addr[22]
port 408 nsew signal output
rlabel metal2 s 115920 36600 115976 37000 6 dcache_mem_addr[23]
port 409 nsew signal output
rlabel metal2 s 28112 36600 28168 37000 6 dcache_mem_addr[2]
port 410 nsew signal output
rlabel metal2 s 33488 36600 33544 37000 6 dcache_mem_addr[3]
port 411 nsew signal output
rlabel metal2 s 38864 36600 38920 37000 6 dcache_mem_addr[4]
port 412 nsew signal output
rlabel metal2 s 44240 36600 44296 37000 6 dcache_mem_addr[5]
port 413 nsew signal output
rlabel metal2 s 49616 36600 49672 37000 6 dcache_mem_addr[6]
port 414 nsew signal output
rlabel metal2 s 54992 36600 55048 37000 6 dcache_mem_addr[7]
port 415 nsew signal output
rlabel metal2 s 60368 36600 60424 37000 6 dcache_mem_addr[8]
port 416 nsew signal output
rlabel metal2 s 65744 36600 65800 37000 6 dcache_mem_addr[9]
port 417 nsew signal output
rlabel metal2 s 3920 36600 3976 37000 6 dcache_mem_cache_enable
port 418 nsew signal output
rlabel metal2 s 4816 36600 4872 37000 6 dcache_mem_exception
port 419 nsew signal input
rlabel metal2 s 14672 36600 14728 37000 6 dcache_mem_i_data[0]
port 420 nsew signal output
rlabel metal2 s 72016 36600 72072 37000 6 dcache_mem_i_data[10]
port 421 nsew signal output
rlabel metal2 s 77392 36600 77448 37000 6 dcache_mem_i_data[11]
port 422 nsew signal output
rlabel metal2 s 82768 36600 82824 37000 6 dcache_mem_i_data[12]
port 423 nsew signal output
rlabel metal2 s 88144 36600 88200 37000 6 dcache_mem_i_data[13]
port 424 nsew signal output
rlabel metal2 s 93520 36600 93576 37000 6 dcache_mem_i_data[14]
port 425 nsew signal output
rlabel metal2 s 98896 36600 98952 37000 6 dcache_mem_i_data[15]
port 426 nsew signal output
rlabel metal2 s 21840 36600 21896 37000 6 dcache_mem_i_data[1]
port 427 nsew signal output
rlabel metal2 s 29008 36600 29064 37000 6 dcache_mem_i_data[2]
port 428 nsew signal output
rlabel metal2 s 34384 36600 34440 37000 6 dcache_mem_i_data[3]
port 429 nsew signal output
rlabel metal2 s 39760 36600 39816 37000 6 dcache_mem_i_data[4]
port 430 nsew signal output
rlabel metal2 s 45136 36600 45192 37000 6 dcache_mem_i_data[5]
port 431 nsew signal output
rlabel metal2 s 50512 36600 50568 37000 6 dcache_mem_i_data[6]
port 432 nsew signal output
rlabel metal2 s 55888 36600 55944 37000 6 dcache_mem_i_data[7]
port 433 nsew signal output
rlabel metal2 s 61264 36600 61320 37000 6 dcache_mem_i_data[8]
port 434 nsew signal output
rlabel metal2 s 66640 36600 66696 37000 6 dcache_mem_i_data[9]
port 435 nsew signal output
rlabel metal2 s 15568 36600 15624 37000 6 dcache_mem_o_data[0]
port 436 nsew signal input
rlabel metal2 s 72912 36600 72968 37000 6 dcache_mem_o_data[10]
port 437 nsew signal input
rlabel metal2 s 78288 36600 78344 37000 6 dcache_mem_o_data[11]
port 438 nsew signal input
rlabel metal2 s 83664 36600 83720 37000 6 dcache_mem_o_data[12]
port 439 nsew signal input
rlabel metal2 s 89040 36600 89096 37000 6 dcache_mem_o_data[13]
port 440 nsew signal input
rlabel metal2 s 94416 36600 94472 37000 6 dcache_mem_o_data[14]
port 441 nsew signal input
rlabel metal2 s 99792 36600 99848 37000 6 dcache_mem_o_data[15]
port 442 nsew signal input
rlabel metal2 s 22736 36600 22792 37000 6 dcache_mem_o_data[1]
port 443 nsew signal input
rlabel metal2 s 29904 36600 29960 37000 6 dcache_mem_o_data[2]
port 444 nsew signal input
rlabel metal2 s 35280 36600 35336 37000 6 dcache_mem_o_data[3]
port 445 nsew signal input
rlabel metal2 s 40656 36600 40712 37000 6 dcache_mem_o_data[4]
port 446 nsew signal input
rlabel metal2 s 46032 36600 46088 37000 6 dcache_mem_o_data[5]
port 447 nsew signal input
rlabel metal2 s 51408 36600 51464 37000 6 dcache_mem_o_data[6]
port 448 nsew signal input
rlabel metal2 s 56784 36600 56840 37000 6 dcache_mem_o_data[7]
port 449 nsew signal input
rlabel metal2 s 62160 36600 62216 37000 6 dcache_mem_o_data[8]
port 450 nsew signal input
rlabel metal2 s 67536 36600 67592 37000 6 dcache_mem_o_data[9]
port 451 nsew signal input
rlabel metal2 s 5712 36600 5768 37000 6 dcache_mem_req
port 452 nsew signal output
rlabel metal2 s 16464 36600 16520 37000 6 dcache_mem_sel[0]
port 453 nsew signal output
rlabel metal2 s 23632 36600 23688 37000 6 dcache_mem_sel[1]
port 454 nsew signal output
rlabel metal2 s 6608 36600 6664 37000 6 dcache_mem_we
port 455 nsew signal output
rlabel metal2 s 7504 36600 7560 37000 6 dcache_rst
port 456 nsew signal output
rlabel metal2 s 8400 36600 8456 37000 6 dcache_wb_4_burst
port 457 nsew signal input
rlabel metal2 s 9296 36600 9352 37000 6 dcache_wb_ack
port 458 nsew signal output
rlabel metal2 s 17360 36600 17416 37000 6 dcache_wb_adr[0]
port 459 nsew signal input
rlabel metal2 s 73808 36600 73864 37000 6 dcache_wb_adr[10]
port 460 nsew signal input
rlabel metal2 s 79184 36600 79240 37000 6 dcache_wb_adr[11]
port 461 nsew signal input
rlabel metal2 s 84560 36600 84616 37000 6 dcache_wb_adr[12]
port 462 nsew signal input
rlabel metal2 s 89936 36600 89992 37000 6 dcache_wb_adr[13]
port 463 nsew signal input
rlabel metal2 s 95312 36600 95368 37000 6 dcache_wb_adr[14]
port 464 nsew signal input
rlabel metal2 s 100688 36600 100744 37000 6 dcache_wb_adr[15]
port 465 nsew signal input
rlabel metal2 s 104272 36600 104328 37000 6 dcache_wb_adr[16]
port 466 nsew signal input
rlabel metal2 s 106064 36600 106120 37000 6 dcache_wb_adr[17]
port 467 nsew signal input
rlabel metal2 s 107856 36600 107912 37000 6 dcache_wb_adr[18]
port 468 nsew signal input
rlabel metal2 s 109648 36600 109704 37000 6 dcache_wb_adr[19]
port 469 nsew signal input
rlabel metal2 s 24528 36600 24584 37000 6 dcache_wb_adr[1]
port 470 nsew signal input
rlabel metal2 s 111440 36600 111496 37000 6 dcache_wb_adr[20]
port 471 nsew signal input
rlabel metal2 s 113232 36600 113288 37000 6 dcache_wb_adr[21]
port 472 nsew signal input
rlabel metal2 s 115024 36600 115080 37000 6 dcache_wb_adr[22]
port 473 nsew signal input
rlabel metal2 s 116816 36600 116872 37000 6 dcache_wb_adr[23]
port 474 nsew signal input
rlabel metal2 s 30800 36600 30856 37000 6 dcache_wb_adr[2]
port 475 nsew signal input
rlabel metal2 s 36176 36600 36232 37000 6 dcache_wb_adr[3]
port 476 nsew signal input
rlabel metal2 s 41552 36600 41608 37000 6 dcache_wb_adr[4]
port 477 nsew signal input
rlabel metal2 s 46928 36600 46984 37000 6 dcache_wb_adr[5]
port 478 nsew signal input
rlabel metal2 s 52304 36600 52360 37000 6 dcache_wb_adr[6]
port 479 nsew signal input
rlabel metal2 s 57680 36600 57736 37000 6 dcache_wb_adr[7]
port 480 nsew signal input
rlabel metal2 s 63056 36600 63112 37000 6 dcache_wb_adr[8]
port 481 nsew signal input
rlabel metal2 s 68432 36600 68488 37000 6 dcache_wb_adr[9]
port 482 nsew signal input
rlabel metal2 s 10192 36600 10248 37000 6 dcache_wb_cyc
port 483 nsew signal input
rlabel metal2 s 11088 36600 11144 37000 6 dcache_wb_err
port 484 nsew signal output
rlabel metal2 s 18256 36600 18312 37000 6 dcache_wb_i_dat[0]
port 485 nsew signal output
rlabel metal2 s 74704 36600 74760 37000 6 dcache_wb_i_dat[10]
port 486 nsew signal output
rlabel metal2 s 80080 36600 80136 37000 6 dcache_wb_i_dat[11]
port 487 nsew signal output
rlabel metal2 s 85456 36600 85512 37000 6 dcache_wb_i_dat[12]
port 488 nsew signal output
rlabel metal2 s 90832 36600 90888 37000 6 dcache_wb_i_dat[13]
port 489 nsew signal output
rlabel metal2 s 96208 36600 96264 37000 6 dcache_wb_i_dat[14]
port 490 nsew signal output
rlabel metal2 s 101584 36600 101640 37000 6 dcache_wb_i_dat[15]
port 491 nsew signal output
rlabel metal2 s 25424 36600 25480 37000 6 dcache_wb_i_dat[1]
port 492 nsew signal output
rlabel metal2 s 31696 36600 31752 37000 6 dcache_wb_i_dat[2]
port 493 nsew signal output
rlabel metal2 s 37072 36600 37128 37000 6 dcache_wb_i_dat[3]
port 494 nsew signal output
rlabel metal2 s 42448 36600 42504 37000 6 dcache_wb_i_dat[4]
port 495 nsew signal output
rlabel metal2 s 47824 36600 47880 37000 6 dcache_wb_i_dat[5]
port 496 nsew signal output
rlabel metal2 s 53200 36600 53256 37000 6 dcache_wb_i_dat[6]
port 497 nsew signal output
rlabel metal2 s 58576 36600 58632 37000 6 dcache_wb_i_dat[7]
port 498 nsew signal output
rlabel metal2 s 63952 36600 64008 37000 6 dcache_wb_i_dat[8]
port 499 nsew signal output
rlabel metal2 s 69328 36600 69384 37000 6 dcache_wb_i_dat[9]
port 500 nsew signal output
rlabel metal2 s 19152 36600 19208 37000 6 dcache_wb_o_dat[0]
port 501 nsew signal input
rlabel metal2 s 75600 36600 75656 37000 6 dcache_wb_o_dat[10]
port 502 nsew signal input
rlabel metal2 s 80976 36600 81032 37000 6 dcache_wb_o_dat[11]
port 503 nsew signal input
rlabel metal2 s 86352 36600 86408 37000 6 dcache_wb_o_dat[12]
port 504 nsew signal input
rlabel metal2 s 91728 36600 91784 37000 6 dcache_wb_o_dat[13]
port 505 nsew signal input
rlabel metal2 s 97104 36600 97160 37000 6 dcache_wb_o_dat[14]
port 506 nsew signal input
rlabel metal2 s 102480 36600 102536 37000 6 dcache_wb_o_dat[15]
port 507 nsew signal input
rlabel metal2 s 26320 36600 26376 37000 6 dcache_wb_o_dat[1]
port 508 nsew signal input
rlabel metal2 s 32592 36600 32648 37000 6 dcache_wb_o_dat[2]
port 509 nsew signal input
rlabel metal2 s 37968 36600 38024 37000 6 dcache_wb_o_dat[3]
port 510 nsew signal input
rlabel metal2 s 43344 36600 43400 37000 6 dcache_wb_o_dat[4]
port 511 nsew signal input
rlabel metal2 s 48720 36600 48776 37000 6 dcache_wb_o_dat[5]
port 512 nsew signal input
rlabel metal2 s 54096 36600 54152 37000 6 dcache_wb_o_dat[6]
port 513 nsew signal input
rlabel metal2 s 59472 36600 59528 37000 6 dcache_wb_o_dat[7]
port 514 nsew signal input
rlabel metal2 s 64848 36600 64904 37000 6 dcache_wb_o_dat[8]
port 515 nsew signal input
rlabel metal2 s 70224 36600 70280 37000 6 dcache_wb_o_dat[9]
port 516 nsew signal input
rlabel metal2 s 20048 36600 20104 37000 6 dcache_wb_sel[0]
port 517 nsew signal input
rlabel metal2 s 27216 36600 27272 37000 6 dcache_wb_sel[1]
port 518 nsew signal input
rlabel metal2 s 11984 36600 12040 37000 6 dcache_wb_stb
port 519 nsew signal input
rlabel metal2 s 12880 36600 12936 37000 6 dcache_wb_we
port 520 nsew signal input
rlabel metal3 s 0 3136 400 3192 6 ic0_mem_ack
port 521 nsew signal input
rlabel metal3 s 0 6496 400 6552 6 ic0_mem_addr[0]
port 522 nsew signal output
rlabel metal3 s 0 20608 400 20664 6 ic0_mem_addr[10]
port 523 nsew signal output
rlabel metal3 s 0 21952 400 22008 6 ic0_mem_addr[11]
port 524 nsew signal output
rlabel metal3 s 0 23296 400 23352 6 ic0_mem_addr[12]
port 525 nsew signal output
rlabel metal3 s 0 24640 400 24696 6 ic0_mem_addr[13]
port 526 nsew signal output
rlabel metal3 s 0 25984 400 26040 6 ic0_mem_addr[14]
port 527 nsew signal output
rlabel metal3 s 0 27328 400 27384 6 ic0_mem_addr[15]
port 528 nsew signal output
rlabel metal3 s 0 8176 400 8232 6 ic0_mem_addr[1]
port 529 nsew signal output
rlabel metal3 s 0 9856 400 9912 6 ic0_mem_addr[2]
port 530 nsew signal output
rlabel metal3 s 0 11200 400 11256 6 ic0_mem_addr[3]
port 531 nsew signal output
rlabel metal3 s 0 12544 400 12600 6 ic0_mem_addr[4]
port 532 nsew signal output
rlabel metal3 s 0 13888 400 13944 6 ic0_mem_addr[5]
port 533 nsew signal output
rlabel metal3 s 0 15232 400 15288 6 ic0_mem_addr[6]
port 534 nsew signal output
rlabel metal3 s 0 16576 400 16632 6 ic0_mem_addr[7]
port 535 nsew signal output
rlabel metal3 s 0 17920 400 17976 6 ic0_mem_addr[8]
port 536 nsew signal output
rlabel metal3 s 0 19264 400 19320 6 ic0_mem_addr[9]
port 537 nsew signal output
rlabel metal3 s 0 3472 400 3528 6 ic0_mem_cache_flush
port 538 nsew signal output
rlabel metal3 s 0 6832 400 6888 6 ic0_mem_data[0]
port 539 nsew signal input
rlabel metal3 s 0 20944 400 21000 6 ic0_mem_data[10]
port 540 nsew signal input
rlabel metal3 s 0 22288 400 22344 6 ic0_mem_data[11]
port 541 nsew signal input
rlabel metal3 s 0 23632 400 23688 6 ic0_mem_data[12]
port 542 nsew signal input
rlabel metal3 s 0 24976 400 25032 6 ic0_mem_data[13]
port 543 nsew signal input
rlabel metal3 s 0 26320 400 26376 6 ic0_mem_data[14]
port 544 nsew signal input
rlabel metal3 s 0 27664 400 27720 6 ic0_mem_data[15]
port 545 nsew signal input
rlabel metal3 s 0 28672 400 28728 6 ic0_mem_data[16]
port 546 nsew signal input
rlabel metal3 s 0 29008 400 29064 6 ic0_mem_data[17]
port 547 nsew signal input
rlabel metal3 s 0 29344 400 29400 6 ic0_mem_data[18]
port 548 nsew signal input
rlabel metal3 s 0 29680 400 29736 6 ic0_mem_data[19]
port 549 nsew signal input
rlabel metal3 s 0 8512 400 8568 6 ic0_mem_data[1]
port 550 nsew signal input
rlabel metal3 s 0 30016 400 30072 6 ic0_mem_data[20]
port 551 nsew signal input
rlabel metal3 s 0 30352 400 30408 6 ic0_mem_data[21]
port 552 nsew signal input
rlabel metal3 s 0 30688 400 30744 6 ic0_mem_data[22]
port 553 nsew signal input
rlabel metal3 s 0 31024 400 31080 6 ic0_mem_data[23]
port 554 nsew signal input
rlabel metal3 s 0 31360 400 31416 6 ic0_mem_data[24]
port 555 nsew signal input
rlabel metal3 s 0 31696 400 31752 6 ic0_mem_data[25]
port 556 nsew signal input
rlabel metal3 s 0 32032 400 32088 6 ic0_mem_data[26]
port 557 nsew signal input
rlabel metal3 s 0 32368 400 32424 6 ic0_mem_data[27]
port 558 nsew signal input
rlabel metal3 s 0 32704 400 32760 6 ic0_mem_data[28]
port 559 nsew signal input
rlabel metal3 s 0 33040 400 33096 6 ic0_mem_data[29]
port 560 nsew signal input
rlabel metal3 s 0 10192 400 10248 6 ic0_mem_data[2]
port 561 nsew signal input
rlabel metal3 s 0 33376 400 33432 6 ic0_mem_data[30]
port 562 nsew signal input
rlabel metal3 s 0 33712 400 33768 6 ic0_mem_data[31]
port 563 nsew signal input
rlabel metal3 s 0 11536 400 11592 6 ic0_mem_data[3]
port 564 nsew signal input
rlabel metal3 s 0 12880 400 12936 6 ic0_mem_data[4]
port 565 nsew signal input
rlabel metal3 s 0 14224 400 14280 6 ic0_mem_data[5]
port 566 nsew signal input
rlabel metal3 s 0 15568 400 15624 6 ic0_mem_data[6]
port 567 nsew signal input
rlabel metal3 s 0 16912 400 16968 6 ic0_mem_data[7]
port 568 nsew signal input
rlabel metal3 s 0 18256 400 18312 6 ic0_mem_data[8]
port 569 nsew signal input
rlabel metal3 s 0 19600 400 19656 6 ic0_mem_data[9]
port 570 nsew signal input
rlabel metal3 s 0 3808 400 3864 6 ic0_mem_ppl_submit
port 571 nsew signal output
rlabel metal3 s 0 4144 400 4200 6 ic0_mem_req
port 572 nsew signal output
rlabel metal3 s 0 4480 400 4536 6 ic0_rst
port 573 nsew signal output
rlabel metal3 s 0 4816 400 4872 6 ic0_wb_ack
port 574 nsew signal output
rlabel metal3 s 0 7168 400 7224 6 ic0_wb_adr[0]
port 575 nsew signal input
rlabel metal3 s 0 21280 400 21336 6 ic0_wb_adr[10]
port 576 nsew signal input
rlabel metal3 s 0 22624 400 22680 6 ic0_wb_adr[11]
port 577 nsew signal input
rlabel metal3 s 0 23968 400 24024 6 ic0_wb_adr[12]
port 578 nsew signal input
rlabel metal3 s 0 25312 400 25368 6 ic0_wb_adr[13]
port 579 nsew signal input
rlabel metal3 s 0 26656 400 26712 6 ic0_wb_adr[14]
port 580 nsew signal input
rlabel metal3 s 0 28000 400 28056 6 ic0_wb_adr[15]
port 581 nsew signal input
rlabel metal3 s 0 8848 400 8904 6 ic0_wb_adr[1]
port 582 nsew signal input
rlabel metal3 s 0 10528 400 10584 6 ic0_wb_adr[2]
port 583 nsew signal input
rlabel metal3 s 0 11872 400 11928 6 ic0_wb_adr[3]
port 584 nsew signal input
rlabel metal3 s 0 13216 400 13272 6 ic0_wb_adr[4]
port 585 nsew signal input
rlabel metal3 s 0 14560 400 14616 6 ic0_wb_adr[5]
port 586 nsew signal input
rlabel metal3 s 0 15904 400 15960 6 ic0_wb_adr[6]
port 587 nsew signal input
rlabel metal3 s 0 17248 400 17304 6 ic0_wb_adr[7]
port 588 nsew signal input
rlabel metal3 s 0 18592 400 18648 6 ic0_wb_adr[8]
port 589 nsew signal input
rlabel metal3 s 0 19936 400 19992 6 ic0_wb_adr[9]
port 590 nsew signal input
rlabel metal3 s 0 5152 400 5208 6 ic0_wb_cyc
port 591 nsew signal input
rlabel metal3 s 0 5488 400 5544 6 ic0_wb_err
port 592 nsew signal output
rlabel metal3 s 0 7504 400 7560 6 ic0_wb_i_dat[0]
port 593 nsew signal output
rlabel metal3 s 0 21616 400 21672 6 ic0_wb_i_dat[10]
port 594 nsew signal output
rlabel metal3 s 0 22960 400 23016 6 ic0_wb_i_dat[11]
port 595 nsew signal output
rlabel metal3 s 0 24304 400 24360 6 ic0_wb_i_dat[12]
port 596 nsew signal output
rlabel metal3 s 0 25648 400 25704 6 ic0_wb_i_dat[13]
port 597 nsew signal output
rlabel metal3 s 0 26992 400 27048 6 ic0_wb_i_dat[14]
port 598 nsew signal output
rlabel metal3 s 0 28336 400 28392 6 ic0_wb_i_dat[15]
port 599 nsew signal output
rlabel metal3 s 0 9184 400 9240 6 ic0_wb_i_dat[1]
port 600 nsew signal output
rlabel metal3 s 0 10864 400 10920 6 ic0_wb_i_dat[2]
port 601 nsew signal output
rlabel metal3 s 0 12208 400 12264 6 ic0_wb_i_dat[3]
port 602 nsew signal output
rlabel metal3 s 0 13552 400 13608 6 ic0_wb_i_dat[4]
port 603 nsew signal output
rlabel metal3 s 0 14896 400 14952 6 ic0_wb_i_dat[5]
port 604 nsew signal output
rlabel metal3 s 0 16240 400 16296 6 ic0_wb_i_dat[6]
port 605 nsew signal output
rlabel metal3 s 0 17584 400 17640 6 ic0_wb_i_dat[7]
port 606 nsew signal output
rlabel metal3 s 0 18928 400 18984 6 ic0_wb_i_dat[8]
port 607 nsew signal output
rlabel metal3 s 0 20272 400 20328 6 ic0_wb_i_dat[9]
port 608 nsew signal output
rlabel metal3 s 0 7840 400 7896 6 ic0_wb_sel[0]
port 609 nsew signal input
rlabel metal3 s 0 9520 400 9576 6 ic0_wb_sel[1]
port 610 nsew signal input
rlabel metal3 s 0 5824 400 5880 6 ic0_wb_stb
port 611 nsew signal input
rlabel metal3 s 0 6160 400 6216 6 ic0_wb_we
port 612 nsew signal input
rlabel metal3 s 119600 3136 120000 3192 6 ic1_mem_ack
port 613 nsew signal input
rlabel metal3 s 119600 6496 120000 6552 6 ic1_mem_addr[0]
port 614 nsew signal output
rlabel metal3 s 119600 20608 120000 20664 6 ic1_mem_addr[10]
port 615 nsew signal output
rlabel metal3 s 119600 21952 120000 22008 6 ic1_mem_addr[11]
port 616 nsew signal output
rlabel metal3 s 119600 23296 120000 23352 6 ic1_mem_addr[12]
port 617 nsew signal output
rlabel metal3 s 119600 24640 120000 24696 6 ic1_mem_addr[13]
port 618 nsew signal output
rlabel metal3 s 119600 25984 120000 26040 6 ic1_mem_addr[14]
port 619 nsew signal output
rlabel metal3 s 119600 27328 120000 27384 6 ic1_mem_addr[15]
port 620 nsew signal output
rlabel metal3 s 119600 8176 120000 8232 6 ic1_mem_addr[1]
port 621 nsew signal output
rlabel metal3 s 119600 9856 120000 9912 6 ic1_mem_addr[2]
port 622 nsew signal output
rlabel metal3 s 119600 11200 120000 11256 6 ic1_mem_addr[3]
port 623 nsew signal output
rlabel metal3 s 119600 12544 120000 12600 6 ic1_mem_addr[4]
port 624 nsew signal output
rlabel metal3 s 119600 13888 120000 13944 6 ic1_mem_addr[5]
port 625 nsew signal output
rlabel metal3 s 119600 15232 120000 15288 6 ic1_mem_addr[6]
port 626 nsew signal output
rlabel metal3 s 119600 16576 120000 16632 6 ic1_mem_addr[7]
port 627 nsew signal output
rlabel metal3 s 119600 17920 120000 17976 6 ic1_mem_addr[8]
port 628 nsew signal output
rlabel metal3 s 119600 19264 120000 19320 6 ic1_mem_addr[9]
port 629 nsew signal output
rlabel metal3 s 119600 3472 120000 3528 6 ic1_mem_cache_flush
port 630 nsew signal output
rlabel metal3 s 119600 6832 120000 6888 6 ic1_mem_data[0]
port 631 nsew signal input
rlabel metal3 s 119600 20944 120000 21000 6 ic1_mem_data[10]
port 632 nsew signal input
rlabel metal3 s 119600 22288 120000 22344 6 ic1_mem_data[11]
port 633 nsew signal input
rlabel metal3 s 119600 23632 120000 23688 6 ic1_mem_data[12]
port 634 nsew signal input
rlabel metal3 s 119600 24976 120000 25032 6 ic1_mem_data[13]
port 635 nsew signal input
rlabel metal3 s 119600 26320 120000 26376 6 ic1_mem_data[14]
port 636 nsew signal input
rlabel metal3 s 119600 27664 120000 27720 6 ic1_mem_data[15]
port 637 nsew signal input
rlabel metal3 s 119600 28672 120000 28728 6 ic1_mem_data[16]
port 638 nsew signal input
rlabel metal3 s 119600 29008 120000 29064 6 ic1_mem_data[17]
port 639 nsew signal input
rlabel metal3 s 119600 29344 120000 29400 6 ic1_mem_data[18]
port 640 nsew signal input
rlabel metal3 s 119600 29680 120000 29736 6 ic1_mem_data[19]
port 641 nsew signal input
rlabel metal3 s 119600 8512 120000 8568 6 ic1_mem_data[1]
port 642 nsew signal input
rlabel metal3 s 119600 30016 120000 30072 6 ic1_mem_data[20]
port 643 nsew signal input
rlabel metal3 s 119600 30352 120000 30408 6 ic1_mem_data[21]
port 644 nsew signal input
rlabel metal3 s 119600 30688 120000 30744 6 ic1_mem_data[22]
port 645 nsew signal input
rlabel metal3 s 119600 31024 120000 31080 6 ic1_mem_data[23]
port 646 nsew signal input
rlabel metal3 s 119600 31360 120000 31416 6 ic1_mem_data[24]
port 647 nsew signal input
rlabel metal3 s 119600 31696 120000 31752 6 ic1_mem_data[25]
port 648 nsew signal input
rlabel metal3 s 119600 32032 120000 32088 6 ic1_mem_data[26]
port 649 nsew signal input
rlabel metal3 s 119600 32368 120000 32424 6 ic1_mem_data[27]
port 650 nsew signal input
rlabel metal3 s 119600 32704 120000 32760 6 ic1_mem_data[28]
port 651 nsew signal input
rlabel metal3 s 119600 33040 120000 33096 6 ic1_mem_data[29]
port 652 nsew signal input
rlabel metal3 s 119600 10192 120000 10248 6 ic1_mem_data[2]
port 653 nsew signal input
rlabel metal3 s 119600 33376 120000 33432 6 ic1_mem_data[30]
port 654 nsew signal input
rlabel metal3 s 119600 33712 120000 33768 6 ic1_mem_data[31]
port 655 nsew signal input
rlabel metal3 s 119600 11536 120000 11592 6 ic1_mem_data[3]
port 656 nsew signal input
rlabel metal3 s 119600 12880 120000 12936 6 ic1_mem_data[4]
port 657 nsew signal input
rlabel metal3 s 119600 14224 120000 14280 6 ic1_mem_data[5]
port 658 nsew signal input
rlabel metal3 s 119600 15568 120000 15624 6 ic1_mem_data[6]
port 659 nsew signal input
rlabel metal3 s 119600 16912 120000 16968 6 ic1_mem_data[7]
port 660 nsew signal input
rlabel metal3 s 119600 18256 120000 18312 6 ic1_mem_data[8]
port 661 nsew signal input
rlabel metal3 s 119600 19600 120000 19656 6 ic1_mem_data[9]
port 662 nsew signal input
rlabel metal3 s 119600 3808 120000 3864 6 ic1_mem_ppl_submit
port 663 nsew signal output
rlabel metal3 s 119600 4144 120000 4200 6 ic1_mem_req
port 664 nsew signal output
rlabel metal3 s 119600 4480 120000 4536 6 ic1_rst
port 665 nsew signal output
rlabel metal3 s 119600 4816 120000 4872 6 ic1_wb_ack
port 666 nsew signal output
rlabel metal3 s 119600 7168 120000 7224 6 ic1_wb_adr[0]
port 667 nsew signal input
rlabel metal3 s 119600 21280 120000 21336 6 ic1_wb_adr[10]
port 668 nsew signal input
rlabel metal3 s 119600 22624 120000 22680 6 ic1_wb_adr[11]
port 669 nsew signal input
rlabel metal3 s 119600 23968 120000 24024 6 ic1_wb_adr[12]
port 670 nsew signal input
rlabel metal3 s 119600 25312 120000 25368 6 ic1_wb_adr[13]
port 671 nsew signal input
rlabel metal3 s 119600 26656 120000 26712 6 ic1_wb_adr[14]
port 672 nsew signal input
rlabel metal3 s 119600 28000 120000 28056 6 ic1_wb_adr[15]
port 673 nsew signal input
rlabel metal3 s 119600 8848 120000 8904 6 ic1_wb_adr[1]
port 674 nsew signal input
rlabel metal3 s 119600 10528 120000 10584 6 ic1_wb_adr[2]
port 675 nsew signal input
rlabel metal3 s 119600 11872 120000 11928 6 ic1_wb_adr[3]
port 676 nsew signal input
rlabel metal3 s 119600 13216 120000 13272 6 ic1_wb_adr[4]
port 677 nsew signal input
rlabel metal3 s 119600 14560 120000 14616 6 ic1_wb_adr[5]
port 678 nsew signal input
rlabel metal3 s 119600 15904 120000 15960 6 ic1_wb_adr[6]
port 679 nsew signal input
rlabel metal3 s 119600 17248 120000 17304 6 ic1_wb_adr[7]
port 680 nsew signal input
rlabel metal3 s 119600 18592 120000 18648 6 ic1_wb_adr[8]
port 681 nsew signal input
rlabel metal3 s 119600 19936 120000 19992 6 ic1_wb_adr[9]
port 682 nsew signal input
rlabel metal3 s 119600 5152 120000 5208 6 ic1_wb_cyc
port 683 nsew signal input
rlabel metal3 s 119600 5488 120000 5544 6 ic1_wb_err
port 684 nsew signal output
rlabel metal3 s 119600 7504 120000 7560 6 ic1_wb_i_dat[0]
port 685 nsew signal output
rlabel metal3 s 119600 21616 120000 21672 6 ic1_wb_i_dat[10]
port 686 nsew signal output
rlabel metal3 s 119600 22960 120000 23016 6 ic1_wb_i_dat[11]
port 687 nsew signal output
rlabel metal3 s 119600 24304 120000 24360 6 ic1_wb_i_dat[12]
port 688 nsew signal output
rlabel metal3 s 119600 25648 120000 25704 6 ic1_wb_i_dat[13]
port 689 nsew signal output
rlabel metal3 s 119600 26992 120000 27048 6 ic1_wb_i_dat[14]
port 690 nsew signal output
rlabel metal3 s 119600 28336 120000 28392 6 ic1_wb_i_dat[15]
port 691 nsew signal output
rlabel metal3 s 119600 9184 120000 9240 6 ic1_wb_i_dat[1]
port 692 nsew signal output
rlabel metal3 s 119600 10864 120000 10920 6 ic1_wb_i_dat[2]
port 693 nsew signal output
rlabel metal3 s 119600 12208 120000 12264 6 ic1_wb_i_dat[3]
port 694 nsew signal output
rlabel metal3 s 119600 13552 120000 13608 6 ic1_wb_i_dat[4]
port 695 nsew signal output
rlabel metal3 s 119600 14896 120000 14952 6 ic1_wb_i_dat[5]
port 696 nsew signal output
rlabel metal3 s 119600 16240 120000 16296 6 ic1_wb_i_dat[6]
port 697 nsew signal output
rlabel metal3 s 119600 17584 120000 17640 6 ic1_wb_i_dat[7]
port 698 nsew signal output
rlabel metal3 s 119600 18928 120000 18984 6 ic1_wb_i_dat[8]
port 699 nsew signal output
rlabel metal3 s 119600 20272 120000 20328 6 ic1_wb_i_dat[9]
port 700 nsew signal output
rlabel metal3 s 119600 7840 120000 7896 6 ic1_wb_sel[0]
port 701 nsew signal input
rlabel metal3 s 119600 9520 120000 9576 6 ic1_wb_sel[1]
port 702 nsew signal input
rlabel metal3 s 119600 5824 120000 5880 6 ic1_wb_stb
port 703 nsew signal input
rlabel metal3 s 119600 6160 120000 6216 6 ic1_wb_we
port 704 nsew signal input
rlabel metal2 s 49056 0 49112 400 6 inner_disable
port 705 nsew signal input
rlabel metal2 s 49280 0 49336 400 6 inner_embed_mode
port 706 nsew signal input
rlabel metal2 s 49504 0 49560 400 6 inner_ext_irq
port 707 nsew signal input
rlabel metal2 s 49728 0 49784 400 6 inner_wb_4_burst
port 708 nsew signal output
rlabel metal2 s 49952 0 50008 400 6 inner_wb_8_burst
port 709 nsew signal output
rlabel metal2 s 50176 0 50232 400 6 inner_wb_ack
port 710 nsew signal input
rlabel metal2 s 51296 0 51352 400 6 inner_wb_adr[0]
port 711 nsew signal output
rlabel metal2 s 58464 0 58520 400 6 inner_wb_adr[10]
port 712 nsew signal output
rlabel metal2 s 59136 0 59192 400 6 inner_wb_adr[11]
port 713 nsew signal output
rlabel metal2 s 59808 0 59864 400 6 inner_wb_adr[12]
port 714 nsew signal output
rlabel metal2 s 60480 0 60536 400 6 inner_wb_adr[13]
port 715 nsew signal output
rlabel metal2 s 61152 0 61208 400 6 inner_wb_adr[14]
port 716 nsew signal output
rlabel metal2 s 61824 0 61880 400 6 inner_wb_adr[15]
port 717 nsew signal output
rlabel metal2 s 62496 0 62552 400 6 inner_wb_adr[16]
port 718 nsew signal output
rlabel metal2 s 62720 0 62776 400 6 inner_wb_adr[17]
port 719 nsew signal output
rlabel metal2 s 62944 0 63000 400 6 inner_wb_adr[18]
port 720 nsew signal output
rlabel metal2 s 63168 0 63224 400 6 inner_wb_adr[19]
port 721 nsew signal output
rlabel metal2 s 52192 0 52248 400 6 inner_wb_adr[1]
port 722 nsew signal output
rlabel metal2 s 63392 0 63448 400 6 inner_wb_adr[20]
port 723 nsew signal output
rlabel metal2 s 63616 0 63672 400 6 inner_wb_adr[21]
port 724 nsew signal output
rlabel metal2 s 63840 0 63896 400 6 inner_wb_adr[22]
port 725 nsew signal output
rlabel metal2 s 64064 0 64120 400 6 inner_wb_adr[23]
port 726 nsew signal output
rlabel metal2 s 53088 0 53144 400 6 inner_wb_adr[2]
port 727 nsew signal output
rlabel metal2 s 53760 0 53816 400 6 inner_wb_adr[3]
port 728 nsew signal output
rlabel metal2 s 54432 0 54488 400 6 inner_wb_adr[4]
port 729 nsew signal output
rlabel metal2 s 55104 0 55160 400 6 inner_wb_adr[5]
port 730 nsew signal output
rlabel metal2 s 55776 0 55832 400 6 inner_wb_adr[6]
port 731 nsew signal output
rlabel metal2 s 56448 0 56504 400 6 inner_wb_adr[7]
port 732 nsew signal output
rlabel metal2 s 57120 0 57176 400 6 inner_wb_adr[8]
port 733 nsew signal output
rlabel metal2 s 57792 0 57848 400 6 inner_wb_adr[9]
port 734 nsew signal output
rlabel metal2 s 50400 0 50456 400 6 inner_wb_cyc
port 735 nsew signal output
rlabel metal2 s 50624 0 50680 400 6 inner_wb_err
port 736 nsew signal input
rlabel metal2 s 51520 0 51576 400 6 inner_wb_i_dat[0]
port 737 nsew signal input
rlabel metal2 s 58688 0 58744 400 6 inner_wb_i_dat[10]
port 738 nsew signal input
rlabel metal2 s 59360 0 59416 400 6 inner_wb_i_dat[11]
port 739 nsew signal input
rlabel metal2 s 60032 0 60088 400 6 inner_wb_i_dat[12]
port 740 nsew signal input
rlabel metal2 s 60704 0 60760 400 6 inner_wb_i_dat[13]
port 741 nsew signal input
rlabel metal2 s 61376 0 61432 400 6 inner_wb_i_dat[14]
port 742 nsew signal input
rlabel metal2 s 62048 0 62104 400 6 inner_wb_i_dat[15]
port 743 nsew signal input
rlabel metal2 s 52416 0 52472 400 6 inner_wb_i_dat[1]
port 744 nsew signal input
rlabel metal2 s 53312 0 53368 400 6 inner_wb_i_dat[2]
port 745 nsew signal input
rlabel metal2 s 53984 0 54040 400 6 inner_wb_i_dat[3]
port 746 nsew signal input
rlabel metal2 s 54656 0 54712 400 6 inner_wb_i_dat[4]
port 747 nsew signal input
rlabel metal2 s 55328 0 55384 400 6 inner_wb_i_dat[5]
port 748 nsew signal input
rlabel metal2 s 56000 0 56056 400 6 inner_wb_i_dat[6]
port 749 nsew signal input
rlabel metal2 s 56672 0 56728 400 6 inner_wb_i_dat[7]
port 750 nsew signal input
rlabel metal2 s 57344 0 57400 400 6 inner_wb_i_dat[8]
port 751 nsew signal input
rlabel metal2 s 58016 0 58072 400 6 inner_wb_i_dat[9]
port 752 nsew signal input
rlabel metal2 s 51744 0 51800 400 6 inner_wb_o_dat[0]
port 753 nsew signal output
rlabel metal2 s 58912 0 58968 400 6 inner_wb_o_dat[10]
port 754 nsew signal output
rlabel metal2 s 59584 0 59640 400 6 inner_wb_o_dat[11]
port 755 nsew signal output
rlabel metal2 s 60256 0 60312 400 6 inner_wb_o_dat[12]
port 756 nsew signal output
rlabel metal2 s 60928 0 60984 400 6 inner_wb_o_dat[13]
port 757 nsew signal output
rlabel metal2 s 61600 0 61656 400 6 inner_wb_o_dat[14]
port 758 nsew signal output
rlabel metal2 s 62272 0 62328 400 6 inner_wb_o_dat[15]
port 759 nsew signal output
rlabel metal2 s 52640 0 52696 400 6 inner_wb_o_dat[1]
port 760 nsew signal output
rlabel metal2 s 53536 0 53592 400 6 inner_wb_o_dat[2]
port 761 nsew signal output
rlabel metal2 s 54208 0 54264 400 6 inner_wb_o_dat[3]
port 762 nsew signal output
rlabel metal2 s 54880 0 54936 400 6 inner_wb_o_dat[4]
port 763 nsew signal output
rlabel metal2 s 55552 0 55608 400 6 inner_wb_o_dat[5]
port 764 nsew signal output
rlabel metal2 s 56224 0 56280 400 6 inner_wb_o_dat[6]
port 765 nsew signal output
rlabel metal2 s 56896 0 56952 400 6 inner_wb_o_dat[7]
port 766 nsew signal output
rlabel metal2 s 57568 0 57624 400 6 inner_wb_o_dat[8]
port 767 nsew signal output
rlabel metal2 s 58240 0 58296 400 6 inner_wb_o_dat[9]
port 768 nsew signal output
rlabel metal2 s 51968 0 52024 400 6 inner_wb_sel[0]
port 769 nsew signal output
rlabel metal2 s 52864 0 52920 400 6 inner_wb_sel[1]
port 770 nsew signal output
rlabel metal2 s 50848 0 50904 400 6 inner_wb_stb
port 771 nsew signal output
rlabel metal2 s 51072 0 51128 400 6 inner_wb_we
port 772 nsew signal output
rlabel metal4 s 2224 1538 2384 35310 6 vccd1
port 773 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 35310 6 vccd1
port 773 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 35310 6 vccd1
port 773 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 35310 6 vccd1
port 773 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 35310 6 vccd1
port 773 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 35310 6 vccd1
port 773 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 35310 6 vccd1
port 773 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 35310 6 vccd1
port 773 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 35310 6 vssd1
port 774 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 35310 6 vssd1
port 774 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 35310 6 vssd1
port 774 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 35310 6 vssd1
port 774 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 35310 6 vssd1
port 774 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 35310 6 vssd1
port 774 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 35310 6 vssd1
port 774 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 35310 6 vssd1
port 774 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 120000 37000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 12425958
string GDS_FILE /home/piotro/caravel_user_project/openlane/inner_interconnect/runs/23_11_15_18_38/results/signoff/interconnect_inner.magic.gds
string GDS_START 480556
<< end >>

