magic
tech sky130B
magscale 1 2
timestamp 1663070775
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 658 1368 39362 37584
<< metal2 >>
rect 662 39200 718 40000
rect 1766 39200 1822 40000
rect 2870 39200 2926 40000
rect 3974 39200 4030 40000
rect 5078 39200 5134 40000
rect 6182 39200 6238 40000
rect 7286 39200 7342 40000
rect 8390 39200 8446 40000
rect 9494 39200 9550 40000
rect 10598 39200 10654 40000
rect 11702 39200 11758 40000
rect 12806 39200 12862 40000
rect 13910 39200 13966 40000
rect 15014 39200 15070 40000
rect 16118 39200 16174 40000
rect 17222 39200 17278 40000
rect 18326 39200 18382 40000
rect 19430 39200 19486 40000
rect 20534 39200 20590 40000
rect 21638 39200 21694 40000
rect 22742 39200 22798 40000
rect 23846 39200 23902 40000
rect 24950 39200 25006 40000
rect 26054 39200 26110 40000
rect 27158 39200 27214 40000
rect 28262 39200 28318 40000
rect 29366 39200 29422 40000
rect 30470 39200 30526 40000
rect 31574 39200 31630 40000
rect 32678 39200 32734 40000
rect 33782 39200 33838 40000
rect 34886 39200 34942 40000
rect 35990 39200 36046 40000
rect 37094 39200 37150 40000
rect 38198 39200 38254 40000
rect 39302 39200 39358 40000
rect 2318 0 2374 800
rect 2870 0 2926 800
rect 3422 0 3478 800
rect 3974 0 4030 800
rect 4526 0 4582 800
rect 5078 0 5134 800
rect 5630 0 5686 800
rect 6182 0 6238 800
rect 6734 0 6790 800
rect 7286 0 7342 800
rect 7838 0 7894 800
rect 8390 0 8446 800
rect 8942 0 8998 800
rect 9494 0 9550 800
rect 10046 0 10102 800
rect 10598 0 10654 800
rect 11150 0 11206 800
rect 11702 0 11758 800
rect 12254 0 12310 800
rect 12806 0 12862 800
rect 13358 0 13414 800
rect 13910 0 13966 800
rect 14462 0 14518 800
rect 15014 0 15070 800
rect 15566 0 15622 800
rect 16118 0 16174 800
rect 16670 0 16726 800
rect 17222 0 17278 800
rect 17774 0 17830 800
rect 18326 0 18382 800
rect 18878 0 18934 800
rect 19430 0 19486 800
rect 19982 0 20038 800
rect 20534 0 20590 800
rect 21086 0 21142 800
rect 21638 0 21694 800
rect 22190 0 22246 800
rect 22742 0 22798 800
rect 23294 0 23350 800
rect 23846 0 23902 800
rect 24398 0 24454 800
rect 24950 0 25006 800
rect 25502 0 25558 800
rect 26054 0 26110 800
rect 26606 0 26662 800
rect 27158 0 27214 800
rect 27710 0 27766 800
rect 28262 0 28318 800
rect 28814 0 28870 800
rect 29366 0 29422 800
rect 29918 0 29974 800
rect 30470 0 30526 800
rect 31022 0 31078 800
rect 31574 0 31630 800
rect 32126 0 32182 800
rect 32678 0 32734 800
rect 33230 0 33286 800
rect 33782 0 33838 800
rect 34334 0 34390 800
rect 34886 0 34942 800
rect 35438 0 35494 800
rect 35990 0 36046 800
rect 36542 0 36598 800
rect 37094 0 37150 800
rect 37646 0 37702 800
<< obsm2 >>
rect 774 39144 1710 39200
rect 1878 39144 2814 39200
rect 2982 39144 3918 39200
rect 4086 39144 5022 39200
rect 5190 39144 6126 39200
rect 6294 39144 7230 39200
rect 7398 39144 8334 39200
rect 8502 39144 9438 39200
rect 9606 39144 10542 39200
rect 10710 39144 11646 39200
rect 11814 39144 12750 39200
rect 12918 39144 13854 39200
rect 14022 39144 14958 39200
rect 15126 39144 16062 39200
rect 16230 39144 17166 39200
rect 17334 39144 18270 39200
rect 18438 39144 19374 39200
rect 19542 39144 20478 39200
rect 20646 39144 21582 39200
rect 21750 39144 22686 39200
rect 22854 39144 23790 39200
rect 23958 39144 24894 39200
rect 25062 39144 25998 39200
rect 26166 39144 27102 39200
rect 27270 39144 28206 39200
rect 28374 39144 29310 39200
rect 29478 39144 30414 39200
rect 30582 39144 31518 39200
rect 31686 39144 32622 39200
rect 32790 39144 33726 39200
rect 33894 39144 34830 39200
rect 34998 39144 35934 39200
rect 36102 39144 37038 39200
rect 37206 39144 38142 39200
rect 38310 39144 39246 39200
rect 664 856 39356 39144
rect 664 734 2262 856
rect 2430 734 2814 856
rect 2982 734 3366 856
rect 3534 734 3918 856
rect 4086 734 4470 856
rect 4638 734 5022 856
rect 5190 734 5574 856
rect 5742 734 6126 856
rect 6294 734 6678 856
rect 6846 734 7230 856
rect 7398 734 7782 856
rect 7950 734 8334 856
rect 8502 734 8886 856
rect 9054 734 9438 856
rect 9606 734 9990 856
rect 10158 734 10542 856
rect 10710 734 11094 856
rect 11262 734 11646 856
rect 11814 734 12198 856
rect 12366 734 12750 856
rect 12918 734 13302 856
rect 13470 734 13854 856
rect 14022 734 14406 856
rect 14574 734 14958 856
rect 15126 734 15510 856
rect 15678 734 16062 856
rect 16230 734 16614 856
rect 16782 734 17166 856
rect 17334 734 17718 856
rect 17886 734 18270 856
rect 18438 734 18822 856
rect 18990 734 19374 856
rect 19542 734 19926 856
rect 20094 734 20478 856
rect 20646 734 21030 856
rect 21198 734 21582 856
rect 21750 734 22134 856
rect 22302 734 22686 856
rect 22854 734 23238 856
rect 23406 734 23790 856
rect 23958 734 24342 856
rect 24510 734 24894 856
rect 25062 734 25446 856
rect 25614 734 25998 856
rect 26166 734 26550 856
rect 26718 734 27102 856
rect 27270 734 27654 856
rect 27822 734 28206 856
rect 28374 734 28758 856
rect 28926 734 29310 856
rect 29478 734 29862 856
rect 30030 734 30414 856
rect 30582 734 30966 856
rect 31134 734 31518 856
rect 31686 734 32070 856
rect 32238 734 32622 856
rect 32790 734 33174 856
rect 33342 734 33726 856
rect 33894 734 34278 856
rect 34446 734 34830 856
rect 34998 734 35382 856
rect 35550 734 35934 856
rect 36102 734 36486 856
rect 36654 734 37038 856
rect 37206 734 37590 856
rect 37758 734 39356 856
<< metal3 >>
rect 0 29928 800 30048
rect 0 9936 800 10056
<< obsm3 >>
rect 800 30128 35246 37569
rect 880 29848 35246 30128
rect 800 10136 35246 29848
rect 880 9856 35246 10136
rect 800 1803 35246 9856
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
<< labels >>
rlabel metal2 s 662 39200 718 40000 6 cw_ack
port 1 nsew signal input
rlabel metal2 s 1766 39200 1822 40000 6 cw_dir
port 2 nsew signal output
rlabel metal2 s 2870 39200 2926 40000 6 cw_err
port 3 nsew signal input
rlabel metal2 s 3974 39200 4030 40000 6 cw_io_i[0]
port 4 nsew signal input
rlabel metal2 s 15014 39200 15070 40000 6 cw_io_i[10]
port 5 nsew signal input
rlabel metal2 s 16118 39200 16174 40000 6 cw_io_i[11]
port 6 nsew signal input
rlabel metal2 s 17222 39200 17278 40000 6 cw_io_i[12]
port 7 nsew signal input
rlabel metal2 s 18326 39200 18382 40000 6 cw_io_i[13]
port 8 nsew signal input
rlabel metal2 s 19430 39200 19486 40000 6 cw_io_i[14]
port 9 nsew signal input
rlabel metal2 s 20534 39200 20590 40000 6 cw_io_i[15]
port 10 nsew signal input
rlabel metal2 s 5078 39200 5134 40000 6 cw_io_i[1]
port 11 nsew signal input
rlabel metal2 s 6182 39200 6238 40000 6 cw_io_i[2]
port 12 nsew signal input
rlabel metal2 s 7286 39200 7342 40000 6 cw_io_i[3]
port 13 nsew signal input
rlabel metal2 s 8390 39200 8446 40000 6 cw_io_i[4]
port 14 nsew signal input
rlabel metal2 s 9494 39200 9550 40000 6 cw_io_i[5]
port 15 nsew signal input
rlabel metal2 s 10598 39200 10654 40000 6 cw_io_i[6]
port 16 nsew signal input
rlabel metal2 s 11702 39200 11758 40000 6 cw_io_i[7]
port 17 nsew signal input
rlabel metal2 s 12806 39200 12862 40000 6 cw_io_i[8]
port 18 nsew signal input
rlabel metal2 s 13910 39200 13966 40000 6 cw_io_i[9]
port 19 nsew signal input
rlabel metal2 s 21638 39200 21694 40000 6 cw_io_o[0]
port 20 nsew signal output
rlabel metal2 s 32678 39200 32734 40000 6 cw_io_o[10]
port 21 nsew signal output
rlabel metal2 s 33782 39200 33838 40000 6 cw_io_o[11]
port 22 nsew signal output
rlabel metal2 s 34886 39200 34942 40000 6 cw_io_o[12]
port 23 nsew signal output
rlabel metal2 s 35990 39200 36046 40000 6 cw_io_o[13]
port 24 nsew signal output
rlabel metal2 s 37094 39200 37150 40000 6 cw_io_o[14]
port 25 nsew signal output
rlabel metal2 s 38198 39200 38254 40000 6 cw_io_o[15]
port 26 nsew signal output
rlabel metal2 s 22742 39200 22798 40000 6 cw_io_o[1]
port 27 nsew signal output
rlabel metal2 s 23846 39200 23902 40000 6 cw_io_o[2]
port 28 nsew signal output
rlabel metal2 s 24950 39200 25006 40000 6 cw_io_o[3]
port 29 nsew signal output
rlabel metal2 s 26054 39200 26110 40000 6 cw_io_o[4]
port 30 nsew signal output
rlabel metal2 s 27158 39200 27214 40000 6 cw_io_o[5]
port 31 nsew signal output
rlabel metal2 s 28262 39200 28318 40000 6 cw_io_o[6]
port 32 nsew signal output
rlabel metal2 s 29366 39200 29422 40000 6 cw_io_o[7]
port 33 nsew signal output
rlabel metal2 s 30470 39200 30526 40000 6 cw_io_o[8]
port 34 nsew signal output
rlabel metal2 s 31574 39200 31630 40000 6 cw_io_o[9]
port 35 nsew signal output
rlabel metal2 s 39302 39200 39358 40000 6 cw_req
port 36 nsew signal output
rlabel metal3 s 0 9936 800 10056 6 i_clk
port 37 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 i_rst
port 38 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 39 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 40 nsew ground bidirectional
rlabel metal2 s 2318 0 2374 800 6 wb_4_burst
port 41 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wb_8_burst
port 42 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wb_ack
port 43 nsew signal output
rlabel metal2 s 3974 0 4030 800 6 wb_adr[0]
port 44 nsew signal input
rlabel metal2 s 9494 0 9550 800 6 wb_adr[10]
port 45 nsew signal input
rlabel metal2 s 10046 0 10102 800 6 wb_adr[11]
port 46 nsew signal input
rlabel metal2 s 10598 0 10654 800 6 wb_adr[12]
port 47 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wb_adr[13]
port 48 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wb_adr[14]
port 49 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 wb_adr[15]
port 50 nsew signal input
rlabel metal2 s 12806 0 12862 800 6 wb_adr[16]
port 51 nsew signal input
rlabel metal2 s 13358 0 13414 800 6 wb_adr[17]
port 52 nsew signal input
rlabel metal2 s 13910 0 13966 800 6 wb_adr[18]
port 53 nsew signal input
rlabel metal2 s 14462 0 14518 800 6 wb_adr[19]
port 54 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wb_adr[1]
port 55 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wb_adr[20]
port 56 nsew signal input
rlabel metal2 s 15566 0 15622 800 6 wb_adr[21]
port 57 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 wb_adr[22]
port 58 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 wb_adr[23]
port 59 nsew signal input
rlabel metal2 s 5078 0 5134 800 6 wb_adr[2]
port 60 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wb_adr[3]
port 61 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wb_adr[4]
port 62 nsew signal input
rlabel metal2 s 6734 0 6790 800 6 wb_adr[5]
port 63 nsew signal input
rlabel metal2 s 7286 0 7342 800 6 wb_adr[6]
port 64 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wb_adr[7]
port 65 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wb_adr[8]
port 66 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wb_adr[9]
port 67 nsew signal input
rlabel metal2 s 17222 0 17278 800 6 wb_cyc
port 68 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wb_err
port 69 nsew signal output
rlabel metal2 s 18326 0 18382 800 6 wb_i_dat[0]
port 70 nsew signal output
rlabel metal2 s 23846 0 23902 800 6 wb_i_dat[10]
port 71 nsew signal output
rlabel metal2 s 24398 0 24454 800 6 wb_i_dat[11]
port 72 nsew signal output
rlabel metal2 s 24950 0 25006 800 6 wb_i_dat[12]
port 73 nsew signal output
rlabel metal2 s 25502 0 25558 800 6 wb_i_dat[13]
port 74 nsew signal output
rlabel metal2 s 26054 0 26110 800 6 wb_i_dat[14]
port 75 nsew signal output
rlabel metal2 s 26606 0 26662 800 6 wb_i_dat[15]
port 76 nsew signal output
rlabel metal2 s 18878 0 18934 800 6 wb_i_dat[1]
port 77 nsew signal output
rlabel metal2 s 19430 0 19486 800 6 wb_i_dat[2]
port 78 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 wb_i_dat[3]
port 79 nsew signal output
rlabel metal2 s 20534 0 20590 800 6 wb_i_dat[4]
port 80 nsew signal output
rlabel metal2 s 21086 0 21142 800 6 wb_i_dat[5]
port 81 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 wb_i_dat[6]
port 82 nsew signal output
rlabel metal2 s 22190 0 22246 800 6 wb_i_dat[7]
port 83 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 wb_i_dat[8]
port 84 nsew signal output
rlabel metal2 s 23294 0 23350 800 6 wb_i_dat[9]
port 85 nsew signal output
rlabel metal2 s 27158 0 27214 800 6 wb_o_dat[0]
port 86 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 wb_o_dat[10]
port 87 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 wb_o_dat[11]
port 88 nsew signal input
rlabel metal2 s 33782 0 33838 800 6 wb_o_dat[12]
port 89 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 wb_o_dat[13]
port 90 nsew signal input
rlabel metal2 s 34886 0 34942 800 6 wb_o_dat[14]
port 91 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wb_o_dat[15]
port 92 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wb_o_dat[1]
port 93 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wb_o_dat[2]
port 94 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 wb_o_dat[3]
port 95 nsew signal input
rlabel metal2 s 29366 0 29422 800 6 wb_o_dat[4]
port 96 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wb_o_dat[5]
port 97 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 wb_o_dat[6]
port 98 nsew signal input
rlabel metal2 s 31022 0 31078 800 6 wb_o_dat[7]
port 99 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 wb_o_dat[8]
port 100 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 wb_o_dat[9]
port 101 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 wb_sel[0]
port 102 nsew signal input
rlabel metal2 s 36542 0 36598 800 6 wb_sel[1]
port 103 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 wb_stb
port 104 nsew signal input
rlabel metal2 s 37646 0 37702 800 6 wb_we
port 105 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1508484
string GDS_FILE /home/piotro/ppcpu_caravel/openlane/wb_compressor/runs/22_09_13_14_04/results/signoff/wb_compressor.magic.gds
string GDS_START 302790
<< end >>

